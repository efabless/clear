magic
tech sky130A
magscale 1 2
timestamp 1625784080
<< locali >>
rect 17509 10591 17543 10761
rect 17451 10557 17543 10591
rect 19349 10047 19383 10217
rect 16129 9027 16163 9129
rect 18797 8823 18831 9061
rect 18153 7735 18187 7905
rect 11437 7191 11471 7293
rect 14565 6103 14599 6409
rect 12265 5627 12299 5797
rect 18153 5151 18187 5253
rect 21097 5219 21131 5321
rect 18613 5083 18647 5185
rect 11437 4607 11471 4777
rect 11989 3587 12023 3689
rect 13553 3519 13587 3689
rect 16405 3383 16439 3553
rect 7389 2907 7423 3077
rect 9597 1819 9631 2057
<< viali >>
rect 18981 20485 19015 20519
rect 19533 20485 19567 20519
rect 20269 20417 20303 20451
rect 5733 20349 5767 20383
rect 6561 20349 6595 20383
rect 17969 20349 18003 20383
rect 21281 20349 21315 20383
rect 18797 20281 18831 20315
rect 19349 20281 19383 20315
rect 20637 20281 20671 20315
rect 20821 20281 20855 20315
rect 21097 20281 21131 20315
rect 5917 20213 5951 20247
rect 17417 20213 17451 20247
rect 17141 20009 17175 20043
rect 17601 20009 17635 20043
rect 20085 20009 20119 20043
rect 18429 19941 18463 19975
rect 17417 19873 17451 19907
rect 18245 19873 18279 19907
rect 20269 19873 20303 19907
rect 20637 19873 20671 19907
rect 20821 19873 20855 19907
rect 21189 19873 21223 19907
rect 21373 19737 21407 19771
rect 19717 19465 19751 19499
rect 20177 19465 20211 19499
rect 20637 19465 20671 19499
rect 6745 19261 6779 19295
rect 12633 19261 12667 19295
rect 19901 19261 19935 19295
rect 20361 19261 20395 19295
rect 20821 19261 20855 19295
rect 6929 19193 6963 19227
rect 21189 19193 21223 19227
rect 21373 19193 21407 19227
rect 12817 19125 12851 19159
rect 11989 18921 12023 18955
rect 18705 18921 18739 18955
rect 20085 18921 20119 18955
rect 20821 18921 20855 18955
rect 11805 18785 11839 18819
rect 18521 18785 18555 18819
rect 19901 18785 19935 18819
rect 20637 18785 20671 18819
rect 21189 18785 21223 18819
rect 21373 18649 21407 18683
rect 20085 18377 20119 18411
rect 12357 18309 12391 18343
rect 9413 18173 9447 18207
rect 12173 18173 12207 18207
rect 19901 18173 19935 18207
rect 21189 18105 21223 18139
rect 21373 18105 21407 18139
rect 9597 18037 9631 18071
rect 20821 17833 20855 17867
rect 8125 17697 8159 17731
rect 20637 17697 20671 17731
rect 21189 17697 21223 17731
rect 21373 17561 21407 17595
rect 8309 17493 8343 17527
rect 12081 17289 12115 17323
rect 19809 17289 19843 17323
rect 20269 17289 20303 17323
rect 20821 17153 20855 17187
rect 11897 17085 11931 17119
rect 19625 17085 19659 17119
rect 20085 17085 20119 17119
rect 20637 17017 20671 17051
rect 21189 17017 21223 17051
rect 21373 17017 21407 17051
rect 18061 16745 18095 16779
rect 20361 16745 20395 16779
rect 20637 16745 20671 16779
rect 21189 16677 21223 16711
rect 17877 16609 17911 16643
rect 20177 16609 20211 16643
rect 20821 16609 20855 16643
rect 21373 16609 21407 16643
rect 20085 16201 20119 16235
rect 20821 16201 20855 16235
rect 19901 15997 19935 16031
rect 20637 15997 20671 16031
rect 21189 15929 21223 15963
rect 21373 15929 21407 15963
rect 14749 15657 14783 15691
rect 20269 15657 20303 15691
rect 20821 15589 20855 15623
rect 14565 15521 14599 15555
rect 20085 15521 20119 15555
rect 20637 15521 20671 15555
rect 21189 15521 21223 15555
rect 21281 15317 21315 15351
rect 12081 15113 12115 15147
rect 20637 15113 20671 15147
rect 11897 14909 11931 14943
rect 20821 14909 20855 14943
rect 21189 14841 21223 14875
rect 21373 14841 21407 14875
rect 9965 14569 9999 14603
rect 20361 14569 20395 14603
rect 20821 14569 20855 14603
rect 9321 14433 9355 14467
rect 9781 14433 9815 14467
rect 20177 14433 20211 14467
rect 20637 14433 20671 14467
rect 21189 14433 21223 14467
rect 9505 14297 9539 14331
rect 21373 14297 21407 14331
rect 19165 14229 19199 14263
rect 19809 14229 19843 14263
rect 19441 14025 19475 14059
rect 11345 13957 11379 13991
rect 19901 13957 19935 13991
rect 20361 13889 20395 13923
rect 11161 13821 11195 13855
rect 17601 13821 17635 13855
rect 18245 13821 18279 13855
rect 19257 13821 19291 13855
rect 19717 13821 19751 13855
rect 21189 13821 21223 13855
rect 18521 13753 18555 13787
rect 18981 13685 19015 13719
rect 13829 13481 13863 13515
rect 20361 13481 20395 13515
rect 20821 13481 20855 13515
rect 17356 13413 17390 13447
rect 21373 13413 21407 13447
rect 13645 13345 13679 13379
rect 17877 13345 17911 13379
rect 18613 13345 18647 13379
rect 19073 13345 19107 13379
rect 20177 13345 20211 13379
rect 20637 13345 20671 13379
rect 21189 13345 21223 13379
rect 17601 13277 17635 13311
rect 18797 13209 18831 13243
rect 19625 13209 19659 13243
rect 16221 13141 16255 13175
rect 18061 13141 18095 13175
rect 19257 13141 19291 13175
rect 16589 12937 16623 12971
rect 19809 12937 19843 12971
rect 20821 12937 20855 12971
rect 21281 12937 21315 12971
rect 20269 12869 20303 12903
rect 16129 12733 16163 12767
rect 16405 12733 16439 12767
rect 17141 12733 17175 12767
rect 19165 12733 19199 12767
rect 19625 12733 19659 12767
rect 20085 12733 20119 12767
rect 20637 12733 20671 12767
rect 21097 12733 21131 12767
rect 15761 12665 15795 12699
rect 17386 12665 17420 12699
rect 18797 12665 18831 12699
rect 18521 12597 18555 12631
rect 19349 12597 19383 12631
rect 20085 12393 20119 12427
rect 21005 12393 21039 12427
rect 18144 12325 18178 12359
rect 21281 12325 21315 12359
rect 15669 12257 15703 12291
rect 15936 12257 15970 12291
rect 17877 12257 17911 12291
rect 19901 12257 19935 12291
rect 20545 12257 20579 12291
rect 20821 12257 20855 12291
rect 17601 12189 17635 12223
rect 14749 12053 14783 12087
rect 15301 12053 15335 12087
rect 17049 12053 17083 12087
rect 19257 12053 19291 12087
rect 20361 12053 20395 12087
rect 18429 11849 18463 11883
rect 14933 11781 14967 11815
rect 16589 11781 16623 11815
rect 15577 11713 15611 11747
rect 17877 11713 17911 11747
rect 15117 11645 15151 11679
rect 16405 11645 16439 11679
rect 17233 11645 17267 11679
rect 18061 11645 18095 11679
rect 20094 11645 20128 11679
rect 20361 11645 20395 11679
rect 21005 11645 21039 11679
rect 1777 11577 1811 11611
rect 1685 11509 1719 11543
rect 2237 11509 2271 11543
rect 14381 11509 14415 11543
rect 15669 11509 15703 11543
rect 15761 11509 15795 11543
rect 16129 11509 16163 11543
rect 17417 11509 17451 11543
rect 17969 11509 18003 11543
rect 18981 11509 19015 11543
rect 20821 11509 20855 11543
rect 21281 11509 21315 11543
rect 13553 11305 13587 11339
rect 14013 11305 14047 11339
rect 16313 11305 16347 11339
rect 17141 11305 17175 11339
rect 17509 11305 17543 11339
rect 18981 11305 19015 11339
rect 19809 11305 19843 11339
rect 20269 11305 20303 11339
rect 20821 11237 20855 11271
rect 13645 11169 13679 11203
rect 14657 11169 14691 11203
rect 14924 11169 14958 11203
rect 18061 11169 18095 11203
rect 18889 11169 18923 11203
rect 20177 11169 20211 11203
rect 13461 11101 13495 11135
rect 16957 11101 16991 11135
rect 17049 11101 17083 11135
rect 19165 11101 19199 11135
rect 20361 11101 20395 11135
rect 16037 11033 16071 11067
rect 18521 11033 18555 11067
rect 18245 10965 18279 10999
rect 21281 10965 21315 10999
rect 14013 10761 14047 10795
rect 15669 10761 15703 10795
rect 17509 10761 17543 10795
rect 12633 10625 12667 10659
rect 17601 10625 17635 10659
rect 12357 10557 12391 10591
rect 14289 10557 14323 10591
rect 14545 10557 14579 10591
rect 15945 10557 15979 10591
rect 16405 10557 16439 10591
rect 17141 10557 17175 10591
rect 17417 10557 17451 10591
rect 17868 10557 17902 10591
rect 19257 10557 19291 10591
rect 19717 10557 19751 10591
rect 19973 10557 20007 10591
rect 12900 10489 12934 10523
rect 12173 10421 12207 10455
rect 16129 10421 16163 10455
rect 16589 10421 16623 10455
rect 17325 10421 17359 10455
rect 18981 10421 19015 10455
rect 19441 10421 19475 10455
rect 21097 10421 21131 10455
rect 11805 10217 11839 10251
rect 13737 10217 13771 10251
rect 15577 10217 15611 10251
rect 16589 10217 16623 10251
rect 19349 10217 19383 10251
rect 20821 10217 20855 10251
rect 12541 10149 12575 10183
rect 14565 10149 14599 10183
rect 18000 10149 18034 10183
rect 12173 10081 12207 10115
rect 12817 10081 12851 10115
rect 13277 10081 13311 10115
rect 15209 10081 15243 10115
rect 16221 10081 16255 10115
rect 18521 10081 18555 10115
rect 19257 10081 19291 10115
rect 19901 10081 19935 10115
rect 20729 10081 20763 10115
rect 15025 10013 15059 10047
rect 15117 10013 15151 10047
rect 15945 10013 15979 10047
rect 16129 10013 16163 10047
rect 18245 10013 18279 10047
rect 19349 10013 19383 10047
rect 20913 10013 20947 10047
rect 13001 9945 13035 9979
rect 20361 9945 20395 9979
rect 13461 9877 13495 9911
rect 16865 9877 16899 9911
rect 19073 9877 19107 9911
rect 20085 9877 20119 9911
rect 16405 9673 16439 9707
rect 11345 9605 11379 9639
rect 11897 9605 11931 9639
rect 17049 9605 17083 9639
rect 12449 9537 12483 9571
rect 18061 9537 18095 9571
rect 20729 9537 20763 9571
rect 11161 9469 11195 9503
rect 13645 9469 13679 9503
rect 14105 9469 14139 9503
rect 14749 9469 14783 9503
rect 15025 9469 15059 9503
rect 17969 9469 18003 9503
rect 19634 9469 19668 9503
rect 19901 9469 19935 9503
rect 21373 9469 21407 9503
rect 12265 9401 12299 9435
rect 12909 9401 12943 9435
rect 15292 9401 15326 9435
rect 17877 9401 17911 9435
rect 12357 9333 12391 9367
rect 13461 9333 13495 9367
rect 14289 9333 14323 9367
rect 14565 9333 14599 9367
rect 17509 9333 17543 9367
rect 18521 9333 18555 9367
rect 20177 9333 20211 9367
rect 20545 9333 20579 9367
rect 20637 9333 20671 9367
rect 21189 9333 21223 9367
rect 10057 9129 10091 9163
rect 11713 9129 11747 9163
rect 15945 9129 15979 9163
rect 16129 9129 16163 9163
rect 17877 9129 17911 9163
rect 12256 9061 12290 9095
rect 16466 9061 16500 9095
rect 18797 9061 18831 9095
rect 9689 8993 9723 9027
rect 10600 8993 10634 9027
rect 14821 8993 14855 9027
rect 16129 8993 16163 9027
rect 16221 8993 16255 9027
rect 18705 8993 18739 9027
rect 9413 8925 9447 8959
rect 9597 8925 9631 8959
rect 10333 8925 10367 8959
rect 11989 8925 12023 8959
rect 14013 8925 14047 8959
rect 14565 8925 14599 8959
rect 19625 8993 19659 9027
rect 21106 8993 21140 9027
rect 21373 8993 21407 9027
rect 18981 8925 19015 8959
rect 19993 8857 20027 8891
rect 13369 8789 13403 8823
rect 17601 8789 17635 8823
rect 18521 8789 18555 8823
rect 18797 8789 18831 8823
rect 8125 8585 8159 8619
rect 11161 8585 11195 8619
rect 17877 8585 17911 8619
rect 20729 8585 20763 8619
rect 16589 8517 16623 8551
rect 18337 8517 18371 8551
rect 17233 8449 17267 8483
rect 18889 8449 18923 8483
rect 9505 8381 9539 8415
rect 9781 8381 9815 8415
rect 10037 8381 10071 8415
rect 12725 8381 12759 8415
rect 12992 8381 13026 8415
rect 16405 8381 16439 8415
rect 18705 8381 18739 8415
rect 19349 8381 19383 8415
rect 19605 8381 19639 8415
rect 9238 8313 9272 8347
rect 14381 8313 14415 8347
rect 16129 8313 16163 8347
rect 17509 8313 17543 8347
rect 18797 8313 18831 8347
rect 21005 8313 21039 8347
rect 12081 8245 12115 8279
rect 12449 8245 12483 8279
rect 14105 8245 14139 8279
rect 17417 8245 17451 8279
rect 8677 8041 8711 8075
rect 9505 8041 9539 8075
rect 10885 8041 10919 8075
rect 11253 8041 11287 8075
rect 14013 8041 14047 8075
rect 15025 8041 15059 8075
rect 16313 8041 16347 8075
rect 20821 8041 20855 8075
rect 14933 7973 14967 8007
rect 15945 7973 15979 8007
rect 17702 7973 17736 8007
rect 20729 7973 20763 8007
rect 10241 7905 10275 7939
rect 11621 7905 11655 7939
rect 11888 7905 11922 7939
rect 13645 7905 13679 7939
rect 15853 7905 15887 7939
rect 17969 7905 18003 7939
rect 18153 7905 18187 7939
rect 18613 7905 18647 7939
rect 20085 7905 20119 7939
rect 10701 7837 10735 7871
rect 10793 7837 10827 7871
rect 13369 7837 13403 7871
rect 13553 7837 13587 7871
rect 15117 7837 15151 7871
rect 15761 7837 15795 7871
rect 14565 7769 14599 7803
rect 18705 7837 18739 7871
rect 18889 7837 18923 7871
rect 20913 7837 20947 7871
rect 19901 7769 19935 7803
rect 10057 7701 10091 7735
rect 13001 7701 13035 7735
rect 16589 7701 16623 7735
rect 18153 7701 18187 7735
rect 18245 7701 18279 7735
rect 20361 7701 20395 7735
rect 9505 7497 9539 7531
rect 9873 7497 9907 7531
rect 11897 7497 11931 7531
rect 16497 7497 16531 7531
rect 17877 7497 17911 7531
rect 19349 7497 19383 7531
rect 21281 7497 21315 7531
rect 10333 7429 10367 7463
rect 15117 7429 15151 7463
rect 19625 7429 19659 7463
rect 8953 7361 8987 7395
rect 10701 7361 10735 7395
rect 12449 7361 12483 7395
rect 14650 7361 14684 7395
rect 15945 7361 15979 7395
rect 17325 7361 17359 7395
rect 18153 7361 18187 7395
rect 18797 7361 18831 7395
rect 20085 7361 20119 7395
rect 20177 7361 20211 7395
rect 8493 7293 8527 7327
rect 10149 7293 10183 7327
rect 11437 7293 11471 7327
rect 12265 7293 12299 7327
rect 14933 7293 14967 7327
rect 19993 7293 20027 7327
rect 21005 7293 21039 7327
rect 10977 7225 11011 7259
rect 12357 7225 12391 7259
rect 13001 7225 13035 7259
rect 14412 7225 14446 7259
rect 9045 7157 9079 7191
rect 9137 7157 9171 7191
rect 10885 7157 10919 7191
rect 11345 7157 11379 7191
rect 11437 7157 11471 7191
rect 13277 7157 13311 7191
rect 15393 7157 15427 7191
rect 16037 7157 16071 7191
rect 16129 7157 16163 7191
rect 17417 7157 17451 7191
rect 17509 7157 17543 7191
rect 18889 7157 18923 7191
rect 18981 7157 19015 7191
rect 20821 7157 20855 7191
rect 8769 6953 8803 6987
rect 10701 6953 10735 6987
rect 12357 6953 12391 6987
rect 9321 6817 9355 6851
rect 9577 6817 9611 6851
rect 11233 6817 11267 6851
rect 12633 6817 12667 6851
rect 13461 6817 13495 6851
rect 14841 6817 14875 6851
rect 15557 6817 15591 6851
rect 17877 6817 17911 6851
rect 18144 6817 18178 6851
rect 20157 6817 20191 6851
rect 10977 6749 11011 6783
rect 13185 6749 13219 6783
rect 13369 6749 13403 6783
rect 15301 6749 15335 6783
rect 17509 6749 17543 6783
rect 19901 6749 19935 6783
rect 12817 6681 12851 6715
rect 13829 6681 13863 6715
rect 16681 6681 16715 6715
rect 17049 6681 17083 6715
rect 7941 6613 7975 6647
rect 8309 6613 8343 6647
rect 14565 6613 14599 6647
rect 15025 6613 15059 6647
rect 19257 6613 19291 6647
rect 21281 6613 21315 6647
rect 10425 6409 10459 6443
rect 11345 6409 11379 6443
rect 13461 6409 13495 6443
rect 13921 6409 13955 6443
rect 14565 6409 14599 6443
rect 14657 6409 14691 6443
rect 18521 6409 18555 6443
rect 20177 6409 20211 6443
rect 12449 6341 12483 6375
rect 12817 6273 12851 6307
rect 7389 6205 7423 6239
rect 9045 6205 9079 6239
rect 10701 6205 10735 6239
rect 11161 6205 11195 6239
rect 12265 6205 12299 6239
rect 13737 6205 13771 6239
rect 14381 6205 14415 6239
rect 7656 6137 7690 6171
rect 9290 6137 9324 6171
rect 13093 6137 13127 6171
rect 21005 6273 21039 6307
rect 16037 6205 16071 6239
rect 16405 6205 16439 6239
rect 17141 6205 17175 6239
rect 17397 6205 17431 6239
rect 18797 6205 18831 6239
rect 20913 6205 20947 6239
rect 15792 6137 15826 6171
rect 19064 6137 19098 6171
rect 20821 6137 20855 6171
rect 8769 6069 8803 6103
rect 10885 6069 10919 6103
rect 11989 6069 12023 6103
rect 13001 6069 13035 6103
rect 14197 6069 14231 6103
rect 14565 6069 14599 6103
rect 16589 6069 16623 6103
rect 20453 6069 20487 6103
rect 8309 5865 8343 5899
rect 8585 5865 8619 5899
rect 13737 5865 13771 5899
rect 15393 5865 15427 5899
rect 16129 5865 16163 5899
rect 16589 5865 16623 5899
rect 17141 5865 17175 5899
rect 20545 5865 20579 5899
rect 9321 5797 9355 5831
rect 11192 5797 11226 5831
rect 12265 5797 12299 5831
rect 15485 5797 15519 5831
rect 18797 5797 18831 5831
rect 21281 5797 21315 5831
rect 6653 5729 6687 5763
rect 7297 5729 7331 5763
rect 7941 5729 7975 5763
rect 8769 5729 8803 5763
rect 9597 5729 9631 5763
rect 11897 5729 11931 5763
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 11437 5661 11471 5695
rect 12624 5729 12658 5763
rect 14841 5729 14875 5763
rect 16497 5729 16531 5763
rect 17509 5729 17543 5763
rect 17601 5729 17635 5763
rect 18889 5729 18923 5763
rect 20453 5729 20487 5763
rect 12357 5661 12391 5695
rect 15301 5661 15335 5695
rect 16773 5661 16807 5695
rect 17693 5661 17727 5695
rect 18705 5661 18739 5695
rect 20637 5661 20671 5695
rect 10057 5593 10091 5627
rect 12081 5593 12115 5627
rect 12265 5593 12299 5627
rect 15853 5593 15887 5627
rect 18153 5593 18187 5627
rect 6837 5525 6871 5559
rect 9781 5525 9815 5559
rect 19257 5525 19291 5559
rect 19809 5525 19843 5559
rect 20085 5525 20119 5559
rect 21189 5525 21223 5559
rect 6929 5321 6963 5355
rect 9321 5321 9355 5355
rect 19625 5321 19659 5355
rect 21097 5321 21131 5355
rect 18153 5253 18187 5287
rect 18521 5253 18555 5287
rect 5733 5185 5767 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 9965 5185 9999 5219
rect 14105 5185 14139 5219
rect 15117 5185 15151 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 21097 5185 21131 5219
rect 21189 5185 21223 5219
rect 13562 5117 13596 5151
rect 13829 5117 13863 5151
rect 16589 5117 16623 5151
rect 17325 5117 17359 5151
rect 18153 5117 18187 5151
rect 18337 5117 18371 5151
rect 18981 5117 19015 5151
rect 19993 5117 20027 5151
rect 20085 5117 20119 5151
rect 20821 5117 20855 5151
rect 6101 5049 6135 5083
rect 8064 5049 8098 5083
rect 10232 5049 10266 5083
rect 15209 5049 15243 5083
rect 17785 5049 17819 5083
rect 17969 5049 18003 5083
rect 18613 5049 18647 5083
rect 18797 5049 18831 5083
rect 20637 5049 20671 5083
rect 6653 4981 6687 5015
rect 8861 4981 8895 5015
rect 8953 4981 8987 5015
rect 9689 4981 9723 5015
rect 11345 4981 11379 5015
rect 12081 4981 12115 5015
rect 12449 4981 12483 5015
rect 14565 4981 14599 5015
rect 15301 4981 15335 5015
rect 15669 4981 15703 5015
rect 15945 4981 15979 5015
rect 16405 4981 16439 5015
rect 17233 4981 17267 5015
rect 5365 4777 5399 4811
rect 5733 4777 5767 4811
rect 6469 4777 6503 4811
rect 8309 4777 8343 4811
rect 9321 4777 9355 4811
rect 11345 4777 11379 4811
rect 11437 4777 11471 4811
rect 11621 4777 11655 4811
rect 11989 4777 12023 4811
rect 13277 4777 13311 4811
rect 15485 4777 15519 4811
rect 15577 4777 15611 4811
rect 15945 4777 15979 4811
rect 19809 4777 19843 4811
rect 9781 4709 9815 4743
rect 4997 4641 5031 4675
rect 7113 4641 7147 4675
rect 7941 4641 7975 4675
rect 8585 4641 8619 4675
rect 9689 4641 9723 4675
rect 10977 4641 11011 4675
rect 13645 4709 13679 4743
rect 16405 4709 16439 4743
rect 16957 4709 16991 4743
rect 17417 4709 17451 4743
rect 20821 4709 20855 4743
rect 13001 4641 13035 4675
rect 14749 4641 14783 4675
rect 18817 4641 18851 4675
rect 19073 4641 19107 4675
rect 20177 4641 20211 4675
rect 21005 4641 21039 4675
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 9965 4573 9999 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 11437 4573 11471 4607
rect 12081 4573 12115 4607
rect 12173 4573 12207 4607
rect 13737 4573 13771 4607
rect 13829 4573 13863 4607
rect 15301 4573 15335 4607
rect 20269 4573 20303 4607
rect 20361 4573 20395 4607
rect 6101 4505 6135 4539
rect 14565 4505 14599 4539
rect 16221 4505 16255 4539
rect 16773 4505 16807 4539
rect 6837 4437 6871 4471
rect 7297 4437 7331 4471
rect 8769 4437 8803 4471
rect 12817 4437 12851 4471
rect 17693 4437 17727 4471
rect 4537 4233 4571 4267
rect 9229 4233 9263 4267
rect 21189 4233 21223 4267
rect 7113 4165 7147 4199
rect 10517 4097 10551 4131
rect 10701 4097 10735 4131
rect 12633 4097 12667 4131
rect 14105 4097 14139 4131
rect 15945 4097 15979 4131
rect 20729 4097 20763 4131
rect 6929 4029 6963 4063
rect 7389 4029 7423 4063
rect 7849 4029 7883 4063
rect 9505 4029 9539 4063
rect 9965 4029 9999 4063
rect 10793 4029 10827 4063
rect 11897 4029 11931 4063
rect 13921 4029 13955 4063
rect 17325 4029 17359 4063
rect 17877 4029 17911 4063
rect 19461 4029 19495 4063
rect 19717 4029 19751 4063
rect 20545 4029 20579 4063
rect 20637 4029 20671 4063
rect 21373 4029 21407 4063
rect 8094 3961 8128 3995
rect 12817 3961 12851 3995
rect 15678 3961 15712 3995
rect 16405 3961 16439 3995
rect 18061 3961 18095 3995
rect 4905 3893 4939 3927
rect 5365 3893 5399 3927
rect 5733 3893 5767 3927
rect 6009 3893 6043 3927
rect 6653 3893 6687 3927
rect 7573 3893 7607 3927
rect 9689 3893 9723 3927
rect 10149 3893 10183 3927
rect 11161 3893 11195 3927
rect 12081 3893 12115 3927
rect 12909 3893 12943 3927
rect 13277 3893 13311 3927
rect 13553 3893 13587 3927
rect 14013 3893 14047 3927
rect 14565 3893 14599 3927
rect 16313 3893 16347 3927
rect 17417 3893 17451 3927
rect 18337 3893 18371 3927
rect 20177 3893 20211 3927
rect 4077 3689 4111 3723
rect 7113 3689 7147 3723
rect 11621 3689 11655 3723
rect 11989 3689 12023 3723
rect 13553 3689 13587 3723
rect 14565 3689 14599 3723
rect 19165 3689 19199 3723
rect 20453 3689 20487 3723
rect 13216 3621 13250 3655
rect 6745 3553 6779 3587
rect 8502 3553 8536 3587
rect 9321 3553 9355 3587
rect 11078 3553 11112 3587
rect 11345 3553 11379 3587
rect 11989 3553 12023 3587
rect 13921 3621 13955 3655
rect 17702 3621 17736 3655
rect 21281 3621 21315 3655
rect 16057 3553 16091 3587
rect 16405 3553 16439 3587
rect 18797 3553 18831 3587
rect 6561 3485 6595 3519
rect 6653 3485 6687 3519
rect 8769 3485 8803 3519
rect 13461 3485 13495 3519
rect 13553 3485 13587 3519
rect 16313 3485 16347 3519
rect 5733 3417 5767 3451
rect 9505 3417 9539 3451
rect 17969 3485 18003 3519
rect 18613 3485 18647 3519
rect 18705 3485 18739 3519
rect 20545 3485 20579 3519
rect 20729 3485 20763 3519
rect 19809 3417 19843 3451
rect 1409 3349 1443 3383
rect 4353 3349 4387 3383
rect 4997 3349 5031 3383
rect 5365 3349 5399 3383
rect 6101 3349 6135 3383
rect 7389 3349 7423 3383
rect 9965 3349 9999 3383
rect 12081 3349 12115 3383
rect 13829 3349 13863 3383
rect 14933 3349 14967 3383
rect 16405 3349 16439 3383
rect 16589 3349 16623 3383
rect 20085 3349 20119 3383
rect 21189 3349 21223 3383
rect 4721 3145 4755 3179
rect 5181 3145 5215 3179
rect 6101 3145 6135 3179
rect 7481 3145 7515 3179
rect 9781 3145 9815 3179
rect 12449 3145 12483 3179
rect 19073 3145 19107 3179
rect 20269 3145 20303 3179
rect 20637 3145 20671 3179
rect 5641 3077 5675 3111
rect 7205 3077 7239 3111
rect 7389 3077 7423 3111
rect 21097 3077 21131 3111
rect 1409 2941 1443 2975
rect 3617 2941 3651 2975
rect 4537 2941 4571 2975
rect 4997 2941 5031 2975
rect 5457 2941 5491 2975
rect 5917 2941 5951 2975
rect 7021 2941 7055 2975
rect 8861 3009 8895 3043
rect 9137 3009 9171 3043
rect 15485 3009 15519 3043
rect 16497 3009 16531 3043
rect 17693 3009 17727 3043
rect 18521 3009 18555 3043
rect 19625 3009 19659 3043
rect 19809 3009 19843 3043
rect 11161 2941 11195 2975
rect 11989 2941 12023 2975
rect 13829 2941 13863 2975
rect 15209 2941 15243 2975
rect 17509 2941 17543 2975
rect 17601 2941 17635 2975
rect 18705 2941 18739 2975
rect 19901 2941 19935 2975
rect 1869 2873 1903 2907
rect 2973 2873 3007 2907
rect 7389 2873 7423 2907
rect 8594 2873 8628 2907
rect 10916 2873 10950 2907
rect 12173 2873 12207 2907
rect 13584 2873 13618 2907
rect 14289 2873 14323 2907
rect 15301 2873 15335 2907
rect 16221 2873 16255 2907
rect 16313 2873 16347 2907
rect 18613 2873 18647 2907
rect 20729 2873 20763 2907
rect 21281 2873 21315 2907
rect 1593 2805 1627 2839
rect 2237 2805 2271 2839
rect 2605 2805 2639 2839
rect 3893 2805 3927 2839
rect 6561 2805 6595 2839
rect 14197 2805 14231 2839
rect 14841 2805 14875 2839
rect 15853 2805 15887 2839
rect 17141 2805 17175 2839
rect 4721 2601 4755 2635
rect 7389 2601 7423 2635
rect 7941 2601 7975 2635
rect 8309 2601 8343 2635
rect 8401 2601 8435 2635
rect 9597 2601 9631 2635
rect 10701 2601 10735 2635
rect 11161 2601 11195 2635
rect 12817 2601 12851 2635
rect 13277 2601 13311 2635
rect 15117 2601 15151 2635
rect 16221 2601 16255 2635
rect 20085 2601 20119 2635
rect 1685 2533 1719 2567
rect 9965 2533 9999 2567
rect 10793 2533 10827 2567
rect 13737 2533 13771 2567
rect 16129 2533 16163 2567
rect 18153 2533 18187 2567
rect 18797 2533 18831 2567
rect 19257 2533 19291 2567
rect 2145 2465 2179 2499
rect 2605 2465 2639 2499
rect 3065 2465 3099 2499
rect 4077 2465 4111 2499
rect 4537 2465 4571 2499
rect 5089 2465 5123 2499
rect 5549 2465 5583 2499
rect 6009 2465 6043 2499
rect 6745 2465 6779 2499
rect 7205 2465 7239 2499
rect 9413 2465 9447 2499
rect 11437 2465 11471 2499
rect 12265 2465 12299 2499
rect 12909 2465 12943 2499
rect 17601 2465 17635 2499
rect 19441 2465 19475 2499
rect 20821 2465 20855 2499
rect 8585 2397 8619 2431
rect 10609 2397 10643 2431
rect 12725 2397 12759 2431
rect 14841 2397 14875 2431
rect 15025 2397 15059 2431
rect 16313 2397 16347 2431
rect 16865 2397 16899 2431
rect 20545 2397 20579 2431
rect 4261 2329 4295 2363
rect 6929 2329 6963 2363
rect 10149 2329 10183 2363
rect 13553 2329 13587 2363
rect 14197 2329 14231 2363
rect 15761 2329 15795 2363
rect 17417 2329 17451 2363
rect 17969 2329 18003 2363
rect 18981 2329 19015 2363
rect 1777 2261 1811 2295
rect 2329 2261 2363 2295
rect 2789 2261 2823 2295
rect 3249 2261 3283 2295
rect 5273 2261 5307 2295
rect 5733 2261 5767 2295
rect 6193 2261 6227 2295
rect 15485 2261 15519 2295
rect 9597 2057 9631 2091
rect 9597 1785 9631 1819
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 18966 20516 18972 20528
rect 18927 20488 18972 20516
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 19518 20516 19524 20528
rect 19479 20488 19524 20516
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20622 20448 20628 20460
rect 20303 20420 20628 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20622 20408 20628 20420
rect 20680 20448 20686 20460
rect 20680 20420 21312 20448
rect 20680 20408 20686 20420
rect 5718 20380 5724 20392
rect 5679 20352 5724 20380
rect 5718 20340 5724 20352
rect 5776 20380 5782 20392
rect 6549 20383 6607 20389
rect 6549 20380 6561 20383
rect 5776 20352 6561 20380
rect 5776 20340 5782 20352
rect 6549 20349 6561 20352
rect 6595 20349 6607 20383
rect 6549 20343 6607 20349
rect 17586 20340 17592 20392
rect 17644 20380 17650 20392
rect 21284 20389 21312 20420
rect 17957 20383 18015 20389
rect 17957 20380 17969 20383
rect 17644 20352 17969 20380
rect 17644 20340 17650 20352
rect 17957 20349 17969 20352
rect 18003 20349 18015 20383
rect 17957 20343 18015 20349
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 18782 20312 18788 20324
rect 18743 20284 18788 20312
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 19337 20315 19395 20321
rect 19337 20281 19349 20315
rect 19383 20312 19395 20315
rect 20070 20312 20076 20324
rect 19383 20284 20076 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 20070 20272 20076 20284
rect 20128 20272 20134 20324
rect 20625 20315 20683 20321
rect 20625 20281 20637 20315
rect 20671 20281 20683 20315
rect 20806 20312 20812 20324
rect 20767 20284 20812 20312
rect 20625 20275 20683 20281
rect 5902 20244 5908 20256
rect 5863 20216 5908 20244
rect 5902 20204 5908 20216
rect 5960 20204 5966 20256
rect 17402 20244 17408 20256
rect 17363 20216 17408 20244
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 20640 20244 20668 20275
rect 20806 20272 20812 20284
rect 20864 20272 20870 20324
rect 21082 20312 21088 20324
rect 21043 20284 21088 20312
rect 21082 20272 21088 20284
rect 21140 20272 21146 20324
rect 18012 20216 20668 20244
rect 18012 20204 18018 20216
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 17218 20040 17224 20052
rect 17175 20012 17224 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 17586 20040 17592 20052
rect 17547 20012 17592 20040
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 18782 20000 18788 20052
rect 18840 20040 18846 20052
rect 20073 20043 20131 20049
rect 20073 20040 20085 20043
rect 18840 20012 20085 20040
rect 18840 20000 18846 20012
rect 20073 20009 20085 20012
rect 20119 20009 20131 20043
rect 20073 20003 20131 20009
rect 17236 19904 17264 20000
rect 18417 19975 18475 19981
rect 18417 19941 18429 19975
rect 18463 19972 18475 19975
rect 18598 19972 18604 19984
rect 18463 19944 18604 19972
rect 18463 19941 18475 19944
rect 18417 19935 18475 19941
rect 18598 19932 18604 19944
rect 18656 19932 18662 19984
rect 17405 19907 17463 19913
rect 17405 19904 17417 19907
rect 17236 19876 17417 19904
rect 17405 19873 17417 19876
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 19702 19904 19708 19916
rect 18279 19876 19708 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 20254 19904 20260 19916
rect 20215 19876 20260 19904
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20622 19904 20628 19916
rect 20583 19876 20628 19904
rect 20622 19864 20628 19876
rect 20680 19864 20686 19916
rect 20806 19904 20812 19916
rect 20767 19876 20812 19904
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 21174 19904 21180 19916
rect 21135 19876 21180 19904
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 21358 19768 21364 19780
rect 21319 19740 21364 19768
rect 21358 19728 21364 19740
rect 21416 19728 21422 19780
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 19702 19496 19708 19508
rect 19663 19468 19708 19496
rect 19702 19456 19708 19468
rect 19760 19456 19766 19508
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 20165 19499 20223 19505
rect 20165 19496 20177 19499
rect 20128 19468 20177 19496
rect 20128 19456 20134 19468
rect 20165 19465 20177 19468
rect 20211 19465 20223 19499
rect 20622 19496 20628 19508
rect 20583 19468 20628 19496
rect 20165 19459 20223 19465
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 5902 19252 5908 19304
rect 5960 19292 5966 19304
rect 6733 19295 6791 19301
rect 6733 19292 6745 19295
rect 5960 19264 6745 19292
rect 5960 19252 5966 19264
rect 6733 19261 6745 19264
rect 6779 19261 6791 19295
rect 6733 19255 6791 19261
rect 11974 19252 11980 19304
rect 12032 19292 12038 19304
rect 12621 19295 12679 19301
rect 12621 19292 12633 19295
rect 12032 19264 12633 19292
rect 12032 19252 12038 19264
rect 12621 19261 12633 19264
rect 12667 19261 12679 19295
rect 12621 19255 12679 19261
rect 18690 19252 18696 19304
rect 18748 19292 18754 19304
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 18748 19264 19901 19292
rect 18748 19252 18754 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 20070 19252 20076 19304
rect 20128 19292 20134 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 20128 19264 20361 19292
rect 20128 19252 20134 19264
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 20806 19292 20812 19304
rect 20767 19264 20812 19292
rect 20349 19255 20407 19261
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 6917 19227 6975 19233
rect 6917 19193 6929 19227
rect 6963 19224 6975 19227
rect 7282 19224 7288 19236
rect 6963 19196 7288 19224
rect 6963 19193 6975 19196
rect 6917 19187 6975 19193
rect 7282 19184 7288 19196
rect 7340 19184 7346 19236
rect 16758 19184 16764 19236
rect 16816 19224 16822 19236
rect 21177 19227 21235 19233
rect 21177 19224 21189 19227
rect 16816 19196 21189 19224
rect 16816 19184 16822 19196
rect 21177 19193 21189 19196
rect 21223 19193 21235 19227
rect 21358 19224 21364 19236
rect 21319 19196 21364 19224
rect 21177 19187 21235 19193
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 12805 19159 12863 19165
rect 12805 19125 12817 19159
rect 12851 19156 12863 19159
rect 17954 19156 17960 19168
rect 12851 19128 17960 19156
rect 12851 19125 12863 19128
rect 12805 19119 12863 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 11974 18952 11980 18964
rect 11935 18924 11980 18952
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 18690 18952 18696 18964
rect 18651 18924 18696 18952
rect 18690 18912 18696 18924
rect 18748 18912 18754 18964
rect 20070 18952 20076 18964
rect 20031 18924 20076 18952
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 20809 18955 20867 18961
rect 20809 18921 20821 18955
rect 20855 18952 20867 18955
rect 21174 18952 21180 18964
rect 20855 18924 21180 18952
rect 20855 18921 20867 18924
rect 20809 18915 20867 18921
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 11793 18819 11851 18825
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 11974 18816 11980 18828
rect 11839 18788 11980 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 11974 18776 11980 18788
rect 12032 18776 12038 18828
rect 18509 18819 18567 18825
rect 18509 18785 18521 18819
rect 18555 18816 18567 18819
rect 18598 18816 18604 18828
rect 18555 18788 18604 18816
rect 18555 18785 18567 18788
rect 18509 18779 18567 18785
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 19610 18776 19616 18828
rect 19668 18816 19674 18828
rect 19889 18819 19947 18825
rect 19889 18816 19901 18819
rect 19668 18788 19901 18816
rect 19668 18776 19674 18788
rect 19889 18785 19901 18788
rect 19935 18785 19947 18819
rect 20622 18816 20628 18828
rect 20583 18788 20628 18816
rect 19889 18779 19947 18785
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 21174 18816 21180 18828
rect 21135 18788 21180 18816
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 21358 18680 21364 18692
rect 21319 18652 21364 18680
rect 21358 18640 21364 18652
rect 21416 18640 21422 18692
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 20073 18411 20131 18417
rect 20073 18377 20085 18411
rect 20119 18408 20131 18411
rect 20254 18408 20260 18420
rect 20119 18380 20260 18408
rect 20119 18377 20131 18380
rect 20073 18371 20131 18377
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 12345 18343 12403 18349
rect 12345 18309 12357 18343
rect 12391 18340 12403 18343
rect 16758 18340 16764 18352
rect 12391 18312 16764 18340
rect 12391 18309 12403 18312
rect 12345 18303 12403 18309
rect 16758 18300 16764 18312
rect 16816 18300 16822 18352
rect 9401 18207 9459 18213
rect 9401 18173 9413 18207
rect 9447 18204 9459 18207
rect 9490 18204 9496 18216
rect 9447 18176 9496 18204
rect 9447 18173 9459 18176
rect 9401 18167 9459 18173
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 12158 18204 12164 18216
rect 12119 18176 12164 18204
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18204 19947 18207
rect 19978 18204 19984 18216
rect 19935 18176 19984 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 20806 18204 20812 18216
rect 20088 18176 20812 18204
rect 20088 18136 20116 18176
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 9600 18108 20116 18136
rect 9600 18077 9628 18108
rect 20254 18096 20260 18148
rect 20312 18136 20318 18148
rect 21177 18139 21235 18145
rect 21177 18136 21189 18139
rect 20312 18108 21189 18136
rect 20312 18096 20318 18108
rect 21177 18105 21189 18108
rect 21223 18105 21235 18139
rect 21358 18136 21364 18148
rect 21319 18108 21364 18136
rect 21177 18099 21235 18105
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 9585 18071 9643 18077
rect 9585 18037 9597 18071
rect 9631 18037 9643 18071
rect 9585 18031 9643 18037
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 20809 17867 20867 17873
rect 20809 17833 20821 17867
rect 20855 17864 20867 17867
rect 21174 17864 21180 17876
rect 20855 17836 21180 17864
rect 20855 17833 20867 17836
rect 20809 17827 20867 17833
rect 21174 17824 21180 17836
rect 21232 17824 21238 17876
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17728 8171 17731
rect 8294 17728 8300 17740
rect 8159 17700 8300 17728
rect 8159 17697 8171 17700
rect 8113 17691 8171 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 20625 17731 20683 17737
rect 20625 17728 20637 17731
rect 19852 17700 20637 17728
rect 19852 17688 19858 17700
rect 20625 17697 20637 17700
rect 20671 17697 20683 17731
rect 20625 17691 20683 17697
rect 21177 17731 21235 17737
rect 21177 17697 21189 17731
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 21192 17660 21220 17691
rect 20404 17632 21220 17660
rect 20404 17620 20410 17632
rect 21358 17592 21364 17604
rect 21319 17564 21364 17592
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 8297 17527 8355 17533
rect 8297 17493 8309 17527
rect 8343 17524 8355 17527
rect 20622 17524 20628 17536
rect 8343 17496 20628 17524
rect 8343 17493 8355 17496
rect 8297 17487 8355 17493
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 12069 17323 12127 17329
rect 12069 17289 12081 17323
rect 12115 17320 12127 17323
rect 12158 17320 12164 17332
rect 12115 17292 12164 17320
rect 12115 17289 12127 17292
rect 12069 17283 12127 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 19794 17320 19800 17332
rect 19755 17292 19800 17320
rect 19794 17280 19800 17292
rect 19852 17280 19858 17332
rect 20254 17320 20260 17332
rect 20215 17292 20260 17320
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 20806 17184 20812 17196
rect 20767 17156 20812 17184
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 11790 17076 11796 17128
rect 11848 17116 11854 17128
rect 11885 17119 11943 17125
rect 11885 17116 11897 17119
rect 11848 17088 11897 17116
rect 11848 17076 11854 17088
rect 11885 17085 11897 17088
rect 11931 17085 11943 17119
rect 11885 17079 11943 17085
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 19613 17119 19671 17125
rect 19613 17116 19625 17119
rect 13872 17088 19625 17116
rect 13872 17076 13878 17088
rect 19613 17085 19625 17088
rect 19659 17085 19671 17119
rect 20070 17116 20076 17128
rect 20031 17088 20076 17116
rect 19613 17079 19671 17085
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20622 17048 20628 17060
rect 20583 17020 20628 17048
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 21174 17048 21180 17060
rect 21135 17020 21180 17048
rect 21174 17008 21180 17020
rect 21232 17008 21238 17060
rect 21361 17051 21419 17057
rect 21361 17017 21373 17051
rect 21407 17048 21419 17051
rect 21450 17048 21456 17060
rect 21407 17020 21456 17048
rect 21407 17017 21419 17020
rect 21361 17011 21419 17017
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 18049 16779 18107 16785
rect 18049 16745 18061 16779
rect 18095 16776 18107 16779
rect 20070 16776 20076 16788
rect 18095 16748 20076 16776
rect 18095 16745 18107 16748
rect 18049 16739 18107 16745
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 20622 16776 20628 16788
rect 20583 16748 20628 16776
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 20254 16668 20260 16720
rect 20312 16708 20318 16720
rect 21177 16711 21235 16717
rect 21177 16708 21189 16711
rect 20312 16680 21189 16708
rect 20312 16668 20318 16680
rect 21177 16677 21189 16680
rect 21223 16677 21235 16711
rect 21177 16671 21235 16677
rect 17678 16600 17684 16652
rect 17736 16640 17742 16652
rect 17865 16643 17923 16649
rect 17865 16640 17877 16643
rect 17736 16612 17877 16640
rect 17736 16600 17742 16612
rect 17865 16609 17877 16612
rect 17911 16609 17923 16643
rect 17865 16603 17923 16609
rect 17954 16600 17960 16652
rect 18012 16640 18018 16652
rect 20162 16640 20168 16652
rect 18012 16612 20024 16640
rect 20123 16612 20168 16640
rect 18012 16600 18018 16612
rect 19996 16572 20024 16612
rect 20162 16600 20168 16612
rect 20220 16600 20226 16652
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 20272 16612 20821 16640
rect 20272 16572 20300 16612
rect 20809 16609 20821 16612
rect 20855 16609 20867 16643
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 20809 16603 20867 16609
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 19996 16544 20300 16572
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 20073 16235 20131 16241
rect 20073 16201 20085 16235
rect 20119 16232 20131 16235
rect 20162 16232 20168 16244
rect 20119 16204 20168 16232
rect 20119 16201 20131 16204
rect 20073 16195 20131 16201
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21174 16232 21180 16244
rect 20855 16204 21180 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 16574 15988 16580 16040
rect 16632 16028 16638 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 16632 16000 19901 16028
rect 16632 15988 16638 16000
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 16022 15920 16028 15972
rect 16080 15960 16086 15972
rect 20640 15960 20668 15991
rect 16080 15932 20668 15960
rect 21177 15963 21235 15969
rect 16080 15920 16086 15932
rect 21177 15929 21189 15963
rect 21223 15929 21235 15963
rect 21358 15960 21364 15972
rect 21319 15932 21364 15960
rect 21177 15923 21235 15929
rect 20438 15852 20444 15904
rect 20496 15892 20502 15904
rect 21192 15892 21220 15923
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 20496 15864 21220 15892
rect 20496 15852 20502 15864
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 17954 15688 17960 15700
rect 14783 15660 17960 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 20254 15688 20260 15700
rect 20215 15660 20260 15688
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 20806 15620 20812 15632
rect 20767 15592 20812 15620
rect 20806 15580 20812 15592
rect 20864 15580 20870 15632
rect 14550 15552 14556 15564
rect 14511 15524 14556 15552
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 20070 15552 20076 15564
rect 20031 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 20622 15552 20628 15564
rect 20583 15524 20628 15552
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 21174 15552 21180 15564
rect 21135 15524 21180 15552
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 12069 15147 12127 15153
rect 12069 15113 12081 15147
rect 12115 15144 12127 15147
rect 16022 15144 16028 15156
rect 12115 15116 16028 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 20622 15144 20628 15156
rect 20583 15116 20628 15144
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 11882 14940 11888 14952
rect 11843 14912 11888 14940
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 20806 14940 20812 14952
rect 20767 14912 20812 14940
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 20346 14832 20352 14884
rect 20404 14872 20410 14884
rect 21177 14875 21235 14881
rect 21177 14872 21189 14875
rect 20404 14844 21189 14872
rect 20404 14832 20410 14844
rect 21177 14841 21189 14844
rect 21223 14841 21235 14875
rect 21177 14835 21235 14841
rect 21361 14875 21419 14881
rect 21361 14841 21373 14875
rect 21407 14872 21419 14875
rect 21450 14872 21456 14884
rect 21407 14844 21456 14872
rect 21407 14841 21419 14844
rect 21361 14835 21419 14841
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 9953 14603 10011 14609
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 20070 14600 20076 14612
rect 9999 14572 20076 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20349 14603 20407 14609
rect 20349 14569 20361 14603
rect 20395 14600 20407 14603
rect 20438 14600 20444 14612
rect 20395 14572 20444 14600
rect 20395 14569 20407 14572
rect 20349 14563 20407 14569
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 20809 14603 20867 14609
rect 20809 14569 20821 14603
rect 20855 14600 20867 14603
rect 21174 14600 21180 14612
rect 20855 14572 21180 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 8846 14424 8852 14476
rect 8904 14464 8910 14476
rect 9309 14467 9367 14473
rect 9309 14464 9321 14467
rect 8904 14436 9321 14464
rect 8904 14424 8910 14436
rect 9309 14433 9321 14436
rect 9355 14433 9367 14467
rect 9766 14464 9772 14476
rect 9727 14436 9772 14464
rect 9309 14427 9367 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 16356 14436 20177 14464
rect 16356 14424 16362 14436
rect 20165 14433 20177 14436
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 20625 14467 20683 14473
rect 20625 14433 20637 14467
rect 20671 14433 20683 14467
rect 21174 14464 21180 14476
rect 21135 14436 21180 14464
rect 20625 14427 20683 14433
rect 17954 14356 17960 14408
rect 18012 14396 18018 14408
rect 20640 14396 20668 14427
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 18012 14368 20668 14396
rect 18012 14356 18018 14368
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 20806 14328 20812 14340
rect 9539 14300 20812 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 21358 14328 21364 14340
rect 21319 14300 21364 14328
rect 21358 14288 21364 14300
rect 21416 14288 21422 14340
rect 18874 14220 18880 14272
rect 18932 14260 18938 14272
rect 19153 14263 19211 14269
rect 19153 14260 19165 14263
rect 18932 14232 19165 14260
rect 18932 14220 18938 14232
rect 19153 14229 19165 14232
rect 19199 14229 19211 14263
rect 19153 14223 19211 14229
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 19797 14263 19855 14269
rect 19797 14260 19809 14263
rect 19300 14232 19809 14260
rect 19300 14220 19306 14232
rect 19797 14229 19809 14232
rect 19843 14229 19855 14263
rect 19797 14223 19855 14229
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 20530 14056 20536 14068
rect 19475 14028 20536 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 11333 13991 11391 13997
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 16298 13988 16304 14000
rect 11379 13960 16304 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 19889 13991 19947 13997
rect 19889 13957 19901 13991
rect 19935 13988 19947 13991
rect 20990 13988 20996 14000
rect 19935 13960 20996 13988
rect 19935 13957 19947 13960
rect 19889 13951 19947 13957
rect 20990 13948 20996 13960
rect 21048 13948 21054 14000
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 17184 13892 20361 13920
rect 17184 13880 17190 13892
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 12158 13852 12164 13864
rect 11195 13824 12164 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 17770 13852 17776 13864
rect 17635 13824 17776 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13852 18291 13855
rect 18690 13852 18696 13864
rect 18279 13824 18696 13852
rect 18279 13821 18291 13824
rect 18233 13815 18291 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 18874 13812 18880 13864
rect 18932 13852 18938 13864
rect 19245 13855 19303 13861
rect 19245 13852 19257 13855
rect 18932 13824 19257 13852
rect 18932 13812 18938 13824
rect 19245 13821 19257 13824
rect 19291 13821 19303 13855
rect 19245 13815 19303 13821
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19392 13824 19717 13852
rect 19392 13812 19398 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 20898 13812 20904 13864
rect 20956 13852 20962 13864
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 20956 13824 21189 13852
rect 20956 13812 20962 13824
rect 21177 13821 21189 13824
rect 21223 13852 21235 13855
rect 21542 13852 21548 13864
rect 21223 13824 21548 13852
rect 21223 13821 21235 13824
rect 21177 13815 21235 13821
rect 21542 13812 21548 13824
rect 21600 13812 21606 13864
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 18506 13784 18512 13796
rect 8628 13756 18512 13784
rect 8628 13744 8634 13756
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 18969 13719 19027 13725
rect 18969 13685 18981 13719
rect 19015 13716 19027 13719
rect 19058 13716 19064 13728
rect 19015 13688 19064 13716
rect 19015 13685 19027 13688
rect 18969 13679 19027 13685
rect 19058 13676 19064 13688
rect 19116 13676 19122 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 17954 13512 17960 13524
rect 13863 13484 17960 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 20346 13512 20352 13524
rect 20307 13484 20352 13512
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 20809 13515 20867 13521
rect 20809 13481 20821 13515
rect 20855 13512 20867 13515
rect 21174 13512 21180 13524
rect 20855 13484 21180 13512
rect 20855 13481 20867 13484
rect 20809 13475 20867 13481
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 17402 13453 17408 13456
rect 17344 13447 17408 13453
rect 17344 13413 17356 13447
rect 17390 13413 17408 13447
rect 17344 13407 17408 13413
rect 17402 13404 17408 13407
rect 17460 13404 17466 13456
rect 18690 13444 18696 13456
rect 17880 13416 18696 13444
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 17880 13385 17908 13416
rect 18690 13404 18696 13416
rect 18748 13404 18754 13456
rect 21358 13444 21364 13456
rect 21319 13416 21364 13444
rect 21358 13404 21364 13416
rect 21416 13404 21422 13456
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13320 13348 13645 13376
rect 13320 13336 13326 13348
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13345 17923 13379
rect 17865 13339 17923 13345
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 18601 13379 18659 13385
rect 18601 13376 18613 13379
rect 18564 13348 18613 13376
rect 18564 13336 18570 13348
rect 18601 13345 18613 13348
rect 18647 13345 18659 13379
rect 19058 13376 19064 13388
rect 19019 13348 19064 13376
rect 18601 13339 18659 13345
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 20162 13376 20168 13388
rect 20123 13348 20168 13376
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 20622 13376 20628 13388
rect 20583 13348 20628 13376
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 21177 13379 21235 13385
rect 21177 13345 21189 13379
rect 21223 13345 21235 13379
rect 21177 13339 21235 13345
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13277 17647 13311
rect 20806 13308 20812 13320
rect 17589 13271 17647 13277
rect 19076 13280 20812 13308
rect 17604 13240 17632 13271
rect 17862 13240 17868 13252
rect 17604 13212 17868 13240
rect 17862 13200 17868 13212
rect 17920 13240 17926 13252
rect 18785 13243 18843 13249
rect 18785 13240 18797 13243
rect 17920 13212 18797 13240
rect 17920 13200 17926 13212
rect 18785 13209 18797 13212
rect 18831 13209 18843 13243
rect 18785 13203 18843 13209
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 16209 13175 16267 13181
rect 16209 13172 16221 13175
rect 16080 13144 16221 13172
rect 16080 13132 16086 13144
rect 16209 13141 16221 13144
rect 16255 13141 16267 13175
rect 16209 13135 16267 13141
rect 18049 13175 18107 13181
rect 18049 13141 18061 13175
rect 18095 13172 18107 13175
rect 19076 13172 19104 13280
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 21082 13268 21088 13320
rect 21140 13308 21146 13320
rect 21192 13308 21220 13339
rect 21140 13280 21220 13308
rect 21140 13268 21146 13280
rect 19150 13200 19156 13252
rect 19208 13240 19214 13252
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 19208 13212 19625 13240
rect 19208 13200 19214 13212
rect 19613 13209 19625 13212
rect 19659 13209 19671 13243
rect 19613 13203 19671 13209
rect 18095 13144 19104 13172
rect 19245 13175 19303 13181
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 19245 13141 19257 13175
rect 19291 13172 19303 13175
rect 20254 13172 20260 13184
rect 19291 13144 20260 13172
rect 19291 13141 19303 13144
rect 19245 13135 19303 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 16577 12971 16635 12977
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 18782 12968 18788 12980
rect 16623 12940 18788 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 19797 12971 19855 12977
rect 19797 12937 19809 12971
rect 19843 12968 19855 12971
rect 20622 12968 20628 12980
rect 19843 12940 20628 12968
rect 19843 12937 19855 12940
rect 19797 12931 19855 12937
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 20809 12971 20867 12977
rect 20809 12937 20821 12971
rect 20855 12968 20867 12971
rect 21082 12968 21088 12980
rect 20855 12940 21088 12968
rect 20855 12937 20867 12940
rect 20809 12931 20867 12937
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 20257 12903 20315 12909
rect 20257 12869 20269 12903
rect 20303 12869 20315 12903
rect 20257 12863 20315 12869
rect 16408 12804 17264 12832
rect 16408 12773 16436 12804
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16393 12767 16451 12773
rect 16393 12764 16405 12767
rect 16163 12736 16405 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16393 12733 16405 12736
rect 16439 12733 16451 12767
rect 16393 12727 16451 12733
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17129 12767 17187 12773
rect 17129 12764 17141 12767
rect 17000 12736 17141 12764
rect 17000 12724 17006 12736
rect 17129 12733 17141 12736
rect 17175 12733 17187 12767
rect 17236 12764 17264 12804
rect 18414 12764 18420 12776
rect 17236 12736 18420 12764
rect 17129 12727 17187 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18966 12724 18972 12776
rect 19024 12764 19030 12776
rect 19150 12764 19156 12776
rect 19024 12736 19156 12764
rect 19024 12724 19030 12736
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12764 19671 12767
rect 19702 12764 19708 12776
rect 19659 12736 19708 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 19702 12724 19708 12736
rect 19760 12724 19766 12776
rect 19886 12724 19892 12776
rect 19944 12764 19950 12776
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 19944 12736 20085 12764
rect 19944 12724 19950 12736
rect 20073 12733 20085 12736
rect 20119 12733 20131 12767
rect 20272 12764 20300 12863
rect 20625 12767 20683 12773
rect 20625 12764 20637 12767
rect 20272 12736 20637 12764
rect 20073 12727 20131 12733
rect 20625 12733 20637 12736
rect 20671 12733 20683 12767
rect 21082 12764 21088 12776
rect 21043 12736 21088 12764
rect 20625 12727 20683 12733
rect 21082 12724 21088 12736
rect 21140 12724 21146 12776
rect 15749 12699 15807 12705
rect 15749 12665 15761 12699
rect 15795 12696 15807 12699
rect 16850 12696 16856 12708
rect 15795 12668 16856 12696
rect 15795 12665 15807 12668
rect 15749 12659 15807 12665
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 17034 12656 17040 12708
rect 17092 12696 17098 12708
rect 17374 12699 17432 12705
rect 17374 12696 17386 12699
rect 17092 12668 17386 12696
rect 17092 12656 17098 12668
rect 17374 12665 17386 12668
rect 17420 12665 17432 12699
rect 17374 12659 17432 12665
rect 18046 12656 18052 12708
rect 18104 12696 18110 12708
rect 18785 12699 18843 12705
rect 18785 12696 18797 12699
rect 18104 12668 18797 12696
rect 18104 12656 18110 12668
rect 18785 12665 18797 12668
rect 18831 12665 18843 12699
rect 18785 12659 18843 12665
rect 18506 12628 18512 12640
rect 18467 12600 18512 12628
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 20622 12628 20628 12640
rect 19383 12600 20628 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20162 12424 20168 12436
rect 20119 12396 20168 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 20993 12427 21051 12433
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 21082 12424 21088 12436
rect 21039 12396 21088 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 15672 12328 16988 12356
rect 14642 12248 14648 12300
rect 14700 12288 14706 12300
rect 15672 12297 15700 12328
rect 16960 12300 16988 12328
rect 17954 12316 17960 12368
rect 18012 12356 18018 12368
rect 18132 12359 18190 12365
rect 18132 12356 18144 12359
rect 18012 12328 18144 12356
rect 18012 12316 18018 12328
rect 18132 12325 18144 12328
rect 18178 12356 18190 12359
rect 18506 12356 18512 12368
rect 18178 12328 18512 12356
rect 18178 12325 18190 12328
rect 18132 12319 18190 12325
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 20898 12316 20904 12368
rect 20956 12356 20962 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 20956 12328 21281 12356
rect 20956 12316 20962 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 15930 12297 15936 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14700 12260 15669 12288
rect 14700 12248 14706 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15924 12288 15936 12297
rect 15891 12260 15936 12288
rect 15657 12251 15715 12257
rect 15924 12251 15936 12260
rect 15930 12248 15936 12251
rect 15988 12248 15994 12300
rect 16942 12248 16948 12300
rect 17000 12288 17006 12300
rect 17310 12288 17316 12300
rect 17000 12260 17316 12288
rect 17000 12248 17006 12260
rect 17310 12248 17316 12260
rect 17368 12288 17374 12300
rect 17862 12288 17868 12300
rect 17368 12260 17868 12288
rect 17368 12248 17374 12260
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 19610 12248 19616 12300
rect 19668 12288 19674 12300
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 19668 12260 19901 12288
rect 19668 12248 19674 12260
rect 19889 12257 19901 12260
rect 19935 12257 19947 12291
rect 20530 12288 20536 12300
rect 20491 12260 20536 12288
rect 19889 12251 19947 12257
rect 20530 12248 20536 12260
rect 20588 12248 20594 12300
rect 20809 12291 20867 12297
rect 20809 12257 20821 12291
rect 20855 12257 20867 12291
rect 20809 12251 20867 12257
rect 17586 12220 17592 12232
rect 17547 12192 17592 12220
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 20824 12220 20852 12251
rect 18932 12192 20852 12220
rect 18932 12180 18938 12192
rect 14734 12084 14740 12096
rect 14695 12056 14740 12084
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15286 12084 15292 12096
rect 15247 12056 15292 12084
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 17000 12056 17049 12084
rect 17000 12044 17006 12056
rect 17037 12053 17049 12056
rect 17083 12053 17095 12087
rect 17037 12047 17095 12053
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18046 12084 18052 12096
rect 17920 12056 18052 12084
rect 17920 12044 17926 12056
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 19242 12084 19248 12096
rect 19203 12056 19248 12084
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 20346 12084 20352 12096
rect 20307 12056 20352 12084
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 18046 11880 18052 11892
rect 13596 11852 18052 11880
rect 13596 11840 13602 11852
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 18598 11880 18604 11892
rect 18463 11852 18604 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 13722 11772 13728 11824
rect 13780 11812 13786 11824
rect 14921 11815 14979 11821
rect 14921 11812 14933 11815
rect 13780 11784 14933 11812
rect 13780 11772 13786 11784
rect 14921 11781 14933 11784
rect 14967 11781 14979 11815
rect 14921 11775 14979 11781
rect 16577 11815 16635 11821
rect 16577 11781 16589 11815
rect 16623 11812 16635 11815
rect 18874 11812 18880 11824
rect 16623 11784 18880 11812
rect 16623 11781 16635 11784
rect 16577 11775 16635 11781
rect 18874 11772 18880 11784
rect 18932 11772 18938 11824
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15838 11744 15844 11756
rect 15611 11716 15844 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 17770 11744 17776 11756
rect 17236 11716 17776 11744
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11676 15163 11679
rect 15286 11676 15292 11688
rect 15151 11648 15292 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 15286 11636 15292 11648
rect 15344 11676 15350 11688
rect 16114 11676 16120 11688
rect 15344 11648 16120 11676
rect 15344 11636 15350 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11676 16451 11679
rect 16482 11676 16488 11688
rect 16439 11648 16488 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 17236 11685 17264 11716
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11744 17923 11747
rect 17954 11744 17960 11756
rect 17911 11716 17960 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 17586 11636 17592 11688
rect 17644 11676 17650 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17644 11648 18061 11676
rect 17644 11636 17650 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 20070 11676 20076 11688
rect 20128 11685 20134 11688
rect 19300 11648 20076 11676
rect 19300 11636 19306 11648
rect 20070 11636 20076 11648
rect 20128 11639 20140 11685
rect 20349 11679 20407 11685
rect 20349 11645 20361 11679
rect 20395 11645 20407 11679
rect 20990 11676 20996 11688
rect 20951 11648 20996 11676
rect 20349 11639 20407 11645
rect 20128 11636 20134 11639
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11577 1823 11611
rect 1765 11571 1823 11577
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 1780 11540 1808 11571
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 17034 11608 17040 11620
rect 9364 11580 17040 11608
rect 9364 11568 9370 11580
rect 17034 11568 17040 11580
rect 17092 11568 17098 11620
rect 19978 11608 19984 11620
rect 17236 11580 19984 11608
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 1780 11512 2237 11540
rect 2225 11509 2237 11512
rect 2271 11540 2283 11543
rect 8662 11540 8668 11552
rect 2271 11512 8668 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 13998 11500 14004 11552
rect 14056 11540 14062 11552
rect 14369 11543 14427 11549
rect 14369 11540 14381 11543
rect 14056 11512 14381 11540
rect 14056 11500 14062 11512
rect 14369 11509 14381 11512
rect 14415 11509 14427 11543
rect 15654 11540 15660 11552
rect 15615 11512 15660 11540
rect 14369 11503 14427 11509
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 16117 11543 16175 11549
rect 15804 11512 15849 11540
rect 15804 11500 15810 11512
rect 16117 11509 16129 11543
rect 16163 11540 16175 11543
rect 17236 11540 17264 11580
rect 19978 11568 19984 11580
rect 20036 11568 20042 11620
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 20364 11608 20392 11639
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 20220 11580 20392 11608
rect 20220 11568 20226 11580
rect 17402 11540 17408 11552
rect 16163 11512 17264 11540
rect 17363 11512 17408 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 17957 11543 18015 11549
rect 17957 11540 17969 11543
rect 17552 11512 17969 11540
rect 17552 11500 17558 11512
rect 17957 11509 17969 11512
rect 18003 11509 18015 11543
rect 17957 11503 18015 11509
rect 18969 11543 19027 11549
rect 18969 11509 18981 11543
rect 19015 11540 19027 11543
rect 19334 11540 19340 11552
rect 19015 11512 19340 11540
rect 19015 11509 19027 11512
rect 18969 11503 19027 11509
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11540 20867 11543
rect 20990 11540 20996 11552
rect 20855 11512 20996 11540
rect 20855 11509 20867 11512
rect 20809 11503 20867 11509
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 21266 11540 21272 11552
rect 21227 11512 21272 11540
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 13538 11336 13544 11348
rect 13499 11308 13544 11336
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 14001 11339 14059 11345
rect 14001 11305 14013 11339
rect 14047 11305 14059 11339
rect 14001 11299 14059 11305
rect 14016 11268 14044 11299
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 15804 11308 16313 11336
rect 15804 11296 15810 11308
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 17092 11308 17141 11336
rect 17092 11296 17098 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 17494 11336 17500 11348
rect 17455 11308 17500 11336
rect 17129 11299 17187 11305
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 18969 11339 19027 11345
rect 18969 11305 18981 11339
rect 19015 11336 19027 11339
rect 19797 11339 19855 11345
rect 19797 11336 19809 11339
rect 19015 11308 19809 11336
rect 19015 11305 19027 11308
rect 18969 11299 19027 11305
rect 19797 11305 19809 11308
rect 19843 11305 19855 11339
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 19797 11299 19855 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 14016 11240 17264 11268
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14642 11200 14648 11212
rect 14603 11172 14648 11200
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 14912 11203 14970 11209
rect 14912 11169 14924 11203
rect 14958 11200 14970 11203
rect 15470 11200 15476 11212
rect 14958 11172 15476 11200
rect 14958 11169 14970 11172
rect 14912 11163 14970 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 16850 11160 16856 11212
rect 16908 11200 16914 11212
rect 16908 11172 17080 11200
rect 16908 11160 16914 11172
rect 17052 11144 17080 11172
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11101 13507 11135
rect 16942 11132 16948 11144
rect 16903 11104 16948 11132
rect 13449 11095 13507 11101
rect 13464 11064 13492 11095
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17034 11092 17040 11144
rect 17092 11132 17098 11144
rect 17236 11132 17264 11240
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 20809 11271 20867 11277
rect 20809 11268 20821 11271
rect 17460 11240 18828 11268
rect 17460 11228 17466 11240
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17920 11172 18061 11200
rect 17920 11160 17926 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 18800 11132 18828 11240
rect 19168 11240 20821 11268
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19168 11200 19196 11240
rect 20809 11237 20821 11240
rect 20855 11237 20867 11271
rect 20809 11231 20867 11237
rect 18923 11172 19196 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19978 11200 19984 11212
rect 19300 11172 19984 11200
rect 19300 11160 19306 11172
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11200 20223 11203
rect 20714 11200 20720 11212
rect 20211 11172 20720 11200
rect 20211 11169 20223 11172
rect 20165 11163 20223 11169
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 19058 11132 19064 11144
rect 17092 11104 17137 11132
rect 17236 11104 18644 11132
rect 18800 11104 19064 11132
rect 17092 11092 17098 11104
rect 13906 11064 13912 11076
rect 13464 11036 13912 11064
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 16025 11067 16083 11073
rect 16025 11064 16037 11067
rect 15896 11036 16037 11064
rect 15896 11024 15902 11036
rect 16025 11033 16037 11036
rect 16071 11033 16083 11067
rect 16025 11027 16083 11033
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 16356 11036 18521 11064
rect 16356 11024 16362 11036
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 18616 11064 18644 11104
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 19153 11135 19211 11141
rect 19153 11101 19165 11135
rect 19199 11132 19211 11135
rect 19334 11132 19340 11144
rect 19199 11104 19340 11132
rect 19199 11101 19211 11104
rect 19153 11095 19211 11101
rect 19334 11092 19340 11104
rect 19392 11132 19398 11144
rect 19794 11132 19800 11144
rect 19392 11104 19800 11132
rect 19392 11092 19398 11104
rect 19794 11092 19800 11104
rect 19852 11092 19858 11144
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 20128 11104 20361 11132
rect 20128 11092 20134 11104
rect 20349 11101 20361 11104
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 19518 11064 19524 11076
rect 18616 11036 19524 11064
rect 18509 11027 18567 11033
rect 19518 11024 19524 11036
rect 19576 11024 19582 11076
rect 18233 10999 18291 11005
rect 18233 10965 18245 10999
rect 18279 10996 18291 10999
rect 19242 10996 19248 11008
rect 18279 10968 19248 10996
rect 18279 10965 18291 10968
rect 18233 10959 18291 10965
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 21266 10996 21272 11008
rect 20772 10968 21272 10996
rect 20772 10956 20778 10968
rect 21266 10956 21272 10968
rect 21324 10956 21330 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13964 10764 14013 10792
rect 13964 10752 13970 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 11698 10616 11704 10668
rect 11756 10656 11762 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 11756 10628 12633 10656
rect 11756 10616 11762 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 14016 10656 14044 10755
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 15528 10764 15669 10792
rect 15528 10752 15534 10764
rect 15657 10761 15669 10764
rect 15703 10761 15715 10795
rect 15657 10755 15715 10761
rect 17497 10795 17555 10801
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 19518 10792 19524 10804
rect 17543 10764 19524 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 17402 10684 17408 10736
rect 17460 10724 17466 10736
rect 17460 10696 17632 10724
rect 17460 10684 17466 10696
rect 17604 10665 17632 10696
rect 17589 10659 17647 10665
rect 14016 10628 14412 10656
rect 12621 10619 12679 10625
rect 12345 10591 12403 10597
rect 12345 10557 12357 10591
rect 12391 10557 12403 10591
rect 12345 10551 12403 10557
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10557 14335 10591
rect 14384 10588 14412 10628
rect 17589 10625 17601 10659
rect 17635 10625 17647 10659
rect 17589 10619 17647 10625
rect 14533 10591 14591 10597
rect 14533 10588 14545 10591
rect 14384 10560 14545 10588
rect 14277 10551 14335 10557
rect 14533 10557 14545 10560
rect 14579 10557 14591 10591
rect 15930 10588 15936 10600
rect 15891 10560 15936 10588
rect 14533 10551 14591 10557
rect 12158 10452 12164 10464
rect 12119 10424 12164 10452
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12360 10452 12388 10551
rect 12894 10529 12900 10532
rect 12888 10520 12900 10529
rect 12855 10492 12900 10520
rect 12888 10483 12900 10492
rect 12894 10480 12900 10483
rect 12952 10480 12958 10532
rect 14292 10520 14320 10551
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 17034 10588 17040 10600
rect 16439 10560 17040 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 17175 10560 17417 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 17405 10557 17417 10560
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 17853 10548 17859 10600
rect 17911 10588 17917 10600
rect 17911 10560 17956 10588
rect 17911 10548 17917 10560
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 19024 10560 19257 10588
rect 19024 10548 19030 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10557 19763 10591
rect 19705 10551 19763 10557
rect 14642 10520 14648 10532
rect 14292 10492 14648 10520
rect 14642 10480 14648 10492
rect 14700 10480 14706 10532
rect 16298 10520 16304 10532
rect 15488 10492 16304 10520
rect 15488 10452 15516 10492
rect 16298 10480 16304 10492
rect 16356 10480 16362 10532
rect 19720 10520 19748 10551
rect 19794 10548 19800 10600
rect 19852 10588 19858 10600
rect 19961 10591 20019 10597
rect 19961 10588 19973 10591
rect 19852 10560 19973 10588
rect 19852 10548 19858 10560
rect 19961 10557 19973 10560
rect 20007 10557 20019 10591
rect 19961 10551 20019 10557
rect 20070 10520 20076 10532
rect 16500 10492 19656 10520
rect 19720 10492 20076 10520
rect 12360 10424 15516 10452
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16500 10452 16528 10492
rect 16163 10424 16528 10452
rect 16577 10455 16635 10461
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16577 10421 16589 10455
rect 16623 10452 16635 10455
rect 16666 10452 16672 10464
rect 16623 10424 16672 10452
rect 16623 10421 16635 10424
rect 16577 10415 16635 10421
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 17313 10455 17371 10461
rect 17313 10421 17325 10455
rect 17359 10452 17371 10455
rect 18690 10452 18696 10464
rect 17359 10424 18696 10452
rect 17359 10421 17371 10424
rect 17313 10415 17371 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 18969 10455 19027 10461
rect 18969 10421 18981 10455
rect 19015 10452 19027 10455
rect 19334 10452 19340 10464
rect 19015 10424 19340 10452
rect 19015 10421 19027 10424
rect 18969 10415 19027 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19628 10452 19656 10492
rect 20070 10480 20076 10492
rect 20128 10480 20134 10532
rect 20898 10452 20904 10464
rect 19484 10424 19529 10452
rect 19628 10424 20904 10452
rect 19484 10412 19490 10424
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 21082 10452 21088 10464
rect 21043 10424 21088 10452
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 11793 10251 11851 10257
rect 11793 10217 11805 10251
rect 11839 10248 11851 10251
rect 13538 10248 13544 10260
rect 11839 10220 13544 10248
rect 11839 10217 11851 10220
rect 11793 10211 11851 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 13688 10220 13737 10248
rect 13688 10208 13694 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 15565 10251 15623 10257
rect 13725 10211 13783 10217
rect 14108 10220 14780 10248
rect 12529 10183 12587 10189
rect 12529 10149 12541 10183
rect 12575 10180 12587 10183
rect 12575 10152 13308 10180
rect 12575 10149 12587 10152
rect 12529 10143 12587 10149
rect 13280 10121 13308 10152
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10112 12219 10115
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12207 10084 12817 10112
rect 12207 10081 12219 10084
rect 12161 10075 12219 10081
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 14108 10112 14136 10220
rect 14553 10183 14611 10189
rect 14553 10149 14565 10183
rect 14599 10180 14611 10183
rect 14642 10180 14648 10192
rect 14599 10152 14648 10180
rect 14599 10149 14611 10152
rect 14553 10143 14611 10149
rect 14642 10140 14648 10152
rect 14700 10140 14706 10192
rect 14752 10180 14780 10220
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 15654 10248 15660 10260
rect 15611 10220 15660 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16574 10248 16580 10260
rect 16535 10220 16580 10248
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 18598 10248 18604 10260
rect 16684 10220 18604 10248
rect 16684 10180 16712 10220
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 19337 10251 19395 10257
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 20070 10248 20076 10260
rect 19383 10220 20076 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20806 10248 20812 10260
rect 20767 10220 20812 10248
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 14752 10152 16712 10180
rect 16758 10140 16764 10192
rect 16816 10180 16822 10192
rect 17402 10180 17408 10192
rect 16816 10152 17408 10180
rect 16816 10140 16822 10152
rect 17402 10140 17408 10152
rect 17460 10180 17466 10192
rect 17988 10183 18046 10189
rect 17460 10152 17724 10180
rect 17460 10140 17466 10152
rect 13311 10084 14136 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 12820 10044 12848 10075
rect 14182 10072 14188 10124
rect 14240 10112 14246 10124
rect 14734 10112 14740 10124
rect 14240 10084 14740 10112
rect 14240 10072 14246 10084
rect 14734 10072 14740 10084
rect 14792 10112 14798 10124
rect 15197 10115 15255 10121
rect 15197 10112 15209 10115
rect 14792 10084 15209 10112
rect 14792 10072 14798 10084
rect 15197 10081 15209 10084
rect 15243 10081 15255 10115
rect 15197 10075 15255 10081
rect 16209 10115 16267 10121
rect 16209 10081 16221 10115
rect 16255 10112 16267 10115
rect 17586 10112 17592 10124
rect 16255 10084 17592 10112
rect 16255 10081 16267 10084
rect 16209 10075 16267 10081
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17696 10112 17724 10152
rect 17988 10149 18000 10183
rect 18034 10180 18046 10183
rect 18034 10152 20024 10180
rect 18034 10149 18046 10152
rect 17988 10143 18046 10149
rect 17696 10084 18276 10112
rect 15013 10047 15071 10053
rect 12820 10016 14780 10044
rect 12989 9979 13047 9985
rect 12989 9945 13001 9979
rect 13035 9976 13047 9979
rect 14642 9976 14648 9988
rect 13035 9948 14648 9976
rect 13035 9945 13047 9948
rect 12989 9939 13047 9945
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 14274 9908 14280 9920
rect 13495 9880 14280 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 14752 9908 14780 10016
rect 15013 10013 15025 10047
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10044 15163 10047
rect 15286 10044 15292 10056
rect 15151 10016 15292 10044
rect 15151 10013 15163 10016
rect 15105 10007 15163 10013
rect 15028 9976 15056 10007
rect 15286 10004 15292 10016
rect 15344 10044 15350 10056
rect 15930 10044 15936 10056
rect 15344 10016 15608 10044
rect 15891 10016 15936 10044
rect 15344 10004 15350 10016
rect 15470 9976 15476 9988
rect 15028 9948 15476 9976
rect 15470 9936 15476 9948
rect 15528 9936 15534 9988
rect 15580 9976 15608 10016
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 16114 10044 16120 10056
rect 16075 10016 16120 10044
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 18248 10053 18276 10084
rect 18322 10072 18328 10124
rect 18380 10112 18386 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18380 10084 18521 10112
rect 18380 10072 18386 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 19242 10112 19248 10124
rect 19203 10084 19248 10112
rect 18509 10075 18567 10081
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 19794 10072 19800 10124
rect 19852 10112 19858 10124
rect 19889 10115 19947 10121
rect 19889 10112 19901 10115
rect 19852 10084 19901 10112
rect 19852 10072 19858 10084
rect 19889 10081 19901 10084
rect 19935 10081 19947 10115
rect 19889 10075 19947 10081
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10044 18291 10047
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 18279 10016 19349 10044
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 19337 10013 19349 10016
rect 19383 10013 19395 10047
rect 19996 10044 20024 10152
rect 20714 10112 20720 10124
rect 20675 10084 20720 10112
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 19996 10016 20913 10044
rect 19337 10007 19395 10013
rect 20901 10013 20913 10016
rect 20947 10044 20959 10047
rect 21082 10044 21088 10056
rect 20947 10016 21088 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 21082 10004 21088 10016
rect 21140 10004 21146 10056
rect 15838 9976 15844 9988
rect 15580 9948 15844 9976
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 17218 9976 17224 9988
rect 15948 9948 17224 9976
rect 15948 9908 15976 9948
rect 17218 9936 17224 9948
rect 17276 9936 17282 9988
rect 18782 9936 18788 9988
rect 18840 9976 18846 9988
rect 20349 9979 20407 9985
rect 20349 9976 20361 9979
rect 18840 9948 20361 9976
rect 18840 9936 18846 9948
rect 20349 9945 20361 9948
rect 20395 9945 20407 9979
rect 20349 9939 20407 9945
rect 16850 9908 16856 9920
rect 14752 9880 15976 9908
rect 16811 9880 16856 9908
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 19058 9908 19064 9920
rect 19019 9880 19064 9908
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 20073 9911 20131 9917
rect 20073 9877 20085 9911
rect 20119 9908 20131 9911
rect 20530 9908 20536 9920
rect 20119 9880 20536 9908
rect 20119 9877 20131 9880
rect 20073 9871 20131 9877
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 15286 9704 15292 9716
rect 13596 9676 15292 9704
rect 13596 9664 13602 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 16390 9704 16396 9716
rect 15988 9676 16396 9704
rect 15988 9664 15994 9676
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 18782 9664 18788 9716
rect 18840 9664 18846 9716
rect 11333 9639 11391 9645
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 11698 9636 11704 9648
rect 11379 9608 11704 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 11882 9636 11888 9648
rect 11843 9608 11888 9636
rect 11882 9596 11888 9608
rect 11940 9596 11946 9648
rect 17034 9636 17040 9648
rect 16947 9608 17040 9636
rect 17034 9596 17040 9608
rect 17092 9636 17098 9648
rect 17954 9636 17960 9648
rect 17092 9608 17960 9636
rect 17092 9596 17098 9608
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12308 9540 12449 9568
rect 12308 9528 12314 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 13648 9540 15148 9568
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 13648 9509 13676 9540
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10100 9472 11161 9500
rect 10100 9460 10106 9472
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 14056 9472 14105 9500
rect 14056 9460 14062 9472
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14734 9500 14740 9512
rect 14695 9472 14740 9500
rect 14093 9463 14151 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15010 9500 15016 9512
rect 14971 9472 15016 9500
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15120 9500 15148 9540
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17862 9568 17868 9580
rect 16908 9540 17868 9568
rect 16908 9528 16914 9540
rect 17862 9528 17868 9540
rect 17920 9568 17926 9580
rect 18049 9571 18107 9577
rect 18049 9568 18061 9571
rect 17920 9540 18061 9568
rect 17920 9528 17926 9540
rect 18049 9537 18061 9540
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 17957 9503 18015 9509
rect 15120 9472 17540 9500
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12299 9404 12909 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 12897 9401 12909 9404
rect 12943 9401 12955 9435
rect 15280 9435 15338 9441
rect 12897 9395 12955 9401
rect 14292 9404 15240 9432
rect 12342 9364 12348 9376
rect 12303 9336 12348 9364
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 14292 9373 14320 9404
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 13044 9336 13461 9364
rect 13044 9324 13050 9336
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 14277 9367 14335 9373
rect 14277 9333 14289 9367
rect 14323 9333 14335 9367
rect 14277 9327 14335 9333
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 14553 9367 14611 9373
rect 14553 9364 14565 9367
rect 14424 9336 14565 9364
rect 14424 9324 14430 9336
rect 14553 9333 14565 9336
rect 14599 9333 14611 9367
rect 15212 9364 15240 9404
rect 15280 9401 15292 9435
rect 15326 9432 15338 9435
rect 15930 9432 15936 9444
rect 15326 9404 15936 9432
rect 15326 9401 15338 9404
rect 15280 9395 15338 9401
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 16298 9364 16304 9376
rect 15212 9336 16304 9364
rect 14553 9327 14611 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 17512 9373 17540 9472
rect 17957 9469 17969 9503
rect 18003 9500 18015 9503
rect 18800 9500 18828 9664
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 19812 9540 20729 9568
rect 18003 9472 18828 9500
rect 18003 9469 18015 9472
rect 17957 9463 18015 9469
rect 18874 9460 18880 9512
rect 18932 9460 18938 9512
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 19622 9503 19680 9509
rect 19622 9500 19634 9503
rect 19392 9472 19634 9500
rect 19392 9460 19398 9472
rect 19622 9469 19634 9472
rect 19668 9500 19680 9503
rect 19812 9500 19840 9540
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 19668 9472 19840 9500
rect 19889 9503 19947 9509
rect 19668 9469 19680 9472
rect 19622 9463 19680 9469
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 20070 9500 20076 9512
rect 19935 9472 20076 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 20622 9460 20628 9512
rect 20680 9500 20686 9512
rect 21361 9503 21419 9509
rect 21361 9500 21373 9503
rect 20680 9472 21373 9500
rect 20680 9460 20686 9472
rect 21361 9469 21373 9472
rect 21407 9469 21419 9503
rect 21361 9463 21419 9469
rect 17865 9435 17923 9441
rect 17865 9401 17877 9435
rect 17911 9432 17923 9435
rect 18138 9432 18144 9444
rect 17911 9404 18144 9432
rect 17911 9401 17923 9404
rect 17865 9395 17923 9401
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18892 9432 18920 9460
rect 18892 9404 20668 9432
rect 17497 9367 17555 9373
rect 17497 9333 17509 9367
rect 17543 9333 17555 9367
rect 17497 9327 17555 9333
rect 18509 9367 18567 9373
rect 18509 9333 18521 9367
rect 18555 9364 18567 9367
rect 18874 9364 18880 9376
rect 18555 9336 18880 9364
rect 18555 9333 18567 9336
rect 18509 9327 18567 9333
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 20640 9373 20668 9404
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 20312 9336 20545 9364
rect 20312 9324 20318 9336
rect 20533 9333 20545 9336
rect 20579 9333 20591 9367
rect 20533 9327 20591 9333
rect 20625 9367 20683 9373
rect 20625 9333 20637 9367
rect 20671 9333 20683 9367
rect 20625 9327 20683 9333
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21177 9367 21235 9373
rect 21177 9364 21189 9367
rect 21140 9336 21189 9364
rect 21140 9324 21146 9336
rect 21177 9333 21189 9336
rect 21223 9333 21235 9367
rect 21177 9327 21235 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 9824 9132 10057 9160
rect 9824 9120 9830 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9129 11759 9163
rect 15930 9160 15936 9172
rect 15891 9132 15936 9160
rect 11701 9123 11759 9129
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 11716 9092 11744 9123
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16117 9163 16175 9169
rect 16117 9129 16129 9163
rect 16163 9160 16175 9163
rect 16758 9160 16764 9172
rect 16163 9132 16764 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 16758 9120 16764 9132
rect 16816 9120 16822 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 17865 9163 17923 9169
rect 17865 9160 17877 9163
rect 17644 9132 17877 9160
rect 17644 9120 17650 9132
rect 17865 9129 17877 9132
rect 17911 9129 17923 9163
rect 17865 9123 17923 9129
rect 12250 9101 12256 9104
rect 12244 9092 12256 9101
rect 8720 9064 11652 9092
rect 11716 9064 12256 9092
rect 8720 9052 8726 9064
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10588 9027 10646 9033
rect 10588 8993 10600 9027
rect 10634 9024 10646 9027
rect 10962 9024 10968 9036
rect 10634 8996 10968 9024
rect 10634 8993 10646 8996
rect 10588 8987 10646 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11624 9024 11652 9064
rect 12244 9055 12256 9064
rect 12250 9052 12256 9055
rect 12308 9052 12314 9104
rect 12406 9064 16344 9092
rect 12406 9024 12434 9064
rect 11624 8996 12434 9024
rect 14090 8984 14096 9036
rect 14148 9024 14154 9036
rect 14809 9027 14867 9033
rect 14809 9024 14821 9027
rect 14148 8996 14821 9024
rect 14148 8984 14154 8996
rect 14809 8993 14821 8996
rect 14855 8993 14867 9027
rect 14809 8987 14867 8993
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 16117 9027 16175 9033
rect 16117 9024 16129 9027
rect 15252 8996 16129 9024
rect 15252 8984 15258 8996
rect 16117 8993 16129 8996
rect 16163 9024 16175 9027
rect 16209 9027 16267 9033
rect 16209 9024 16221 9027
rect 16163 8996 16221 9024
rect 16163 8993 16175 8996
rect 16117 8987 16175 8993
rect 16209 8993 16221 8996
rect 16255 8993 16267 9027
rect 16316 9024 16344 9064
rect 16390 9052 16396 9104
rect 16448 9101 16454 9104
rect 16448 9095 16512 9101
rect 16448 9061 16466 9095
rect 16500 9061 16512 9095
rect 16448 9055 16512 9061
rect 18785 9095 18843 9101
rect 18785 9061 18797 9095
rect 18831 9092 18843 9095
rect 18966 9092 18972 9104
rect 18831 9064 18972 9092
rect 18831 9061 18843 9064
rect 18785 9055 18843 9061
rect 16448 9052 16454 9055
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 19334 9052 19340 9104
rect 19392 9092 19398 9104
rect 20070 9092 20076 9104
rect 19392 9064 20076 9092
rect 19392 9052 19398 9064
rect 20070 9052 20076 9064
rect 20128 9092 20134 9104
rect 20128 9064 21404 9092
rect 20128 9052 20134 9064
rect 18690 9024 18696 9036
rect 16316 8996 17540 9024
rect 18651 8996 18696 9024
rect 16209 8987 16267 8993
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 8168 8928 9413 8956
rect 8168 8916 8174 8928
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9582 8956 9588 8968
rect 9543 8928 9588 8956
rect 9401 8919 9459 8925
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10336 8820 10364 8919
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 11756 8928 11989 8956
rect 11756 8916 11762 8928
rect 11977 8925 11989 8928
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 14001 8959 14059 8965
rect 14001 8925 14013 8959
rect 14047 8956 14059 8959
rect 14458 8956 14464 8968
rect 14047 8928 14464 8956
rect 14047 8925 14059 8928
rect 14001 8919 14059 8925
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 11716 8820 11744 8916
rect 13354 8820 13360 8832
rect 9824 8792 11744 8820
rect 13315 8792 13360 8820
rect 9824 8780 9830 8792
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 14568 8820 14596 8919
rect 17512 8888 17540 8996
rect 18690 8984 18696 8996
rect 18748 8984 18754 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 18800 8996 19625 9024
rect 17770 8916 17776 8968
rect 17828 8956 17834 8968
rect 18800 8956 18828 8996
rect 19613 8993 19625 8996
rect 19659 9024 19671 9027
rect 20254 9024 20260 9036
rect 19659 8996 20260 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 20254 8984 20260 8996
rect 20312 9024 20318 9036
rect 20622 9024 20628 9036
rect 20312 8996 20628 9024
rect 20312 8984 20318 8996
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 21376 9033 21404 9064
rect 21094 9027 21152 9033
rect 21094 9024 21106 9027
rect 20772 8996 21106 9024
rect 20772 8984 20778 8996
rect 21094 8993 21106 8996
rect 21140 8993 21152 9027
rect 21094 8987 21152 8993
rect 21361 9027 21419 9033
rect 21361 8993 21373 9027
rect 21407 8993 21419 9027
rect 21361 8987 21419 8993
rect 18966 8956 18972 8968
rect 17828 8928 18828 8956
rect 18927 8928 18972 8956
rect 17828 8916 17834 8928
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 19981 8891 20039 8897
rect 19981 8888 19993 8891
rect 17512 8860 19993 8888
rect 19981 8857 19993 8860
rect 20027 8888 20039 8891
rect 20070 8888 20076 8900
rect 20027 8860 20076 8888
rect 20027 8857 20039 8860
rect 19981 8851 20039 8857
rect 20070 8848 20076 8860
rect 20128 8848 20134 8900
rect 15194 8820 15200 8832
rect 14568 8792 15200 8820
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 17586 8820 17592 8832
rect 17547 8792 17592 8820
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18509 8823 18567 8829
rect 18509 8820 18521 8823
rect 18104 8792 18521 8820
rect 18104 8780 18110 8792
rect 18509 8789 18521 8792
rect 18555 8789 18567 8823
rect 18509 8783 18567 8789
rect 18598 8780 18604 8832
rect 18656 8820 18662 8832
rect 18785 8823 18843 8829
rect 18785 8820 18797 8823
rect 18656 8792 18797 8820
rect 18656 8780 18662 8792
rect 18785 8789 18797 8792
rect 18831 8789 18843 8823
rect 18785 8783 18843 8789
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 8110 8616 8116 8628
rect 8071 8588 8116 8616
rect 8110 8576 8116 8588
rect 8168 8616 8174 8628
rect 8168 8588 9812 8616
rect 8168 8576 8174 8588
rect 9784 8480 9812 8588
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 11020 8588 11161 8616
rect 11020 8576 11026 8588
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 11149 8579 11207 8585
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 14792 8588 17448 8616
rect 14792 8576 14798 8588
rect 16577 8551 16635 8557
rect 16577 8517 16589 8551
rect 16623 8548 16635 8551
rect 17310 8548 17316 8560
rect 16623 8520 17316 8548
rect 16623 8517 16635 8520
rect 16577 8511 16635 8517
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 17420 8548 17448 8588
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 17736 8588 17877 8616
rect 17736 8576 17742 8588
rect 17865 8585 17877 8588
rect 17911 8585 17923 8619
rect 20714 8616 20720 8628
rect 20675 8588 20720 8616
rect 17865 8579 17923 8585
rect 20714 8576 20720 8588
rect 20772 8576 20778 8628
rect 18325 8551 18383 8557
rect 18325 8548 18337 8551
rect 17420 8520 18337 8548
rect 18325 8517 18337 8520
rect 18371 8517 18383 8551
rect 18325 8511 18383 8517
rect 9784 8452 9904 8480
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9766 8412 9772 8424
rect 9539 8384 9772 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9876 8412 9904 8452
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 16816 8452 17233 8480
rect 16816 8440 16822 8452
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 18874 8480 18880 8492
rect 18835 8452 18880 8480
rect 17221 8443 17279 8449
rect 18874 8440 18880 8452
rect 18932 8480 18938 8492
rect 18932 8452 19472 8480
rect 18932 8440 18938 8452
rect 10025 8415 10083 8421
rect 10025 8412 10037 8415
rect 9876 8384 10037 8412
rect 10025 8381 10037 8384
rect 10071 8381 10083 8415
rect 10025 8375 10083 8381
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12066 8412 12072 8424
rect 11940 8384 12072 8412
rect 11940 8372 11946 8384
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12710 8412 12716 8424
rect 12671 8384 12716 8412
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 12980 8415 13038 8421
rect 12980 8381 12992 8415
rect 13026 8412 13038 8415
rect 13354 8412 13360 8424
rect 13026 8384 13360 8412
rect 13026 8381 13038 8384
rect 12980 8375 13038 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 15194 8372 15200 8424
rect 15252 8412 15258 8424
rect 16393 8415 16451 8421
rect 16393 8412 16405 8415
rect 15252 8384 16405 8412
rect 15252 8372 15258 8384
rect 16393 8381 16405 8384
rect 16439 8381 16451 8415
rect 16393 8375 16451 8381
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8412 18751 8415
rect 18966 8412 18972 8424
rect 18739 8384 18972 8412
rect 18739 8381 18751 8384
rect 18693 8375 18751 8381
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19334 8412 19340 8424
rect 19295 8384 19340 8412
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 19444 8412 19472 8452
rect 19593 8415 19651 8421
rect 19593 8412 19605 8415
rect 19444 8384 19605 8412
rect 19593 8381 19605 8384
rect 19639 8381 19651 8415
rect 19593 8375 19651 8381
rect 9214 8344 9220 8356
rect 9272 8353 9278 8356
rect 9184 8316 9220 8344
rect 9214 8304 9220 8316
rect 9272 8307 9284 8353
rect 9272 8304 9278 8307
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 10192 8316 14381 8344
rect 10192 8304 10198 8316
rect 14369 8313 14381 8316
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 16117 8347 16175 8353
rect 16117 8313 16129 8347
rect 16163 8344 16175 8347
rect 17126 8344 17132 8356
rect 16163 8316 17132 8344
rect 16163 8313 16175 8316
rect 16117 8307 16175 8313
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17497 8347 17555 8353
rect 17497 8313 17509 8347
rect 17543 8344 17555 8347
rect 18138 8344 18144 8356
rect 17543 8316 18144 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 18785 8347 18843 8353
rect 18785 8313 18797 8347
rect 18831 8344 18843 8347
rect 20162 8344 20168 8356
rect 18831 8316 20168 8344
rect 18831 8313 18843 8316
rect 18785 8307 18843 8313
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 20254 8304 20260 8356
rect 20312 8344 20318 8356
rect 20993 8347 21051 8353
rect 20993 8344 21005 8347
rect 20312 8316 21005 8344
rect 20312 8304 20318 8316
rect 20993 8313 21005 8316
rect 21039 8313 21051 8347
rect 20993 8307 21051 8313
rect 12066 8276 12072 8288
rect 12027 8248 12072 8276
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 12434 8276 12440 8288
rect 12395 8248 12440 8276
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 14090 8276 14096 8288
rect 14051 8248 14096 8276
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 8662 8072 8668 8084
rect 8623 8044 8668 8072
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9674 8072 9680 8084
rect 9539 8044 9680 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 9784 8044 10885 8072
rect 8478 7964 8484 8016
rect 8536 8004 8542 8016
rect 9784 8004 9812 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 12342 8072 12348 8084
rect 11287 8044 12348 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 14001 8075 14059 8081
rect 14001 8041 14013 8075
rect 14047 8072 14059 8075
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14047 8044 15025 8072
rect 14047 8041 14059 8044
rect 14001 8035 14059 8041
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 16114 8032 16120 8084
rect 16172 8072 16178 8084
rect 16301 8075 16359 8081
rect 16301 8072 16313 8075
rect 16172 8044 16313 8072
rect 16172 8032 16178 8044
rect 16301 8041 16313 8044
rect 16347 8041 16359 8075
rect 16301 8035 16359 8041
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 20809 8075 20867 8081
rect 20809 8072 20821 8075
rect 16448 8044 20821 8072
rect 16448 8032 16454 8044
rect 20809 8041 20821 8044
rect 20855 8041 20867 8075
rect 20809 8035 20867 8041
rect 10962 8004 10968 8016
rect 8536 7976 9812 8004
rect 10704 7976 10968 8004
rect 8536 7964 8542 7976
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10192 7908 10241 7936
rect 10192 7896 10198 7908
rect 10229 7905 10241 7908
rect 10275 7905 10287 7939
rect 10229 7899 10287 7905
rect 10704 7877 10732 7976
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 11716 7976 12388 8004
rect 11716 7948 11744 7976
rect 12360 7948 12388 7976
rect 14458 7964 14464 8016
rect 14516 8004 14522 8016
rect 14921 8007 14979 8013
rect 14921 8004 14933 8007
rect 14516 7976 14933 8004
rect 14516 7964 14522 7976
rect 14921 7973 14933 7976
rect 14967 7973 14979 8007
rect 14921 7967 14979 7973
rect 15746 7964 15752 8016
rect 15804 8004 15810 8016
rect 15933 8007 15991 8013
rect 15933 8004 15945 8007
rect 15804 7976 15945 8004
rect 15804 7964 15810 7976
rect 15933 7973 15945 7976
rect 15979 7973 15991 8007
rect 15933 7967 15991 7973
rect 17586 7964 17592 8016
rect 17644 8004 17650 8016
rect 17690 8007 17748 8013
rect 17690 8004 17702 8007
rect 17644 7976 17702 8004
rect 17644 7964 17650 7976
rect 17690 7973 17702 7976
rect 17736 7973 17748 8007
rect 17690 7967 17748 7973
rect 17788 7976 18920 8004
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7936 11667 7939
rect 11698 7936 11704 7948
rect 11655 7908 11704 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 11876 7939 11934 7945
rect 11876 7905 11888 7939
rect 11922 7936 11934 7939
rect 12158 7936 12164 7948
rect 11922 7908 12164 7936
rect 11922 7905 11934 7908
rect 11876 7899 11934 7905
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12342 7896 12348 7948
rect 12400 7896 12406 7948
rect 13630 7936 13636 7948
rect 13591 7908 13636 7936
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15838 7936 15844 7948
rect 15712 7908 15844 7936
rect 15712 7896 15718 7908
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 17788 7936 17816 7976
rect 16040 7908 17816 7936
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 10870 7868 10876 7880
rect 10827 7840 10876 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14148 7840 15117 7868
rect 14148 7828 14154 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 14550 7800 14556 7812
rect 14511 7772 14556 7800
rect 14550 7760 14556 7772
rect 14608 7760 14614 7812
rect 15764 7800 15792 7831
rect 15930 7800 15936 7812
rect 15764 7772 15936 7800
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 10042 7732 10048 7744
rect 10003 7704 10048 7732
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12952 7704 13001 7732
rect 12952 7692 12958 7704
rect 12989 7701 13001 7704
rect 13035 7732 13047 7735
rect 16040 7732 16068 7908
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 17957 7939 18015 7945
rect 17957 7936 17969 7939
rect 17920 7908 17969 7936
rect 17920 7896 17926 7908
rect 17957 7905 17969 7908
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 18141 7939 18199 7945
rect 18141 7905 18153 7939
rect 18187 7936 18199 7939
rect 18230 7936 18236 7948
rect 18187 7908 18236 7936
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 18601 7939 18659 7945
rect 18601 7936 18613 7939
rect 18564 7908 18613 7936
rect 18564 7896 18570 7908
rect 18601 7905 18613 7908
rect 18647 7905 18659 7939
rect 18601 7899 18659 7905
rect 18693 7871 18751 7877
rect 18064 7840 18644 7868
rect 13035 7704 16068 7732
rect 16577 7735 16635 7741
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 16577 7701 16589 7735
rect 16623 7732 16635 7735
rect 16758 7732 16764 7744
rect 16623 7704 16764 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 16942 7692 16948 7744
rect 17000 7732 17006 7744
rect 18064 7732 18092 7840
rect 18506 7760 18512 7812
rect 18564 7760 18570 7812
rect 18616 7800 18644 7840
rect 18693 7837 18705 7871
rect 18739 7868 18751 7871
rect 18782 7868 18788 7880
rect 18739 7840 18788 7868
rect 18739 7837 18751 7840
rect 18693 7831 18751 7837
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 18892 7877 18920 7976
rect 20622 7964 20628 8016
rect 20680 8004 20686 8016
rect 20717 8007 20775 8013
rect 20717 8004 20729 8007
rect 20680 7976 20729 8004
rect 20680 7964 20686 7976
rect 20717 7973 20729 7976
rect 20763 7973 20775 8007
rect 20717 7967 20775 7973
rect 19978 7896 19984 7948
rect 20036 7936 20042 7948
rect 20073 7939 20131 7945
rect 20073 7936 20085 7939
rect 20036 7908 20085 7936
rect 20036 7896 20042 7908
rect 20073 7905 20085 7908
rect 20119 7905 20131 7939
rect 20073 7899 20131 7905
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7837 18935 7871
rect 18877 7831 18935 7837
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 18616 7772 19901 7800
rect 19889 7769 19901 7772
rect 19935 7769 19947 7803
rect 19889 7763 19947 7769
rect 20714 7760 20720 7812
rect 20772 7800 20778 7812
rect 20916 7800 20944 7831
rect 20772 7772 20944 7800
rect 20772 7760 20778 7772
rect 17000 7704 18092 7732
rect 18141 7735 18199 7741
rect 17000 7692 17006 7704
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18233 7735 18291 7741
rect 18233 7732 18245 7735
rect 18187 7704 18245 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18233 7701 18245 7704
rect 18279 7701 18291 7735
rect 18524 7732 18552 7760
rect 18782 7732 18788 7744
rect 18524 7704 18788 7732
rect 18233 7695 18291 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 20070 7692 20076 7744
rect 20128 7732 20134 7744
rect 20349 7735 20407 7741
rect 20349 7732 20361 7735
rect 20128 7704 20361 7732
rect 20128 7692 20134 7704
rect 20349 7701 20361 7704
rect 20395 7701 20407 7735
rect 20349 7695 20407 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 9490 7528 9496 7540
rect 9451 7500 9496 7528
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 11146 7528 11152 7540
rect 9907 7500 11152 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 11974 7528 11980 7540
rect 11931 7500 11980 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 12710 7528 12716 7540
rect 12400 7500 12716 7528
rect 12400 7488 12406 7500
rect 12710 7488 12716 7500
rect 12768 7528 12774 7540
rect 16482 7528 16488 7540
rect 12768 7500 14688 7528
rect 16443 7500 16488 7528
rect 12768 7488 12774 7500
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 10367 7432 13676 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9398 7392 9404 7404
rect 8987 7364 9404 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 10686 7392 10692 7404
rect 10647 7364 10692 7392
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 12158 7352 12164 7404
rect 12216 7392 12222 7404
rect 12437 7395 12495 7401
rect 12437 7392 12449 7395
rect 12216 7364 12449 7392
rect 12216 7352 12222 7364
rect 12437 7361 12449 7364
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 8527 7296 10149 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 10137 7293 10149 7296
rect 10183 7324 10195 7327
rect 11425 7327 11483 7333
rect 11425 7324 11437 7327
rect 10183 7296 11437 7324
rect 10183 7293 10195 7296
rect 10137 7287 10195 7293
rect 11425 7293 11437 7296
rect 11471 7293 11483 7327
rect 11425 7287 11483 7293
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12253 7327 12311 7333
rect 12253 7324 12265 7327
rect 12124 7296 12265 7324
rect 12124 7284 12130 7296
rect 12253 7293 12265 7296
rect 12299 7293 12311 7327
rect 13648 7324 13676 7432
rect 14660 7401 14688 7500
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 17402 7488 17408 7540
rect 17460 7528 17466 7540
rect 17865 7531 17923 7537
rect 17865 7528 17877 7531
rect 17460 7500 17877 7528
rect 17460 7488 17466 7500
rect 17865 7497 17877 7500
rect 17911 7497 17923 7531
rect 17865 7491 17923 7497
rect 19337 7531 19395 7537
rect 19337 7497 19349 7531
rect 19383 7528 19395 7531
rect 19886 7528 19892 7540
rect 19383 7500 19892 7528
rect 19383 7497 19395 7500
rect 19337 7491 19395 7497
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 21269 7531 21327 7537
rect 21269 7528 21281 7531
rect 20772 7500 21281 7528
rect 20772 7488 20778 7500
rect 21269 7497 21281 7500
rect 21315 7497 21327 7531
rect 21269 7491 21327 7497
rect 15105 7463 15163 7469
rect 15105 7429 15117 7463
rect 15151 7460 15163 7463
rect 18506 7460 18512 7472
rect 15151 7432 18512 7460
rect 15151 7429 15163 7432
rect 15105 7423 15163 7429
rect 18506 7420 18512 7432
rect 18564 7420 18570 7472
rect 19518 7420 19524 7472
rect 19576 7460 19582 7472
rect 19613 7463 19671 7469
rect 19613 7460 19625 7463
rect 19576 7432 19625 7460
rect 19576 7420 19582 7432
rect 19613 7429 19625 7432
rect 19659 7429 19671 7463
rect 19613 7423 19671 7429
rect 14638 7395 14696 7401
rect 14638 7361 14650 7395
rect 14684 7361 14696 7395
rect 15933 7395 15991 7401
rect 14638 7355 14696 7361
rect 14752 7364 15056 7392
rect 14752 7324 14780 7364
rect 13648 7296 14780 7324
rect 12253 7287 12311 7293
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 14884 7296 14933 7324
rect 14884 7284 14890 7296
rect 14921 7293 14933 7296
rect 14967 7293 14979 7327
rect 15028 7324 15056 7364
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 16574 7392 16580 7404
rect 15979 7364 16580 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7392 17371 7395
rect 17586 7392 17592 7404
rect 17359 7364 17592 7392
rect 17359 7361 17371 7364
rect 17313 7355 17371 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 18138 7392 18144 7404
rect 18099 7364 18144 7392
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7392 18843 7395
rect 20070 7392 20076 7404
rect 18831 7364 19840 7392
rect 20031 7364 20076 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 19812 7336 19840 7364
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20220 7364 20265 7392
rect 20220 7352 20226 7364
rect 19242 7324 19248 7336
rect 15028 7296 19248 7324
rect 14921 7287 14979 7293
rect 19242 7284 19248 7296
rect 19300 7284 19306 7336
rect 19794 7284 19800 7336
rect 19852 7284 19858 7336
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7324 20039 7327
rect 20254 7324 20260 7336
rect 20027 7296 20260 7324
rect 20027 7293 20039 7296
rect 19981 7287 20039 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 20993 7327 21051 7333
rect 20993 7293 21005 7327
rect 21039 7293 21051 7327
rect 20993 7287 21051 7293
rect 10226 7216 10232 7268
rect 10284 7256 10290 7268
rect 10965 7259 11023 7265
rect 10965 7256 10977 7259
rect 10284 7228 10977 7256
rect 10284 7216 10290 7228
rect 10965 7225 10977 7228
rect 11011 7225 11023 7259
rect 12345 7259 12403 7265
rect 12345 7256 12357 7259
rect 10965 7219 11023 7225
rect 11348 7228 12357 7256
rect 9030 7188 9036 7200
rect 8991 7160 9036 7188
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 10870 7188 10876 7200
rect 9180 7160 9225 7188
rect 10831 7160 10876 7188
rect 9180 7148 9186 7160
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 11348 7197 11376 7228
rect 12345 7225 12357 7228
rect 12391 7225 12403 7259
rect 12345 7219 12403 7225
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12989 7259 13047 7265
rect 12989 7256 13001 7259
rect 12676 7228 13001 7256
rect 12676 7216 12682 7228
rect 12989 7225 13001 7228
rect 13035 7256 13047 7259
rect 13538 7256 13544 7268
rect 13035 7228 13544 7256
rect 13035 7225 13047 7228
rect 12989 7219 13047 7225
rect 13538 7216 13544 7228
rect 13596 7216 13602 7268
rect 14400 7259 14458 7265
rect 14400 7225 14412 7259
rect 14446 7256 14458 7259
rect 16758 7256 16764 7268
rect 14446 7228 16764 7256
rect 14446 7225 14458 7228
rect 14400 7219 14458 7225
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 18138 7256 18144 7268
rect 16868 7228 18144 7256
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 11425 7191 11483 7197
rect 11425 7157 11437 7191
rect 11471 7188 11483 7191
rect 12802 7188 12808 7200
rect 11471 7160 12808 7188
rect 11471 7157 11483 7160
rect 11425 7151 11483 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13078 7148 13084 7200
rect 13136 7188 13142 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 13136 7160 13277 7188
rect 13136 7148 13142 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 15381 7191 15439 7197
rect 15381 7188 15393 7191
rect 14608 7160 15393 7188
rect 14608 7148 14614 7160
rect 15381 7157 15393 7160
rect 15427 7188 15439 7191
rect 15654 7188 15660 7200
rect 15427 7160 15660 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15896 7160 16037 7188
rect 15896 7148 15902 7160
rect 16025 7157 16037 7160
rect 16071 7157 16083 7191
rect 16025 7151 16083 7157
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 16172 7160 16217 7188
rect 16172 7148 16178 7160
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 16868 7188 16896 7228
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 21008 7256 21036 7287
rect 19208 7228 21036 7256
rect 19208 7216 19214 7228
rect 16356 7160 16896 7188
rect 16356 7148 16362 7160
rect 17034 7148 17040 7200
rect 17092 7188 17098 7200
rect 17402 7188 17408 7200
rect 17092 7160 17408 7188
rect 17092 7148 17098 7160
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17494 7148 17500 7200
rect 17552 7188 17558 7200
rect 18874 7188 18880 7200
rect 17552 7160 17597 7188
rect 18835 7160 18880 7188
rect 17552 7148 17558 7160
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 18969 7191 19027 7197
rect 18969 7157 18981 7191
rect 19015 7188 19027 7191
rect 19242 7188 19248 7200
rect 19015 7160 19248 7188
rect 19015 7157 19027 7160
rect 18969 7151 19027 7157
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 20806 7188 20812 7200
rect 20767 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 8757 6987 8815 6993
rect 8757 6953 8769 6987
rect 8803 6984 8815 6987
rect 9122 6984 9128 6996
rect 8803 6956 9128 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 10686 6984 10692 6996
rect 9232 6956 9812 6984
rect 10647 6956 10692 6984
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 9232 6916 9260 6956
rect 9784 6916 9812 6956
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12216 6956 12357 6984
rect 12216 6944 12222 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12345 6947 12403 6953
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 17954 6984 17960 6996
rect 12860 6956 17960 6984
rect 12860 6944 12866 6956
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 17494 6916 17500 6928
rect 5224 6888 9260 6916
rect 9324 6888 9720 6916
rect 9784 6888 17500 6916
rect 5224 6876 5230 6888
rect 9324 6857 9352 6888
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 9565 6851 9623 6857
rect 9565 6848 9577 6851
rect 9456 6820 9577 6848
rect 9456 6808 9462 6820
rect 9565 6817 9577 6820
rect 9611 6817 9623 6851
rect 9692 6848 9720 6888
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 17586 6876 17592 6928
rect 17644 6916 17650 6928
rect 17644 6888 19334 6916
rect 17644 6876 17650 6888
rect 9692 6820 10640 6848
rect 9565 6811 9623 6817
rect 10612 6780 10640 6820
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 11221 6851 11279 6857
rect 11221 6848 11233 6851
rect 10744 6820 11233 6848
rect 10744 6808 10750 6820
rect 11221 6817 11233 6820
rect 11267 6817 11279 6851
rect 12618 6848 12624 6860
rect 12579 6820 12624 6848
rect 11221 6811 11279 6817
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 14829 6851 14887 6857
rect 14829 6848 14841 6851
rect 14332 6820 14841 6848
rect 14332 6808 14338 6820
rect 14829 6817 14841 6820
rect 14875 6817 14887 6851
rect 14829 6811 14887 6817
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15545 6851 15603 6857
rect 15545 6848 15557 6851
rect 15436 6820 15557 6848
rect 15436 6808 15442 6820
rect 15545 6817 15557 6820
rect 15591 6817 15603 6851
rect 15545 6811 15603 6817
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16758 6848 16764 6860
rect 16080 6820 16764 6848
rect 16080 6808 16086 6820
rect 16758 6808 16764 6820
rect 16816 6848 16822 6860
rect 17862 6848 17868 6860
rect 16816 6820 17540 6848
rect 17775 6820 17868 6848
rect 16816 6808 16822 6820
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10612 6752 10977 6780
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 13170 6780 13176 6792
rect 13131 6752 13176 6780
rect 10965 6743 11023 6749
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6644 7987 6647
rect 8202 6644 8208 6656
rect 7975 6616 8208 6644
rect 7975 6613 7987 6616
rect 7929 6607 7987 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 9490 6644 9496 6656
rect 8343 6616 9496 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 10980 6644 11008 6743
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 13354 6780 13360 6792
rect 13315 6752 13360 6780
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 14734 6780 14740 6792
rect 13648 6752 14740 6780
rect 12805 6715 12863 6721
rect 12805 6681 12817 6715
rect 12851 6712 12863 6715
rect 13648 6712 13676 6752
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 15286 6780 15292 6792
rect 15247 6752 15292 6780
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 17512 6789 17540 6820
rect 17497 6783 17555 6789
rect 16356 6752 17080 6780
rect 16356 6740 16362 6752
rect 13814 6712 13820 6724
rect 12851 6684 13676 6712
rect 13775 6684 13820 6712
rect 12851 6681 12863 6684
rect 12805 6675 12863 6681
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 16574 6672 16580 6724
rect 16632 6712 16638 6724
rect 17052 6721 17080 6752
rect 17497 6749 17509 6783
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 16632 6684 16681 6712
rect 16632 6672 16638 6684
rect 16669 6681 16681 6684
rect 16715 6681 16727 6715
rect 16669 6675 16727 6681
rect 17037 6715 17095 6721
rect 17037 6681 17049 6715
rect 17083 6681 17095 6715
rect 17037 6675 17095 6681
rect 17126 6672 17132 6724
rect 17184 6712 17190 6724
rect 17788 6712 17816 6820
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 18138 6857 18144 6860
rect 18132 6811 18144 6857
rect 18196 6848 18202 6860
rect 19306 6848 19334 6888
rect 19518 6848 19524 6860
rect 18196 6820 18232 6848
rect 19306 6820 19524 6848
rect 18138 6808 18144 6811
rect 18196 6808 18202 6820
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 19794 6808 19800 6860
rect 19852 6848 19858 6860
rect 20145 6851 20203 6857
rect 20145 6848 20157 6851
rect 19852 6820 20157 6848
rect 19852 6808 19858 6820
rect 20145 6817 20157 6820
rect 20191 6817 20203 6851
rect 20145 6811 20203 6817
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 17184 6684 17816 6712
rect 17184 6672 17190 6684
rect 12342 6644 12348 6656
rect 10980 6616 12348 6644
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 14550 6644 14556 6656
rect 12492 6616 14556 6644
rect 12492 6604 12498 6616
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6644 15071 6647
rect 16298 6644 16304 6656
rect 15059 6616 16304 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 17788 6644 17816 6684
rect 19076 6752 19901 6780
rect 19076 6644 19104 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 17788 6616 19104 6644
rect 19245 6647 19303 6653
rect 19245 6613 19257 6647
rect 19291 6644 19303 6647
rect 19334 6644 19340 6656
rect 19291 6616 19340 6644
rect 19291 6613 19303 6616
rect 19245 6607 19303 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 21266 6644 21272 6656
rect 21227 6616 21272 6644
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 9456 6412 10425 6440
rect 9456 6400 9462 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11698 6440 11704 6452
rect 11379 6412 11704 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 13446 6440 13452 6452
rect 13407 6412 13452 6440
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 13955 6412 14565 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 14645 6443 14703 6449
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 15378 6440 15384 6452
rect 14691 6412 15384 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 18138 6400 18144 6452
rect 18196 6440 18202 6452
rect 18509 6443 18567 6449
rect 18509 6440 18521 6443
rect 18196 6412 18521 6440
rect 18196 6400 18202 6412
rect 18509 6409 18521 6412
rect 18555 6440 18567 6443
rect 18555 6412 19748 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 12437 6375 12495 6381
rect 12437 6341 12449 6375
rect 12483 6372 12495 6375
rect 14734 6372 14740 6384
rect 12483 6344 14740 6372
rect 12483 6341 12495 6344
rect 12437 6335 12495 6341
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 19720 6372 19748 6412
rect 19794 6400 19800 6452
rect 19852 6440 19858 6452
rect 20165 6443 20223 6449
rect 20165 6440 20177 6443
rect 19852 6412 20177 6440
rect 19852 6400 19858 6412
rect 20165 6409 20177 6412
rect 20211 6409 20223 6443
rect 20165 6403 20223 6409
rect 20622 6372 20628 6384
rect 19720 6344 20628 6372
rect 20622 6332 20628 6344
rect 20680 6372 20686 6384
rect 20680 6344 21036 6372
rect 20680 6332 20686 6344
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 12805 6307 12863 6313
rect 12805 6304 12817 6307
rect 12676 6276 12817 6304
rect 12676 6264 12682 6276
rect 12805 6273 12817 6276
rect 12851 6304 12863 6307
rect 13078 6304 13084 6316
rect 12851 6276 13084 6304
rect 12851 6273 12863 6276
rect 12805 6267 12863 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 21008 6313 21036 6344
rect 20993 6307 21051 6313
rect 16632 6276 17264 6304
rect 16632 6264 16638 6276
rect 7377 6239 7435 6245
rect 7377 6205 7389 6239
rect 7423 6236 7435 6239
rect 8662 6236 8668 6248
rect 7423 6208 8668 6236
rect 7423 6205 7435 6208
rect 7377 6199 7435 6205
rect 8662 6196 8668 6208
rect 8720 6236 8726 6248
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8720 6208 9045 6236
rect 8720 6196 8726 6208
rect 9033 6205 9045 6208
rect 9079 6205 9091 6239
rect 10686 6236 10692 6248
rect 10647 6208 10692 6236
rect 9033 6199 9091 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 11146 6236 11152 6248
rect 11107 6208 11152 6236
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 11698 6196 11704 6248
rect 11756 6236 11762 6248
rect 12253 6239 12311 6245
rect 12253 6236 12265 6239
rect 11756 6208 12265 6236
rect 11756 6196 11762 6208
rect 12253 6205 12265 6208
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 12434 6196 12440 6248
rect 12492 6196 12498 6248
rect 13722 6236 13728 6248
rect 13683 6208 13728 6236
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 13998 6196 14004 6248
rect 14056 6236 14062 6248
rect 14366 6236 14372 6248
rect 14056 6208 14228 6236
rect 14327 6208 14372 6236
rect 14056 6196 14062 6208
rect 7650 6177 7656 6180
rect 7644 6168 7656 6177
rect 7611 6140 7656 6168
rect 7644 6131 7656 6140
rect 7650 6128 7656 6131
rect 7708 6128 7714 6180
rect 9278 6171 9336 6177
rect 9278 6168 9290 6171
rect 8772 6140 9290 6168
rect 8772 6112 8800 6140
rect 9278 6137 9290 6140
rect 9324 6137 9336 6171
rect 9278 6131 9336 6137
rect 9766 6128 9772 6180
rect 9824 6168 9830 6180
rect 12452 6168 12480 6196
rect 9824 6140 12480 6168
rect 13081 6171 13139 6177
rect 9824 6128 9830 6140
rect 13081 6137 13093 6171
rect 13127 6168 13139 6171
rect 14090 6168 14096 6180
rect 13127 6140 14096 6168
rect 13127 6137 13139 6140
rect 13081 6131 13139 6137
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 14200 6168 14228 6208
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 15286 6196 15292 6248
rect 15344 6236 15350 6248
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15344 6208 16037 6236
rect 15344 6196 15350 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16390 6236 16396 6248
rect 16351 6208 16396 6236
rect 16025 6199 16083 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 17126 6236 17132 6248
rect 16540 6208 16896 6236
rect 17087 6208 17132 6236
rect 16540 6196 16546 6208
rect 15780 6171 15838 6177
rect 14200 6140 15700 6168
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 8570 6100 8576 6112
rect 7156 6072 8576 6100
rect 7156 6060 7162 6072
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 8754 6100 8760 6112
rect 8715 6072 8760 6100
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 10870 6100 10876 6112
rect 10831 6072 10876 6100
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11977 6103 12035 6109
rect 11977 6069 11989 6103
rect 12023 6100 12035 6103
rect 12066 6100 12072 6112
rect 12023 6072 12072 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12989 6103 13047 6109
rect 12989 6100 13001 6103
rect 12768 6072 13001 6100
rect 12768 6060 12774 6072
rect 12989 6069 13001 6072
rect 13035 6069 13047 6103
rect 14182 6100 14188 6112
rect 14143 6072 14188 6100
rect 12989 6063 13047 6069
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 15562 6100 15568 6112
rect 14599 6072 15568 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 15672 6100 15700 6140
rect 15780 6137 15792 6171
rect 15826 6168 15838 6171
rect 16206 6168 16212 6180
rect 15826 6140 16212 6168
rect 15826 6137 15838 6140
rect 15780 6131 15838 6137
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 16868 6168 16896 6208
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17236 6236 17264 6276
rect 20993 6273 21005 6307
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 17385 6239 17443 6245
rect 17385 6236 17397 6239
rect 17236 6208 17397 6236
rect 17385 6205 17397 6208
rect 17431 6205 17443 6239
rect 17385 6199 17443 6205
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 17920 6208 18797 6236
rect 17920 6196 17926 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 18785 6199 18843 6205
rect 19444 6208 20913 6236
rect 18690 6168 18696 6180
rect 16868 6140 18696 6168
rect 18690 6128 18696 6140
rect 18748 6128 18754 6180
rect 19052 6171 19110 6177
rect 19052 6137 19064 6171
rect 19098 6168 19110 6171
rect 19334 6168 19340 6180
rect 19098 6140 19340 6168
rect 19098 6137 19110 6140
rect 19052 6131 19110 6137
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 16482 6100 16488 6112
rect 15672 6072 16488 6100
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 16577 6103 16635 6109
rect 16577 6069 16589 6103
rect 16623 6100 16635 6103
rect 17218 6100 17224 6112
rect 16623 6072 17224 6100
rect 16623 6069 16635 6072
rect 16577 6063 16635 6069
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 17586 6060 17592 6112
rect 17644 6100 17650 6112
rect 19444 6100 19472 6208
rect 20901 6205 20913 6208
rect 20947 6205 20959 6239
rect 20901 6199 20959 6205
rect 19518 6128 19524 6180
rect 19576 6168 19582 6180
rect 20809 6171 20867 6177
rect 20809 6168 20821 6171
rect 19576 6140 20821 6168
rect 19576 6128 19582 6140
rect 20809 6137 20821 6140
rect 20855 6137 20867 6171
rect 20809 6131 20867 6137
rect 17644 6072 19472 6100
rect 17644 6060 17650 6072
rect 20162 6060 20168 6112
rect 20220 6100 20226 6112
rect 20441 6103 20499 6109
rect 20441 6100 20453 6103
rect 20220 6072 20453 6100
rect 20220 6060 20226 6072
rect 20441 6069 20453 6072
rect 20487 6069 20499 6103
rect 20441 6063 20499 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 10042 5896 10048 5908
rect 9232 5868 10048 5896
rect 9232 5828 9260 5868
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 13228 5868 13737 5896
rect 13228 5856 13234 5868
rect 13725 5865 13737 5868
rect 13771 5865 13783 5899
rect 13725 5859 13783 5865
rect 15381 5899 15439 5905
rect 15381 5865 15393 5899
rect 15427 5896 15439 5899
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15427 5868 16129 5896
rect 15427 5865 15439 5868
rect 15381 5859 15439 5865
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 16577 5899 16635 5905
rect 16577 5896 16589 5899
rect 16540 5868 16589 5896
rect 16540 5856 16546 5868
rect 16577 5865 16589 5868
rect 16623 5865 16635 5899
rect 16577 5859 16635 5865
rect 17129 5899 17187 5905
rect 17129 5865 17141 5899
rect 17175 5865 17187 5899
rect 17129 5859 17187 5865
rect 6656 5800 9260 5828
rect 9309 5831 9367 5837
rect 6656 5769 6684 5800
rect 9309 5797 9321 5831
rect 9355 5828 9367 5831
rect 10686 5828 10692 5840
rect 9355 5800 10692 5828
rect 9355 5797 9367 5800
rect 9309 5791 9367 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 11238 5837 11244 5840
rect 11180 5831 11244 5837
rect 11180 5797 11192 5831
rect 11226 5797 11244 5831
rect 11180 5791 11244 5797
rect 11238 5788 11244 5791
rect 11296 5788 11302 5840
rect 12253 5831 12311 5837
rect 12253 5797 12265 5831
rect 12299 5828 12311 5831
rect 15194 5828 15200 5840
rect 12299 5800 15200 5828
rect 12299 5797 12311 5800
rect 12253 5791 12311 5797
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 15473 5831 15531 5837
rect 15473 5797 15485 5831
rect 15519 5828 15531 5831
rect 17144 5828 17172 5859
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 18656 5868 19334 5896
rect 18656 5856 18662 5868
rect 15519 5800 17172 5828
rect 15519 5797 15531 5800
rect 15473 5791 15531 5797
rect 17678 5788 17684 5840
rect 17736 5788 17742 5840
rect 17862 5788 17868 5840
rect 17920 5828 17926 5840
rect 18785 5831 18843 5837
rect 18785 5828 18797 5831
rect 17920 5800 18797 5828
rect 17920 5788 17926 5800
rect 18785 5797 18797 5800
rect 18831 5797 18843 5831
rect 19306 5828 19334 5868
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 20533 5899 20591 5905
rect 20533 5896 20545 5899
rect 19576 5868 20545 5896
rect 19576 5856 19582 5868
rect 20533 5865 20545 5868
rect 20579 5865 20591 5899
rect 20533 5859 20591 5865
rect 21269 5831 21327 5837
rect 21269 5828 21281 5831
rect 19306 5800 21281 5828
rect 18785 5791 18843 5797
rect 21269 5797 21281 5800
rect 21315 5797 21327 5831
rect 21269 5791 21327 5797
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 7285 5763 7343 5769
rect 7285 5729 7297 5763
rect 7331 5760 7343 5763
rect 7929 5763 7987 5769
rect 7929 5760 7941 5763
rect 7331 5732 7941 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 7929 5729 7941 5732
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 8757 5763 8815 5769
rect 8757 5729 8769 5763
rect 8803 5729 8815 5763
rect 8757 5723 8815 5729
rect 7650 5692 7656 5704
rect 7611 5664 7656 5692
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5692 7895 5695
rect 8294 5692 8300 5704
rect 7883 5664 8300 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8772 5692 8800 5723
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9585 5763 9643 5769
rect 9585 5760 9597 5763
rect 9548 5732 9597 5760
rect 9548 5720 9554 5732
rect 9585 5729 9597 5732
rect 9631 5729 9643 5763
rect 9585 5723 9643 5729
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 12066 5760 12072 5772
rect 11931 5732 12072 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 12618 5769 12624 5772
rect 12612 5760 12624 5769
rect 12579 5732 12624 5760
rect 12612 5723 12624 5732
rect 12618 5720 12624 5723
rect 12676 5720 12682 5772
rect 14829 5763 14887 5769
rect 14829 5729 14841 5763
rect 14875 5760 14887 5763
rect 15562 5760 15568 5772
rect 14875 5732 15568 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 16482 5760 16488 5772
rect 16443 5732 16488 5760
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 17494 5760 17500 5772
rect 16592 5732 17500 5760
rect 10134 5692 10140 5704
rect 8772 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5692 11483 5695
rect 12342 5692 12348 5704
rect 11471 5664 12348 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15378 5692 15384 5704
rect 15335 5664 15384 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 16592 5692 16620 5732
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5760 17647 5763
rect 17696 5760 17724 5788
rect 18877 5763 18935 5769
rect 17635 5732 18828 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 15681 5664 16620 5692
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 10045 5627 10103 5633
rect 10045 5624 10057 5627
rect 8444 5596 10057 5624
rect 8444 5584 8450 5596
rect 10045 5593 10057 5596
rect 10091 5593 10103 5627
rect 10045 5587 10103 5593
rect 12069 5627 12127 5633
rect 12069 5593 12081 5627
rect 12115 5624 12127 5627
rect 12253 5627 12311 5633
rect 12253 5624 12265 5627
rect 12115 5596 12265 5624
rect 12115 5593 12127 5596
rect 12069 5587 12127 5593
rect 12253 5593 12265 5596
rect 12299 5593 12311 5627
rect 12253 5587 12311 5593
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 15681 5624 15709 5664
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 16816 5664 17693 5692
rect 16816 5652 16822 5664
rect 17681 5661 17693 5664
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5661 18751 5695
rect 18800 5692 18828 5732
rect 18877 5729 18889 5763
rect 18923 5760 18935 5763
rect 20346 5760 20352 5772
rect 18923 5732 20352 5760
rect 18923 5729 18935 5732
rect 18877 5723 18935 5729
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 20441 5763 20499 5769
rect 20441 5729 20453 5763
rect 20487 5729 20499 5763
rect 20441 5723 20499 5729
rect 20070 5692 20076 5704
rect 18800 5664 20076 5692
rect 18693 5655 18751 5661
rect 15838 5624 15844 5636
rect 14516 5596 15709 5624
rect 15799 5596 15844 5624
rect 14516 5584 14522 5596
rect 15838 5584 15844 5596
rect 15896 5584 15902 5636
rect 17034 5584 17040 5636
rect 17092 5624 17098 5636
rect 18141 5627 18199 5633
rect 18141 5624 18153 5627
rect 17092 5596 18153 5624
rect 17092 5584 17098 5596
rect 18141 5593 18153 5596
rect 18187 5593 18199 5627
rect 18708 5624 18736 5655
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 19334 5624 19340 5636
rect 18708 5596 19340 5624
rect 18141 5587 18199 5593
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 7742 5556 7748 5568
rect 6871 5528 7748 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 9766 5556 9772 5568
rect 9727 5528 9772 5556
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 17954 5556 17960 5568
rect 10744 5528 17960 5556
rect 10744 5516 10750 5528
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 18156 5556 18184 5587
rect 19334 5584 19340 5596
rect 19392 5624 19398 5636
rect 20254 5624 20260 5636
rect 19392 5596 20260 5624
rect 19392 5584 19398 5596
rect 20254 5584 20260 5596
rect 20312 5584 20318 5636
rect 18782 5556 18788 5568
rect 18156 5528 18788 5556
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 19242 5556 19248 5568
rect 19203 5528 19248 5556
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19797 5559 19855 5565
rect 19797 5525 19809 5559
rect 19843 5556 19855 5559
rect 19886 5556 19892 5568
rect 19843 5528 19892 5556
rect 19843 5525 19855 5528
rect 19797 5519 19855 5525
rect 19886 5516 19892 5528
rect 19944 5516 19950 5568
rect 20070 5556 20076 5568
rect 20031 5528 20076 5556
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 20456 5556 20484 5723
rect 20622 5692 20628 5704
rect 20583 5664 20628 5692
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 20622 5556 20628 5568
rect 20456 5528 20628 5556
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 21177 5559 21235 5565
rect 21177 5525 21189 5559
rect 21223 5556 21235 5559
rect 21358 5556 21364 5568
rect 21223 5528 21364 5556
rect 21223 5525 21235 5528
rect 21177 5519 21235 5525
rect 21358 5516 21364 5528
rect 21416 5516 21422 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 7650 5352 7656 5364
rect 6963 5324 7656 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 8662 5352 8668 5364
rect 7984 5324 8668 5352
rect 7984 5312 7990 5324
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 7282 5216 7288 5228
rect 5767 5188 7288 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 8312 5225 8340 5324
rect 8662 5312 8668 5324
rect 8720 5352 8726 5364
rect 8938 5352 8944 5364
rect 8720 5324 8944 5352
rect 8720 5312 8726 5324
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 9088 5324 9321 5352
rect 9088 5312 9094 5324
rect 9309 5321 9321 5324
rect 9355 5321 9367 5355
rect 9309 5315 9367 5321
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 9674 5352 9680 5364
rect 9456 5324 9680 5352
rect 9456 5312 9462 5324
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 9916 5324 10916 5352
rect 9916 5312 9922 5324
rect 9766 5284 9772 5296
rect 8404 5256 9772 5284
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 8404 5148 8432 5256
rect 9766 5244 9772 5256
rect 9824 5244 9830 5296
rect 10888 5284 10916 5324
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 17954 5352 17960 5364
rect 11204 5324 17960 5352
rect 11204 5312 11210 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 19613 5355 19671 5361
rect 19613 5352 19625 5355
rect 18932 5324 19625 5352
rect 18932 5312 18938 5324
rect 19613 5321 19625 5324
rect 19659 5321 19671 5355
rect 19613 5315 19671 5321
rect 19996 5324 20300 5352
rect 10888 5256 12434 5284
rect 8754 5216 8760 5228
rect 8715 5188 8760 5216
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 8996 5188 9965 5216
rect 8996 5176 9002 5188
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 5868 5120 8432 5148
rect 12406 5148 12434 5256
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 18141 5287 18199 5293
rect 18141 5284 18153 5287
rect 14792 5256 18153 5284
rect 14792 5244 14798 5256
rect 18141 5253 18153 5256
rect 18187 5253 18199 5287
rect 18141 5247 18199 5253
rect 18509 5287 18567 5293
rect 18509 5253 18521 5287
rect 18555 5284 18567 5287
rect 19996 5284 20024 5324
rect 18555 5256 20024 5284
rect 18555 5253 18567 5256
rect 18509 5247 18567 5253
rect 20070 5244 20076 5296
rect 20128 5244 20134 5296
rect 20272 5284 20300 5324
rect 20346 5312 20352 5364
rect 20404 5352 20410 5364
rect 21085 5355 21143 5361
rect 21085 5352 21097 5355
rect 20404 5324 21097 5352
rect 20404 5312 20410 5324
rect 21085 5321 21097 5324
rect 21131 5321 21143 5355
rect 21085 5315 21143 5321
rect 21542 5284 21548 5296
rect 20272 5256 21548 5284
rect 21542 5244 21548 5256
rect 21600 5244 21606 5296
rect 14090 5216 14096 5228
rect 14051 5188 14096 5216
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5216 15163 5219
rect 15930 5216 15936 5228
rect 15151 5188 15936 5216
rect 15151 5185 15163 5188
rect 15105 5179 15163 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 18601 5219 18659 5225
rect 16540 5188 18552 5216
rect 16540 5176 16546 5188
rect 13078 5148 13084 5160
rect 12406 5120 13084 5148
rect 5868 5108 5874 5120
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13170 5108 13176 5160
rect 13228 5148 13234 5160
rect 13550 5151 13608 5157
rect 13550 5148 13562 5151
rect 13228 5120 13562 5148
rect 13228 5108 13234 5120
rect 13550 5117 13562 5120
rect 13596 5117 13608 5151
rect 13550 5111 13608 5117
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5148 13875 5151
rect 13998 5148 14004 5160
rect 13863 5120 14004 5148
rect 13863 5117 13875 5120
rect 13817 5111 13875 5117
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5148 16635 5151
rect 16666 5148 16672 5160
rect 16623 5120 16672 5148
rect 16623 5117 16635 5120
rect 16577 5111 16635 5117
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 17276 5120 17325 5148
rect 17276 5108 17282 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5148 18199 5151
rect 18325 5151 18383 5157
rect 18325 5148 18337 5151
rect 18187 5120 18337 5148
rect 18187 5117 18199 5120
rect 18141 5111 18199 5117
rect 18325 5117 18337 5120
rect 18371 5117 18383 5151
rect 18524 5148 18552 5188
rect 18601 5185 18613 5219
rect 18647 5216 18659 5219
rect 19334 5216 19340 5228
rect 18647 5188 19340 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 19334 5176 19340 5188
rect 19392 5176 19398 5228
rect 18969 5151 19027 5157
rect 18524 5120 18920 5148
rect 18325 5111 18383 5117
rect 5350 5040 5356 5092
rect 5408 5080 5414 5092
rect 6089 5083 6147 5089
rect 6089 5080 6101 5083
rect 5408 5052 6101 5080
rect 5408 5040 5414 5052
rect 6089 5049 6101 5052
rect 6135 5080 6147 5083
rect 8052 5083 8110 5089
rect 6135 5052 7236 5080
rect 6135 5049 6147 5052
rect 6089 5043 6147 5049
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6914 5012 6920 5024
rect 6687 4984 6920 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 7208 5012 7236 5052
rect 8052 5049 8064 5083
rect 8098 5080 8110 5083
rect 8386 5080 8392 5092
rect 8098 5052 8392 5080
rect 8098 5049 8110 5052
rect 8052 5043 8110 5049
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 10220 5083 10278 5089
rect 8720 5052 10088 5080
rect 8720 5040 8726 5052
rect 8202 5012 8208 5024
rect 7208 4984 8208 5012
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 8941 5015 8999 5021
rect 8941 4981 8953 5015
rect 8987 5012 8999 5015
rect 9030 5012 9036 5024
rect 8987 4984 9036 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 9766 5012 9772 5024
rect 9723 4984 9772 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10060 5012 10088 5052
rect 10220 5049 10232 5083
rect 10266 5080 10278 5083
rect 10686 5080 10692 5092
rect 10266 5052 10692 5080
rect 10266 5049 10278 5052
rect 10220 5043 10278 5049
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 15194 5080 15200 5092
rect 15107 5052 15200 5080
rect 15194 5040 15200 5052
rect 15252 5080 15258 5092
rect 16482 5080 16488 5092
rect 15252 5052 16488 5080
rect 15252 5040 15258 5052
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 17773 5083 17831 5089
rect 17773 5049 17785 5083
rect 17819 5049 17831 5083
rect 17773 5043 17831 5049
rect 17957 5083 18015 5089
rect 17957 5049 17969 5083
rect 18003 5080 18015 5083
rect 18601 5083 18659 5089
rect 18601 5080 18613 5083
rect 18003 5052 18613 5080
rect 18003 5049 18015 5052
rect 17957 5043 18015 5049
rect 18601 5049 18613 5052
rect 18647 5049 18659 5083
rect 18782 5080 18788 5092
rect 18743 5052 18788 5080
rect 18601 5043 18659 5049
rect 11146 5012 11152 5024
rect 10060 4984 11152 5012
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 12032 4984 12081 5012
rect 12032 4972 12038 4984
rect 12069 4981 12081 4984
rect 12115 4981 12127 5015
rect 12069 4975 12127 4981
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12492 4984 12537 5012
rect 12492 4972 12498 4984
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 14553 5015 14611 5021
rect 14553 5012 14565 5015
rect 14516 4984 14565 5012
rect 14516 4972 14522 4984
rect 14553 4981 14565 4984
rect 14599 4981 14611 5015
rect 14553 4975 14611 4981
rect 15289 5015 15347 5021
rect 15289 4981 15301 5015
rect 15335 5012 15347 5015
rect 15378 5012 15384 5024
rect 15335 4984 15384 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 15528 4984 15669 5012
rect 15528 4972 15534 4984
rect 15657 4981 15669 4984
rect 15703 4981 15715 5015
rect 15930 5012 15936 5024
rect 15891 4984 15936 5012
rect 15657 4975 15715 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 16390 5012 16396 5024
rect 16351 4984 16396 5012
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 17221 5015 17279 5021
rect 17221 5012 17233 5015
rect 16724 4984 17233 5012
rect 16724 4972 16730 4984
rect 17221 4981 17233 4984
rect 17267 4981 17279 5015
rect 17788 5012 17816 5043
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 18892 5080 18920 5120
rect 18969 5117 18981 5151
rect 19015 5148 19027 5151
rect 19058 5148 19064 5160
rect 19015 5120 19064 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 19058 5108 19064 5120
rect 19116 5108 19122 5160
rect 19978 5148 19984 5160
rect 19939 5120 19984 5148
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 20088 5157 20116 5244
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21177 5219 21235 5225
rect 21177 5216 21189 5219
rect 21131 5188 21189 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 21177 5185 21189 5188
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5117 20131 5151
rect 20180 5148 20208 5179
rect 20254 5148 20260 5160
rect 20180 5120 20260 5148
rect 20073 5111 20131 5117
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20548 5120 20821 5148
rect 19334 5080 19340 5092
rect 18892 5052 19340 5080
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 19426 5040 19432 5092
rect 19484 5080 19490 5092
rect 20548 5080 20576 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20809 5111 20867 5117
rect 19484 5052 20576 5080
rect 20625 5083 20683 5089
rect 19484 5040 19490 5052
rect 20625 5049 20637 5083
rect 20671 5049 20683 5083
rect 20625 5043 20683 5049
rect 19794 5012 19800 5024
rect 17788 4984 19800 5012
rect 17221 4975 17279 4981
rect 19794 4972 19800 4984
rect 19852 4972 19858 5024
rect 19978 4972 19984 5024
rect 20036 5012 20042 5024
rect 20640 5012 20668 5043
rect 20036 4984 20668 5012
rect 20036 4972 20042 4984
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 5350 4808 5356 4820
rect 5311 4780 5356 4808
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 5810 4808 5816 4820
rect 5767 4780 5816 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 8294 4808 8300 4820
rect 6503 4780 8156 4808
rect 8255 4780 8300 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 7098 4672 7104 4684
rect 5031 4644 7104 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 7432 4644 7941 4672
rect 7432 4632 7438 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 8128 4672 8156 4780
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 9582 4808 9588 4820
rect 9355 4780 9588 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11425 4811 11483 4817
rect 11425 4808 11437 4811
rect 11379 4780 11437 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11425 4777 11437 4780
rect 11471 4777 11483 4811
rect 11425 4771 11483 4777
rect 11609 4811 11667 4817
rect 11609 4777 11621 4811
rect 11655 4808 11667 4811
rect 11790 4808 11796 4820
rect 11655 4780 11796 4808
rect 11655 4777 11667 4780
rect 11609 4771 11667 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 11974 4808 11980 4820
rect 11935 4780 11980 4808
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 13265 4811 13323 4817
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 13354 4808 13360 4820
rect 13311 4780 13360 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 15470 4808 15476 4820
rect 15431 4780 15476 4808
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 15933 4811 15991 4817
rect 15620 4780 15665 4808
rect 15620 4768 15626 4780
rect 15933 4777 15945 4811
rect 15979 4808 15991 4811
rect 16114 4808 16120 4820
rect 15979 4780 16120 4808
rect 15979 4777 15991 4780
rect 15933 4771 15991 4777
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 19150 4808 19156 4820
rect 18892 4780 19156 4808
rect 8846 4700 8852 4752
rect 8904 4740 8910 4752
rect 9490 4740 9496 4752
rect 8904 4712 9496 4740
rect 8904 4700 8910 4712
rect 9490 4700 9496 4712
rect 9548 4740 9554 4752
rect 9769 4743 9827 4749
rect 9769 4740 9781 4743
rect 9548 4712 9781 4740
rect 9548 4700 9554 4712
rect 9769 4709 9781 4712
rect 9815 4709 9827 4743
rect 10686 4740 10692 4752
rect 10599 4712 10692 4740
rect 9769 4703 9827 4709
rect 10686 4700 10692 4712
rect 10744 4740 10750 4752
rect 12434 4740 12440 4752
rect 10744 4712 12440 4740
rect 10744 4700 10750 4712
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 13633 4743 13691 4749
rect 13633 4709 13645 4743
rect 13679 4740 13691 4743
rect 13722 4740 13728 4752
rect 13679 4712 13728 4740
rect 13679 4709 13691 4712
rect 13633 4703 13691 4709
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 16390 4740 16396 4752
rect 16351 4712 16396 4740
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 16942 4740 16948 4752
rect 16903 4712 16948 4740
rect 16942 4700 16948 4712
rect 17000 4700 17006 4752
rect 17405 4743 17463 4749
rect 17405 4709 17417 4743
rect 17451 4740 17463 4743
rect 18690 4740 18696 4752
rect 17451 4712 18696 4740
rect 17451 4709 17463 4712
rect 17405 4703 17463 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 8573 4675 8631 4681
rect 8573 4672 8585 4675
rect 8128 4644 8585 4672
rect 7929 4635 7987 4641
rect 8573 4641 8585 4644
rect 8619 4672 8631 4675
rect 8662 4672 8668 4684
rect 8619 4644 8668 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9398 4672 9404 4684
rect 8772 4644 9404 4672
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8772 4604 8800 4644
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9674 4672 9680 4684
rect 9635 4644 9680 4672
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 7883 4576 8800 4604
rect 9953 4607 10011 4613
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 10134 4604 10140 4616
rect 9999 4576 10140 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 6089 4539 6147 4545
rect 6089 4505 6101 4539
rect 6135 4536 6147 4539
rect 7190 4536 7196 4548
rect 6135 4508 7196 4536
rect 6135 4505 6147 4508
rect 6089 4499 6147 4505
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 7760 4536 7788 4567
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10704 4613 10732 4700
rect 10962 4672 10968 4684
rect 10923 4644 10968 4672
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 11330 4632 11336 4684
rect 11388 4672 11394 4684
rect 12986 4672 12992 4684
rect 11388 4644 12204 4672
rect 12947 4644 12992 4672
rect 11388 4632 11394 4644
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4573 10747 4607
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10689 4567 10747 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 12176 4613 12204 4644
rect 12986 4632 12992 4644
rect 13044 4632 13050 4684
rect 13078 4632 13084 4684
rect 13136 4672 13142 4684
rect 14090 4672 14096 4684
rect 13136 4644 14096 4672
rect 13136 4632 13142 4644
rect 13740 4613 13768 4644
rect 14090 4632 14096 4644
rect 14148 4672 14154 4684
rect 14550 4672 14556 4684
rect 14148 4644 14556 4672
rect 14148 4632 14154 4644
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 14734 4672 14740 4684
rect 14695 4644 14740 4672
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 18805 4675 18863 4681
rect 18805 4641 18817 4675
rect 18851 4672 18863 4675
rect 18892 4672 18920 4780
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 19702 4768 19708 4820
rect 19760 4808 19766 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19760 4780 19809 4808
rect 19760 4768 19766 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 20990 4808 20996 4820
rect 19797 4771 19855 4777
rect 19904 4780 20996 4808
rect 19242 4700 19248 4752
rect 19300 4740 19306 4752
rect 19904 4740 19932 4780
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 20809 4743 20867 4749
rect 20809 4740 20821 4743
rect 19300 4712 19932 4740
rect 19996 4712 20821 4740
rect 19300 4700 19306 4712
rect 18851 4644 18920 4672
rect 18851 4641 18863 4644
rect 18805 4635 18863 4641
rect 18966 4632 18972 4684
rect 19024 4672 19030 4684
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 19024 4644 19073 4672
rect 19024 4632 19030 4644
rect 19061 4641 19073 4644
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 12069 4607 12127 4613
rect 12069 4604 12081 4607
rect 11471 4576 12081 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 12069 4573 12081 4576
rect 12115 4573 12127 4607
rect 12069 4567 12127 4573
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4573 13783 4607
rect 13725 4567 13783 4573
rect 13817 4607 13875 4613
rect 13817 4573 13829 4607
rect 13863 4573 13875 4607
rect 15286 4604 15292 4616
rect 15247 4576 15292 4604
rect 13817 4567 13875 4573
rect 8386 4536 8392 4548
rect 7760 4508 8392 4536
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 8496 4508 9674 4536
rect 6822 4468 6828 4480
rect 6783 4440 6828 4468
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 8496 4468 8524 4508
rect 7331 4440 8524 4468
rect 8757 4471 8815 4477
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 9306 4468 9312 4480
rect 8803 4440 9312 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 9646 4468 9674 4508
rect 12618 4496 12624 4548
rect 12676 4536 12682 4548
rect 13832 4536 13860 4567
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19996 4604 20024 4712
rect 20809 4709 20821 4712
rect 20855 4709 20867 4743
rect 20809 4703 20867 4709
rect 20162 4672 20168 4684
rect 20123 4644 20168 4672
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 20530 4632 20536 4684
rect 20588 4672 20594 4684
rect 20993 4675 21051 4681
rect 20993 4672 21005 4675
rect 20588 4644 21005 4672
rect 20588 4632 20594 4644
rect 20993 4641 21005 4644
rect 21039 4641 21051 4675
rect 20993 4635 21051 4641
rect 20254 4604 20260 4616
rect 19392 4576 20024 4604
rect 20215 4576 20260 4604
rect 19392 4564 19398 4576
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 20349 4607 20407 4613
rect 20349 4573 20361 4607
rect 20395 4573 20407 4607
rect 20349 4567 20407 4573
rect 12676 4508 13860 4536
rect 12676 4496 12682 4508
rect 14366 4496 14372 4548
rect 14424 4536 14430 4548
rect 14553 4539 14611 4545
rect 14553 4536 14565 4539
rect 14424 4508 14565 4536
rect 14424 4496 14430 4508
rect 14553 4505 14565 4508
rect 14599 4505 14611 4539
rect 14553 4499 14611 4505
rect 15470 4496 15476 4548
rect 15528 4536 15534 4548
rect 16209 4539 16267 4545
rect 16209 4536 16221 4539
rect 15528 4508 16221 4536
rect 15528 4496 15534 4508
rect 16209 4505 16221 4508
rect 16255 4505 16267 4539
rect 16758 4536 16764 4548
rect 16719 4508 16764 4536
rect 16209 4499 16267 4505
rect 16758 4496 16764 4508
rect 16816 4496 16822 4548
rect 17954 4536 17960 4548
rect 16868 4508 17960 4536
rect 12526 4468 12532 4480
rect 9646 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12802 4468 12808 4480
rect 12763 4440 12808 4468
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 13538 4428 13544 4480
rect 13596 4468 13602 4480
rect 16868 4468 16896 4508
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 17678 4468 17684 4480
rect 13596 4440 16896 4468
rect 17591 4440 17684 4468
rect 13596 4428 13602 4440
rect 17678 4428 17684 4440
rect 17736 4468 17742 4480
rect 20364 4468 20392 4567
rect 17736 4440 20392 4468
rect 17736 4428 17742 4440
rect 20622 4428 20628 4480
rect 20680 4468 20686 4480
rect 21266 4468 21272 4480
rect 20680 4440 21272 4468
rect 20680 4428 20686 4440
rect 21266 4428 21272 4440
rect 21324 4468 21330 4480
rect 21450 4468 21456 4480
rect 21324 4440 21456 4468
rect 21324 4428 21330 4440
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 5350 4264 5356 4276
rect 4571 4236 5356 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 6822 4224 6828 4276
rect 6880 4264 6886 4276
rect 8938 4264 8944 4276
rect 6880 4236 8944 4264
rect 6880 4224 6886 4236
rect 8938 4224 8944 4236
rect 8996 4264 9002 4276
rect 9214 4264 9220 4276
rect 8996 4236 9076 4264
rect 9175 4236 9220 4264
rect 8996 4224 9002 4236
rect 7101 4199 7159 4205
rect 7101 4165 7113 4199
rect 7147 4165 7159 4199
rect 9048 4196 9076 4236
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 14734 4224 14740 4276
rect 14792 4264 14798 4276
rect 21177 4267 21235 4273
rect 21177 4264 21189 4267
rect 14792 4236 21189 4264
rect 14792 4224 14798 4236
rect 21177 4233 21189 4236
rect 21223 4233 21235 4267
rect 21177 4227 21235 4233
rect 9490 4196 9496 4208
rect 9048 4168 9496 4196
rect 7101 4159 7159 4165
rect 7116 4128 7144 4159
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 13722 4196 13728 4208
rect 9646 4168 13728 4196
rect 9646 4128 9674 4168
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 19702 4156 19708 4208
rect 19760 4156 19766 4208
rect 20622 4156 20628 4208
rect 20680 4196 20686 4208
rect 21266 4196 21272 4208
rect 20680 4168 20760 4196
rect 20680 4156 20686 4168
rect 7116 4100 7972 4128
rect 6914 4060 6920 4072
rect 6827 4032 6920 4060
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7248 4032 7389 4060
rect 7248 4020 7254 4032
rect 7377 4029 7389 4032
rect 7423 4060 7435 4063
rect 7558 4060 7564 4072
rect 7423 4032 7564 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7708 4032 7849 4060
rect 7708 4020 7714 4032
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 7944 4060 7972 4100
rect 9416 4100 9674 4128
rect 9416 4060 9444 4100
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10100 4100 10517 4128
rect 10100 4088 10106 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 11054 4128 11060 4140
rect 10735 4100 11060 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12400 4100 12633 4128
rect 12400 4088 12406 4100
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 13872 4100 14105 4128
rect 13872 4088 13878 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4128 15991 4131
rect 16022 4128 16028 4140
rect 15979 4100 16028 4128
rect 15979 4097 15991 4100
rect 15933 4091 15991 4097
rect 16022 4088 16028 4100
rect 16080 4128 16086 4140
rect 16298 4128 16304 4140
rect 16080 4100 16304 4128
rect 16080 4088 16086 4100
rect 16298 4088 16304 4100
rect 16356 4128 16362 4140
rect 17126 4128 17132 4140
rect 16356 4100 17132 4128
rect 16356 4088 16362 4100
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 18046 4128 18052 4140
rect 17880 4100 18052 4128
rect 7944 4032 9444 4060
rect 7837 4023 7895 4029
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 9548 4032 9593 4060
rect 9548 4020 9554 4032
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9824 4032 9965 4060
rect 9824 4020 9830 4032
rect 9953 4029 9965 4032
rect 9999 4060 10011 4063
rect 10134 4060 10140 4072
rect 9999 4032 10140 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 11606 4060 11612 4072
rect 10827 4032 11612 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 11885 4063 11943 4069
rect 11885 4029 11897 4063
rect 11931 4060 11943 4063
rect 11974 4060 11980 4072
rect 11931 4032 11980 4060
rect 11931 4029 11943 4032
rect 11885 4023 11943 4029
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13780 4032 13921 4060
rect 13780 4020 13786 4032
rect 13909 4029 13921 4032
rect 13955 4060 13967 4063
rect 15194 4060 15200 4072
rect 13955 4032 15200 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 17310 4060 17316 4072
rect 17271 4032 17316 4060
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 17880 4069 17908 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 19720 4128 19748 4156
rect 20732 4137 20760 4168
rect 20824 4168 21272 4196
rect 20717 4131 20775 4137
rect 20717 4128 20729 4131
rect 19628 4100 20729 4128
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4029 17923 4063
rect 17865 4023 17923 4029
rect 18690 4020 18696 4072
rect 18748 4060 18754 4072
rect 19150 4060 19156 4072
rect 18748 4032 19156 4060
rect 18748 4020 18754 4032
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 19449 4063 19507 4069
rect 19449 4029 19461 4063
rect 19495 4060 19507 4063
rect 19628 4060 19656 4100
rect 20717 4097 20729 4100
rect 20763 4097 20775 4131
rect 20717 4091 20775 4097
rect 19495 4032 19656 4060
rect 19705 4063 19763 4069
rect 19495 4029 19507 4032
rect 19449 4023 19507 4029
rect 19705 4029 19717 4063
rect 19751 4029 19763 4063
rect 20530 4060 20536 4072
rect 20491 4032 20536 4060
rect 19705 4023 19763 4029
rect 6932 3992 6960 4020
rect 7282 3992 7288 4004
rect 6932 3964 7288 3992
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 8082 3995 8140 4001
rect 8082 3992 8094 3995
rect 7524 3964 8094 3992
rect 7524 3952 7530 3964
rect 8082 3961 8094 3964
rect 8128 3961 8140 3995
rect 10594 3992 10600 4004
rect 8082 3955 8140 3961
rect 9600 3964 10600 3992
rect 4890 3924 4896 3936
rect 4851 3896 4896 3924
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 5994 3924 6000 3936
rect 5955 3896 6000 3924
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 6730 3924 6736 3936
rect 6687 3896 6736 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7561 3927 7619 3933
rect 7561 3893 7573 3927
rect 7607 3924 7619 3927
rect 9600 3924 9628 3964
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 11698 3992 11704 4004
rect 11072 3964 11704 3992
rect 7607 3896 9628 3924
rect 9677 3927 9735 3933
rect 7607 3893 7619 3896
rect 7561 3887 7619 3893
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 10042 3924 10048 3936
rect 9723 3896 10048 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3924 10195 3927
rect 11072 3924 11100 3964
rect 11698 3952 11704 3964
rect 11756 3952 11762 4004
rect 12805 3995 12863 4001
rect 12805 3961 12817 3995
rect 12851 3992 12863 3995
rect 12851 3964 13584 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 10183 3896 11100 3924
rect 11149 3927 11207 3933
rect 10183 3893 10195 3896
rect 10137 3887 10195 3893
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11882 3924 11888 3936
rect 11195 3896 11888 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12069 3927 12127 3933
rect 12069 3893 12081 3927
rect 12115 3924 12127 3927
rect 12618 3924 12624 3936
rect 12115 3896 12624 3924
rect 12115 3893 12127 3896
rect 12069 3887 12127 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13262 3924 13268 3936
rect 12952 3896 12997 3924
rect 13223 3896 13268 3924
rect 12952 3884 12958 3896
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13556 3933 13584 3964
rect 15286 3952 15292 4004
rect 15344 3992 15350 4004
rect 15666 3995 15724 4001
rect 15666 3992 15678 3995
rect 15344 3964 15678 3992
rect 15344 3952 15350 3964
rect 15666 3961 15678 3964
rect 15712 3961 15724 3995
rect 15666 3955 15724 3961
rect 16393 3995 16451 4001
rect 16393 3961 16405 3995
rect 16439 3992 16451 3995
rect 16850 3992 16856 4004
rect 16439 3964 16856 3992
rect 16439 3961 16451 3964
rect 16393 3955 16451 3961
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 18049 3995 18107 4001
rect 18049 3961 18061 3995
rect 18095 3992 18107 3995
rect 18138 3992 18144 4004
rect 18095 3964 18144 3992
rect 18095 3961 18107 3964
rect 18049 3955 18107 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18248 3964 19196 3992
rect 13541 3927 13599 3933
rect 13541 3893 13553 3927
rect 13587 3893 13599 3927
rect 13541 3887 13599 3893
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 14090 3924 14096 3936
rect 14047 3896 14096 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14550 3924 14556 3936
rect 14511 3896 14556 3924
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 14700 3896 16313 3924
rect 14700 3884 14706 3896
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 16301 3887 16359 3893
rect 17405 3927 17463 3933
rect 17405 3893 17417 3927
rect 17451 3924 17463 3927
rect 18248 3924 18276 3964
rect 17451 3896 18276 3924
rect 18325 3927 18383 3933
rect 17451 3893 17463 3896
rect 17405 3887 17463 3893
rect 18325 3893 18337 3927
rect 18371 3924 18383 3927
rect 18598 3924 18604 3936
rect 18371 3896 18604 3924
rect 18371 3893 18383 3896
rect 18325 3887 18383 3893
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 19168 3924 19196 3964
rect 19242 3952 19248 4004
rect 19300 3992 19306 4004
rect 19720 3992 19748 4023
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20625 4063 20683 4069
rect 20625 4029 20637 4063
rect 20671 4060 20683 4063
rect 20824 4060 20852 4168
rect 21266 4156 21272 4168
rect 21324 4156 21330 4208
rect 20671 4032 20852 4060
rect 20671 4029 20683 4032
rect 20625 4023 20683 4029
rect 20898 4020 20904 4072
rect 20956 4060 20962 4072
rect 21361 4063 21419 4069
rect 21361 4060 21373 4063
rect 20956 4032 21373 4060
rect 20956 4020 20962 4032
rect 21361 4029 21373 4032
rect 21407 4029 21419 4063
rect 21361 4023 21419 4029
rect 20990 3992 20996 4004
rect 19300 3964 19748 3992
rect 19812 3964 20996 3992
rect 19300 3952 19306 3964
rect 19812 3924 19840 3964
rect 20990 3952 20996 3964
rect 21048 3952 21054 4004
rect 19168 3896 19840 3924
rect 20070 3884 20076 3936
rect 20128 3924 20134 3936
rect 20165 3927 20223 3933
rect 20165 3924 20177 3927
rect 20128 3896 20177 3924
rect 20128 3884 20134 3896
rect 20165 3893 20177 3896
rect 20211 3893 20223 3927
rect 20165 3887 20223 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 4065 3723 4123 3729
rect 4065 3689 4077 3723
rect 4111 3720 4123 3723
rect 7006 3720 7012 3732
rect 4111 3692 7012 3720
rect 4111 3689 4123 3692
rect 4065 3683 4123 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 8754 3720 8760 3732
rect 7147 3692 8760 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 11606 3720 11612 3732
rect 11567 3692 11612 3720
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11977 3723 12035 3729
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 12434 3720 12440 3732
rect 12023 3692 12440 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12434 3680 12440 3692
rect 12492 3720 12498 3732
rect 13541 3723 13599 3729
rect 13541 3720 13553 3723
rect 12492 3692 13553 3720
rect 12492 3680 12498 3692
rect 13541 3689 13553 3692
rect 13587 3689 13599 3723
rect 13541 3683 13599 3689
rect 14458 3680 14464 3732
rect 14516 3720 14522 3732
rect 14553 3723 14611 3729
rect 14553 3720 14565 3723
rect 14516 3692 14565 3720
rect 14516 3680 14522 3692
rect 14553 3689 14565 3692
rect 14599 3689 14611 3723
rect 14553 3683 14611 3689
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 16758 3720 16764 3732
rect 16080 3692 16764 3720
rect 16080 3680 16086 3692
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 19153 3723 19211 3729
rect 17604 3692 17954 3720
rect 7466 3652 7472 3664
rect 6564 3624 7472 3652
rect 6564 3525 6592 3624
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 9214 3652 9220 3664
rect 8404 3624 9220 3652
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 8404 3584 8432 3624
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 13204 3655 13262 3661
rect 10100 3624 12434 3652
rect 10100 3612 10106 3624
rect 6779 3556 8432 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 8478 3544 8484 3596
rect 8536 3593 8542 3596
rect 8536 3584 8548 3593
rect 9309 3587 9367 3593
rect 8536 3556 8581 3584
rect 8536 3547 8548 3556
rect 9309 3553 9321 3587
rect 9355 3553 9367 3587
rect 9309 3547 9367 3553
rect 8536 3544 8542 3547
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 7742 3516 7748 3528
rect 6687 3488 7748 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 8754 3516 8760 3528
rect 8715 3488 8760 3516
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 5721 3451 5779 3457
rect 5721 3417 5733 3451
rect 5767 3448 5779 3451
rect 5767 3420 7880 3448
rect 5767 3417 5779 3420
rect 5721 3411 5779 3417
rect 1210 3340 1216 3392
rect 1268 3380 1274 3392
rect 1397 3383 1455 3389
rect 1397 3380 1409 3383
rect 1268 3352 1409 3380
rect 1268 3340 1274 3352
rect 1397 3349 1409 3352
rect 1443 3349 1455 3383
rect 4338 3380 4344 3392
rect 4299 3352 4344 3380
rect 1397 3343 1455 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5074 3380 5080 3392
rect 5031 3352 5080 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3380 5411 3383
rect 5534 3380 5540 3392
rect 5399 3352 5540 3380
rect 5399 3349 5411 3352
rect 5353 3343 5411 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 6089 3383 6147 3389
rect 6089 3349 6101 3383
rect 6135 3380 6147 3383
rect 7006 3380 7012 3392
rect 6135 3352 7012 3380
rect 6135 3349 6147 3352
rect 6089 3343 6147 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7377 3383 7435 3389
rect 7377 3349 7389 3383
rect 7423 3380 7435 3383
rect 7466 3380 7472 3392
rect 7423 3352 7472 3380
rect 7423 3349 7435 3352
rect 7377 3343 7435 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7852 3380 7880 3420
rect 8846 3380 8852 3392
rect 7852 3352 8852 3380
rect 8846 3340 8852 3352
rect 8904 3380 8910 3392
rect 9324 3380 9352 3547
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 10594 3584 10600 3596
rect 9824 3556 10600 3584
rect 9824 3544 9830 3556
rect 10594 3544 10600 3556
rect 10652 3584 10658 3596
rect 11066 3587 11124 3593
rect 11066 3584 11078 3587
rect 10652 3556 11078 3584
rect 10652 3544 10658 3556
rect 11066 3553 11078 3556
rect 11112 3553 11124 3587
rect 11066 3547 11124 3553
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 11296 3556 11345 3584
rect 11296 3544 11302 3556
rect 11333 3553 11345 3556
rect 11379 3584 11391 3587
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11379 3556 11989 3584
rect 11379 3553 11391 3556
rect 11333 3547 11391 3553
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 12406 3584 12434 3624
rect 13204 3621 13216 3655
rect 13250 3652 13262 3655
rect 13814 3652 13820 3664
rect 13250 3624 13820 3652
rect 13250 3621 13262 3624
rect 13204 3615 13262 3621
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 13909 3655 13967 3661
rect 13909 3621 13921 3655
rect 13955 3652 13967 3655
rect 14182 3652 14188 3664
rect 13955 3624 14188 3652
rect 13955 3621 13967 3624
rect 13909 3615 13967 3621
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 16206 3612 16212 3664
rect 16264 3652 16270 3664
rect 17604 3652 17632 3692
rect 16264 3624 17632 3652
rect 16264 3612 16270 3624
rect 17678 3612 17684 3664
rect 17736 3661 17742 3664
rect 17736 3652 17748 3661
rect 17926 3652 17954 3692
rect 19153 3689 19165 3723
rect 19199 3720 19211 3723
rect 20162 3720 20168 3732
rect 19199 3692 20168 3720
rect 19199 3689 19211 3692
rect 19153 3683 19211 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20441 3723 20499 3729
rect 20441 3689 20453 3723
rect 20487 3720 20499 3723
rect 20714 3720 20720 3732
rect 20487 3692 20720 3720
rect 20487 3689 20499 3692
rect 20441 3683 20499 3689
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 19426 3652 19432 3664
rect 17736 3624 17781 3652
rect 17926 3624 19432 3652
rect 17736 3615 17748 3624
rect 17736 3612 17742 3615
rect 19426 3612 19432 3624
rect 19484 3612 19490 3664
rect 19886 3612 19892 3664
rect 19944 3652 19950 3664
rect 21269 3655 21327 3661
rect 21269 3652 21281 3655
rect 19944 3624 20208 3652
rect 19944 3612 19950 3624
rect 15102 3584 15108 3596
rect 12406 3556 15108 3584
rect 11977 3547 12035 3553
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 16045 3587 16103 3593
rect 16045 3553 16057 3587
rect 16091 3584 16103 3587
rect 16393 3587 16451 3593
rect 16393 3584 16405 3587
rect 16091 3556 16405 3584
rect 16091 3553 16103 3556
rect 16045 3547 16103 3553
rect 16393 3553 16405 3556
rect 16439 3553 16451 3587
rect 16393 3547 16451 3553
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 18785 3587 18843 3593
rect 16908 3556 18092 3584
rect 16908 3544 16914 3556
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3516 13507 3519
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13495 3488 13553 3516
rect 13495 3485 13507 3488
rect 13449 3479 13507 3485
rect 13541 3485 13553 3488
rect 13587 3516 13599 3519
rect 13998 3516 14004 3528
rect 13587 3488 14004 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 16298 3516 16304 3528
rect 16259 3488 16304 3516
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 9493 3451 9551 3457
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 16316 3448 16344 3476
rect 9539 3420 10456 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 9950 3380 9956 3392
rect 8904 3352 9352 3380
rect 9911 3352 9956 3380
rect 8904 3340 8910 3352
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10428 3380 10456 3420
rect 13648 3420 15424 3448
rect 16316 3420 17080 3448
rect 11882 3380 11888 3392
rect 10428 3352 11888 3380
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 12066 3380 12072 3392
rect 12027 3352 12072 3380
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12158 3340 12164 3392
rect 12216 3380 12222 3392
rect 13648 3380 13676 3420
rect 13814 3380 13820 3392
rect 12216 3352 13676 3380
rect 13775 3352 13820 3380
rect 12216 3340 12222 3352
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 14921 3383 14979 3389
rect 14921 3349 14933 3383
rect 14967 3380 14979 3383
rect 15286 3380 15292 3392
rect 14967 3352 15292 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15396 3380 15424 3420
rect 16114 3380 16120 3392
rect 15396 3352 16120 3380
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 16393 3383 16451 3389
rect 16393 3349 16405 3383
rect 16439 3380 16451 3383
rect 16574 3380 16580 3392
rect 16439 3352 16580 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 17052 3380 17080 3420
rect 17972 3380 18000 3479
rect 18064 3448 18092 3556
rect 18785 3553 18797 3587
rect 18831 3584 18843 3587
rect 20070 3584 20076 3596
rect 18831 3556 20076 3584
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 20180 3584 20208 3624
rect 20364 3624 21281 3652
rect 20364 3596 20392 3624
rect 21269 3621 21281 3624
rect 21315 3621 21327 3655
rect 21269 3615 21327 3621
rect 20346 3584 20352 3596
rect 20180 3556 20352 3584
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20806 3584 20812 3596
rect 20456 3556 20812 3584
rect 18598 3516 18604 3528
rect 18559 3488 18604 3516
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 19058 3516 19064 3528
rect 18739 3488 19064 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 20456 3516 20484 3556
rect 20806 3544 20812 3556
rect 20864 3544 20870 3596
rect 19168 3488 20484 3516
rect 19168 3448 19196 3488
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20717 3519 20775 3525
rect 20588 3488 20633 3516
rect 20588 3476 20594 3488
rect 20717 3485 20729 3519
rect 20763 3516 20775 3519
rect 21450 3516 21456 3528
rect 20763 3488 21456 3516
rect 20763 3485 20775 3488
rect 20717 3479 20775 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 18064 3420 19196 3448
rect 19797 3451 19855 3457
rect 19797 3417 19809 3451
rect 19843 3448 19855 3451
rect 21266 3448 21272 3460
rect 19843 3420 21272 3448
rect 19843 3417 19855 3420
rect 19797 3411 19855 3417
rect 21266 3408 21272 3420
rect 21324 3408 21330 3460
rect 18966 3380 18972 3392
rect 17052 3352 18972 3380
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 19886 3340 19892 3392
rect 19944 3380 19950 3392
rect 20073 3383 20131 3389
rect 20073 3380 20085 3383
rect 19944 3352 20085 3380
rect 19944 3340 19950 3352
rect 20073 3349 20085 3352
rect 20119 3349 20131 3383
rect 20073 3343 20131 3349
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 21177 3383 21235 3389
rect 21177 3380 21189 3383
rect 20496 3352 21189 3380
rect 20496 3340 20502 3352
rect 21177 3349 21189 3352
rect 21223 3349 21235 3383
rect 21177 3343 21235 3349
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 4798 3176 4804 3188
rect 4755 3148 4804 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 6086 3176 6092 3188
rect 6047 3148 6092 3176
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 7469 3179 7527 3185
rect 7469 3145 7481 3179
rect 7515 3176 7527 3179
rect 8478 3176 8484 3188
rect 7515 3148 8484 3176
rect 7515 3145 7527 3148
rect 7469 3139 7527 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10502 3176 10508 3188
rect 10100 3148 10508 3176
rect 10100 3136 10106 3148
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 12158 3176 12164 3188
rect 10928 3148 12164 3176
rect 10928 3136 10934 3148
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 13906 3176 13912 3188
rect 12483 3148 13912 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 19058 3176 19064 3188
rect 16172 3148 18828 3176
rect 19019 3148 19064 3176
rect 16172 3136 16178 3148
rect 5626 3108 5632 3120
rect 5587 3080 5632 3108
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 7193 3111 7251 3117
rect 7193 3077 7205 3111
rect 7239 3108 7251 3111
rect 7377 3111 7435 3117
rect 7377 3108 7389 3111
rect 7239 3080 7389 3108
rect 7239 3077 7251 3080
rect 7193 3071 7251 3077
rect 7377 3077 7389 3080
rect 7423 3077 7435 3111
rect 18690 3108 18696 3120
rect 7377 3071 7435 3077
rect 8864 3080 9674 3108
rect 8864 3049 8892 3080
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9214 3040 9220 3052
rect 9171 3012 9220 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 1210 2932 1216 2984
rect 1268 2972 1274 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 1268 2944 1409 2972
rect 1268 2932 1274 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 3970 2972 3976 2984
rect 3651 2944 3976 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 3970 2932 3976 2944
rect 4028 2972 4034 2984
rect 4525 2975 4583 2981
rect 4525 2972 4537 2975
rect 4028 2944 4537 2972
rect 4028 2932 4034 2944
rect 4525 2941 4537 2944
rect 4571 2941 4583 2975
rect 4525 2935 4583 2941
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 4985 2975 5043 2981
rect 4985 2972 4997 2975
rect 4948 2944 4997 2972
rect 4948 2932 4954 2944
rect 4985 2941 4997 2944
rect 5031 2941 5043 2975
rect 4985 2935 5043 2941
rect 5074 2932 5080 2984
rect 5132 2972 5138 2984
rect 5350 2972 5356 2984
rect 5132 2944 5356 2972
rect 5132 2932 5138 2944
rect 5350 2932 5356 2944
rect 5408 2972 5414 2984
rect 5445 2975 5503 2981
rect 5445 2972 5457 2975
rect 5408 2944 5457 2972
rect 5408 2932 5414 2944
rect 5445 2941 5457 2944
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 5905 2975 5963 2981
rect 5905 2972 5917 2975
rect 5776 2944 5917 2972
rect 5776 2932 5782 2944
rect 5905 2941 5917 2944
rect 5951 2941 5963 2975
rect 7006 2972 7012 2984
rect 6967 2944 7012 2972
rect 5905 2935 5963 2941
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 7282 2972 7288 2984
rect 7064 2944 7288 2972
rect 7064 2932 7070 2944
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8754 2972 8760 2984
rect 7708 2944 8760 2972
rect 7708 2932 7714 2944
rect 8754 2932 8760 2944
rect 8812 2972 8818 2984
rect 8864 2972 8892 3003
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 9646 3040 9674 3080
rect 13832 3080 18696 3108
rect 13832 3040 13860 3080
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 18800 3108 18828 3148
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 20254 3176 20260 3188
rect 20215 3148 20260 3176
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 20622 3176 20628 3188
rect 20583 3148 20628 3176
rect 20622 3136 20628 3148
rect 20680 3136 20686 3188
rect 19518 3108 19524 3120
rect 18800 3080 19524 3108
rect 19518 3068 19524 3080
rect 19576 3108 19582 3120
rect 21085 3111 21143 3117
rect 21085 3108 21097 3111
rect 19576 3080 21097 3108
rect 19576 3068 19582 3080
rect 21085 3077 21097 3080
rect 21131 3077 21143 3111
rect 21085 3071 21143 3077
rect 13998 3040 14004 3052
rect 9646 3012 10180 3040
rect 8812 2944 8892 2972
rect 8812 2932 8818 2944
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 10042 2972 10048 2984
rect 9364 2944 10048 2972
rect 9364 2932 9370 2944
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10152 2972 10180 3012
rect 13740 3012 13860 3040
rect 13924 3012 14004 3040
rect 11149 2975 11207 2981
rect 11149 2972 11161 2975
rect 10152 2944 11161 2972
rect 11149 2941 11161 2944
rect 11195 2972 11207 2975
rect 11238 2972 11244 2984
rect 11195 2944 11244 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2972 12035 2975
rect 12802 2972 12808 2984
rect 12023 2944 12808 2972
rect 12023 2941 12035 2944
rect 11977 2935 12035 2941
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 13740 2972 13768 3012
rect 13188 2944 13768 2972
rect 13817 2975 13875 2981
rect 198 2864 204 2916
rect 256 2904 262 2916
rect 1670 2904 1676 2916
rect 256 2876 1676 2904
rect 256 2864 262 2876
rect 1670 2864 1676 2876
rect 1728 2904 1734 2916
rect 1857 2907 1915 2913
rect 1857 2904 1869 2907
rect 1728 2876 1869 2904
rect 1728 2864 1734 2876
rect 1857 2873 1869 2876
rect 1903 2873 1915 2907
rect 1857 2867 1915 2873
rect 2314 2864 2320 2916
rect 2372 2904 2378 2916
rect 2961 2907 3019 2913
rect 2961 2904 2973 2907
rect 2372 2876 2973 2904
rect 2372 2864 2378 2876
rect 2961 2873 2973 2876
rect 3007 2904 3019 2907
rect 3050 2904 3056 2916
rect 3007 2876 3056 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 7377 2907 7435 2913
rect 7377 2873 7389 2907
rect 7423 2904 7435 2907
rect 8202 2904 8208 2916
rect 7423 2876 8208 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8582 2907 8640 2913
rect 8582 2873 8594 2907
rect 8628 2904 8640 2907
rect 9950 2904 9956 2916
rect 8628 2876 9956 2904
rect 8628 2873 8640 2876
rect 8582 2867 8640 2873
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 10904 2907 10962 2913
rect 10904 2873 10916 2907
rect 10950 2904 10962 2907
rect 12066 2904 12072 2916
rect 10950 2876 12072 2904
rect 10950 2873 10962 2876
rect 10904 2867 10962 2873
rect 12066 2864 12072 2876
rect 12124 2864 12130 2916
rect 12161 2907 12219 2913
rect 12161 2873 12173 2907
rect 12207 2904 12219 2907
rect 12710 2904 12716 2916
rect 12207 2876 12716 2904
rect 12207 2873 12219 2876
rect 12161 2867 12219 2873
rect 12710 2864 12716 2876
rect 12768 2864 12774 2916
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 2222 2836 2228 2848
rect 2183 2808 2228 2836
rect 2222 2796 2228 2808
rect 2280 2796 2286 2848
rect 2590 2836 2596 2848
rect 2551 2808 2596 2836
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 3878 2836 3884 2848
rect 3839 2808 3884 2836
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 6546 2836 6552 2848
rect 6507 2808 6552 2836
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 8662 2796 8668 2848
rect 8720 2836 8726 2848
rect 10042 2836 10048 2848
rect 8720 2808 10048 2836
rect 8720 2796 8726 2808
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 13188 2836 13216 2944
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 13924 2972 13952 3012
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 15286 3000 15292 3052
rect 15344 3040 15350 3052
rect 15473 3043 15531 3049
rect 15473 3040 15485 3043
rect 15344 3012 15485 3040
rect 15344 3000 15350 3012
rect 15473 3009 15485 3012
rect 15519 3040 15531 3043
rect 16298 3040 16304 3052
rect 15519 3012 16304 3040
rect 15519 3009 15531 3012
rect 15473 3003 15531 3009
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 16485 3043 16543 3049
rect 16485 3009 16497 3043
rect 16531 3040 16543 3043
rect 16574 3040 16580 3052
rect 16531 3012 16580 3040
rect 16531 3009 16543 3012
rect 16485 3003 16543 3009
rect 16574 3000 16580 3012
rect 16632 3040 16638 3052
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 16632 3012 17693 3040
rect 16632 3000 16638 3012
rect 17681 3009 17693 3012
rect 17727 3009 17739 3043
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 17681 3003 17739 3009
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 18656 3012 19625 3040
rect 18656 3000 18662 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19794 3040 19800 3052
rect 19755 3012 19800 3040
rect 19613 3003 19671 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 21358 3040 21364 3052
rect 20496 3012 21364 3040
rect 20496 3000 20502 3012
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 14550 2972 14556 2984
rect 13863 2944 13952 2972
rect 14016 2944 14556 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 13572 2907 13630 2913
rect 13572 2873 13584 2907
rect 13618 2904 13630 2907
rect 14016 2904 14044 2944
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 15930 2972 15936 2984
rect 15243 2944 15936 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 16172 2944 16344 2972
rect 16172 2932 16178 2944
rect 13618 2876 14044 2904
rect 14277 2907 14335 2913
rect 13618 2873 13630 2876
rect 13572 2867 13630 2873
rect 14277 2873 14289 2907
rect 14323 2904 14335 2907
rect 14323 2876 15056 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 10192 2808 13216 2836
rect 10192 2796 10198 2808
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 14185 2839 14243 2845
rect 14185 2836 14197 2839
rect 13320 2808 14197 2836
rect 13320 2796 13326 2808
rect 14185 2805 14197 2808
rect 14231 2805 14243 2839
rect 14185 2799 14243 2805
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14792 2808 14841 2836
rect 14792 2796 14798 2808
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 15028 2836 15056 2876
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 15289 2907 15347 2913
rect 15289 2904 15301 2907
rect 15160 2876 15301 2904
rect 15160 2864 15166 2876
rect 15289 2873 15301 2876
rect 15335 2873 15347 2907
rect 16206 2904 16212 2916
rect 16167 2876 16212 2904
rect 15289 2867 15347 2873
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 16316 2913 16344 2944
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 17460 2944 17509 2972
rect 17460 2932 17466 2944
rect 17497 2941 17509 2944
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 18414 2972 18420 2984
rect 17644 2944 18420 2972
rect 17644 2932 17650 2944
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 18693 2975 18751 2981
rect 18693 2941 18705 2975
rect 18739 2972 18751 2975
rect 19702 2972 19708 2984
rect 18739 2944 18828 2972
rect 18739 2941 18751 2944
rect 18693 2935 18751 2941
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2873 16359 2907
rect 16301 2867 16359 2873
rect 16482 2864 16488 2916
rect 16540 2904 16546 2916
rect 18601 2907 18659 2913
rect 18601 2904 18613 2907
rect 16540 2876 18613 2904
rect 16540 2864 16546 2876
rect 18601 2873 18613 2876
rect 18647 2873 18659 2907
rect 18800 2904 18828 2944
rect 19067 2944 19708 2972
rect 18966 2904 18972 2916
rect 18800 2876 18972 2904
rect 18601 2867 18659 2873
rect 18966 2864 18972 2876
rect 19024 2864 19030 2916
rect 15562 2836 15568 2848
rect 15028 2808 15568 2836
rect 14829 2799 14887 2805
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 15838 2836 15844 2848
rect 15799 2808 15844 2836
rect 15838 2796 15844 2808
rect 15896 2796 15902 2848
rect 17126 2836 17132 2848
rect 17087 2808 17132 2836
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 18506 2796 18512 2848
rect 18564 2836 18570 2848
rect 19067 2836 19095 2944
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 19886 2972 19892 2984
rect 19847 2944 19892 2972
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 22646 2972 22652 2984
rect 20680 2944 22652 2972
rect 20680 2932 20686 2944
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 19150 2864 19156 2916
rect 19208 2904 19214 2916
rect 20717 2907 20775 2913
rect 20717 2904 20729 2907
rect 19208 2876 20729 2904
rect 19208 2864 19214 2876
rect 20717 2873 20729 2876
rect 20763 2873 20775 2907
rect 21266 2904 21272 2916
rect 21227 2876 21272 2904
rect 20717 2867 20775 2873
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 18564 2808 19095 2836
rect 18564 2796 18570 2808
rect 19426 2796 19432 2848
rect 19484 2836 19490 2848
rect 20530 2836 20536 2848
rect 19484 2808 20536 2836
rect 19484 2796 19490 2808
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 7377 2635 7435 2641
rect 4755 2604 7328 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 1670 2564 1676 2576
rect 1631 2536 1676 2564
rect 1670 2524 1676 2536
rect 1728 2524 1734 2576
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2496 2191 2499
rect 2222 2496 2228 2508
rect 2179 2468 2228 2496
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2590 2496 2596 2508
rect 2551 2468 2596 2496
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 3050 2496 3056 2508
rect 3011 2468 3056 2496
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 3878 2456 3884 2508
rect 3936 2496 3942 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3936 2468 4077 2496
rect 3936 2456 3942 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4338 2456 4344 2508
rect 4396 2496 4402 2508
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 4396 2468 4537 2496
rect 4396 2456 4402 2468
rect 4525 2465 4537 2468
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 5077 2499 5135 2505
rect 5077 2465 5089 2499
rect 5123 2496 5135 2499
rect 5166 2496 5172 2508
rect 5123 2468 5172 2496
rect 5123 2465 5135 2468
rect 5077 2459 5135 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5994 2496 6000 2508
rect 5955 2468 6000 2496
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6546 2456 6552 2508
rect 6604 2496 6610 2508
rect 6733 2499 6791 2505
rect 6733 2496 6745 2499
rect 6604 2468 6745 2496
rect 6604 2456 6610 2468
rect 6733 2465 6745 2468
rect 6779 2465 6791 2499
rect 6733 2459 6791 2465
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6972 2468 7205 2496
rect 6972 2456 6978 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7300 2496 7328 2604
rect 7377 2601 7389 2635
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 7392 2564 7420 2595
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 7800 2604 7941 2632
rect 7800 2592 7806 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 7929 2595 7987 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 9398 2632 9404 2644
rect 8435 2604 9404 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 10689 2635 10747 2641
rect 9631 2604 10272 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 9674 2564 9680 2576
rect 7392 2536 9680 2564
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 9858 2524 9864 2576
rect 9916 2564 9922 2576
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9916 2536 9965 2564
rect 9916 2524 9922 2536
rect 9953 2533 9965 2536
rect 9999 2533 10011 2567
rect 10244 2564 10272 2604
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 10870 2632 10876 2644
rect 10735 2604 10876 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 11112 2604 11161 2632
rect 11112 2592 11118 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 11940 2604 12817 2632
rect 11940 2592 11946 2604
rect 12805 2601 12817 2604
rect 12851 2601 12863 2635
rect 12805 2595 12863 2601
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 12952 2604 13277 2632
rect 12952 2592 12958 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13265 2595 13323 2601
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 15105 2635 15163 2641
rect 15105 2632 15117 2635
rect 14792 2604 15117 2632
rect 14792 2592 14798 2604
rect 15105 2601 15117 2604
rect 15151 2601 15163 2635
rect 15105 2595 15163 2601
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 16209 2635 16267 2641
rect 16209 2632 16221 2635
rect 15896 2604 16221 2632
rect 15896 2592 15902 2604
rect 16209 2601 16221 2604
rect 16255 2601 16267 2635
rect 16209 2595 16267 2601
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 16540 2604 18184 2632
rect 16540 2592 16546 2604
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 10244 2536 10793 2564
rect 9953 2527 10011 2533
rect 10781 2533 10793 2536
rect 10827 2533 10839 2567
rect 10781 2527 10839 2533
rect 12618 2524 12624 2576
rect 12676 2564 12682 2576
rect 13725 2567 13783 2573
rect 13725 2564 13737 2567
rect 12676 2536 13737 2564
rect 12676 2524 12682 2536
rect 13725 2533 13737 2536
rect 13771 2533 13783 2567
rect 13725 2527 13783 2533
rect 16117 2567 16175 2573
rect 16117 2533 16129 2567
rect 16163 2564 16175 2567
rect 17126 2564 17132 2576
rect 16163 2536 17132 2564
rect 16163 2533 16175 2536
rect 16117 2527 16175 2533
rect 17126 2524 17132 2536
rect 17184 2524 17190 2576
rect 18156 2573 18184 2604
rect 18414 2592 18420 2644
rect 18472 2632 18478 2644
rect 20070 2632 20076 2644
rect 18472 2604 19288 2632
rect 20031 2604 20076 2632
rect 18472 2592 18478 2604
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2533 18199 2567
rect 18141 2527 18199 2533
rect 18598 2524 18604 2576
rect 18656 2564 18662 2576
rect 19260 2573 19288 2604
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 18785 2567 18843 2573
rect 18785 2564 18797 2567
rect 18656 2536 18797 2564
rect 18656 2524 18662 2536
rect 18785 2533 18797 2536
rect 18831 2533 18843 2567
rect 18785 2527 18843 2533
rect 19245 2567 19303 2573
rect 19245 2533 19257 2567
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 7300 2468 7788 2496
rect 7193 2459 7251 2465
rect 7374 2428 7380 2440
rect 4264 2400 7380 2428
rect 4264 2369 4292 2400
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7760 2428 7788 2468
rect 7834 2456 7840 2508
rect 7892 2496 7898 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 7892 2468 9413 2496
rect 7892 2456 7898 2468
rect 9401 2465 9413 2468
rect 9447 2496 9459 2499
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 9447 2468 11437 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 12253 2499 12311 2505
rect 12253 2465 12265 2499
rect 12299 2496 12311 2499
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12299 2468 12909 2496
rect 12299 2465 12311 2468
rect 12253 2459 12311 2465
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 16390 2456 16396 2508
rect 16448 2496 16454 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 16448 2468 17601 2496
rect 16448 2456 16454 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19116 2468 19441 2496
rect 19116 2456 19122 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 20809 2499 20867 2505
rect 20809 2496 20821 2499
rect 20772 2468 20821 2496
rect 20772 2456 20778 2468
rect 20809 2465 20821 2468
rect 20855 2465 20867 2499
rect 20809 2459 20867 2465
rect 7760 2400 8524 2428
rect 4249 2363 4307 2369
rect 4249 2329 4261 2363
rect 4295 2329 4307 2363
rect 6917 2363 6975 2369
rect 4249 2323 4307 2329
rect 4632 2332 6776 2360
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 2317 2295 2375 2301
rect 2317 2261 2329 2295
rect 2363 2292 2375 2295
rect 2498 2292 2504 2304
rect 2363 2264 2504 2292
rect 2363 2261 2375 2264
rect 2317 2255 2375 2261
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 2777 2295 2835 2301
rect 2777 2261 2789 2295
rect 2823 2292 2835 2295
rect 3142 2292 3148 2304
rect 2823 2264 3148 2292
rect 2823 2261 2835 2264
rect 2777 2255 2835 2261
rect 3142 2252 3148 2264
rect 3200 2252 3206 2304
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 4632 2292 4660 2332
rect 5258 2292 5264 2304
rect 3283 2264 4660 2292
rect 5219 2264 5264 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 5718 2292 5724 2304
rect 5679 2264 5724 2292
rect 5718 2252 5724 2264
rect 5776 2252 5782 2304
rect 6178 2292 6184 2304
rect 6139 2264 6184 2292
rect 6178 2252 6184 2264
rect 6236 2252 6242 2304
rect 6748 2292 6776 2332
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 8386 2360 8392 2372
rect 6963 2332 8392 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 8496 2360 8524 2400
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 10594 2428 10600 2440
rect 8628 2400 8673 2428
rect 10555 2400 10600 2428
rect 8628 2388 8634 2400
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 13906 2428 13912 2440
rect 12759 2400 13912 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 14550 2388 14556 2440
rect 14608 2428 14614 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14608 2400 14841 2428
rect 14608 2388 14614 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 15059 2400 15792 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 10137 2363 10195 2369
rect 8496 2332 9168 2360
rect 9030 2292 9036 2304
rect 6748 2264 9036 2292
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 9140 2292 9168 2332
rect 10137 2329 10149 2363
rect 10183 2360 10195 2363
rect 12158 2360 12164 2372
rect 10183 2332 12164 2360
rect 10183 2329 10195 2332
rect 10137 2323 10195 2329
rect 12158 2320 12164 2332
rect 12216 2320 12222 2372
rect 15764 2369 15792 2400
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16853 2431 16911 2437
rect 16356 2400 16401 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 20530 2428 20536 2440
rect 16899 2400 20536 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 13541 2363 13599 2369
rect 13541 2360 13553 2363
rect 12406 2332 13553 2360
rect 10962 2292 10968 2304
rect 9140 2264 10968 2292
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11698 2252 11704 2304
rect 11756 2292 11762 2304
rect 12406 2292 12434 2332
rect 13541 2329 13553 2332
rect 13587 2329 13599 2363
rect 13541 2323 13599 2329
rect 14185 2363 14243 2369
rect 14185 2329 14197 2363
rect 14231 2360 14243 2363
rect 15749 2363 15807 2369
rect 14231 2332 15700 2360
rect 14231 2329 14243 2332
rect 14185 2323 14243 2329
rect 11756 2264 12434 2292
rect 15473 2295 15531 2301
rect 11756 2252 11762 2264
rect 15473 2261 15485 2295
rect 15519 2292 15531 2295
rect 15562 2292 15568 2304
rect 15519 2264 15568 2292
rect 15519 2261 15531 2264
rect 15473 2255 15531 2261
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 15672 2292 15700 2332
rect 15749 2329 15761 2363
rect 15795 2329 15807 2363
rect 15749 2323 15807 2329
rect 15838 2320 15844 2372
rect 15896 2360 15902 2372
rect 16482 2360 16488 2372
rect 15896 2332 16488 2360
rect 15896 2320 15902 2332
rect 16482 2320 16488 2332
rect 16540 2320 16546 2372
rect 17126 2320 17132 2372
rect 17184 2360 17190 2372
rect 17405 2363 17463 2369
rect 17405 2360 17417 2363
rect 17184 2332 17417 2360
rect 17184 2320 17190 2332
rect 17405 2329 17417 2332
rect 17451 2329 17463 2363
rect 17405 2323 17463 2329
rect 17678 2320 17684 2372
rect 17736 2360 17742 2372
rect 17957 2363 18015 2369
rect 17957 2360 17969 2363
rect 17736 2332 17969 2360
rect 17736 2320 17742 2332
rect 17957 2329 17969 2332
rect 18003 2329 18015 2363
rect 17957 2323 18015 2329
rect 18969 2363 19027 2369
rect 18969 2329 18981 2363
rect 19015 2360 19027 2363
rect 20622 2360 20628 2372
rect 19015 2332 20628 2360
rect 19015 2329 19027 2332
rect 18969 2323 19027 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 19058 2292 19064 2304
rect 15672 2264 19064 2292
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 1762 2048 1768 2100
rect 1820 2088 1826 2100
rect 1820 2060 2774 2088
rect 1820 2048 1826 2060
rect 2746 2020 2774 2060
rect 7558 2048 7564 2100
rect 7616 2088 7622 2100
rect 9585 2091 9643 2097
rect 9585 2088 9597 2091
rect 7616 2060 9597 2088
rect 7616 2048 7622 2060
rect 9585 2057 9597 2060
rect 9631 2057 9643 2091
rect 9585 2051 9643 2057
rect 15562 2048 15568 2100
rect 15620 2088 15626 2100
rect 19610 2088 19616 2100
rect 15620 2060 19616 2088
rect 15620 2048 15626 2060
rect 19610 2048 19616 2060
rect 19668 2048 19674 2100
rect 17586 2020 17592 2032
rect 2746 1992 17592 2020
rect 17586 1980 17592 1992
rect 17644 1980 17650 2032
rect 6178 1912 6184 1964
rect 6236 1952 6242 1964
rect 18966 1952 18972 1964
rect 6236 1924 18972 1952
rect 6236 1912 6242 1924
rect 18966 1912 18972 1924
rect 19024 1912 19030 1964
rect 2498 1844 2504 1896
rect 2556 1884 2562 1896
rect 2556 1856 2774 1884
rect 2556 1844 2562 1856
rect 1762 1776 1768 1828
rect 1820 1816 1826 1828
rect 2590 1816 2596 1828
rect 1820 1788 2596 1816
rect 1820 1776 1826 1788
rect 2590 1776 2596 1788
rect 2648 1776 2654 1828
rect 658 1708 664 1760
rect 716 1748 722 1760
rect 2222 1748 2228 1760
rect 716 1720 2228 1748
rect 716 1708 722 1720
rect 2222 1708 2228 1720
rect 2280 1708 2286 1760
rect 2746 1612 2774 1856
rect 5258 1844 5264 1896
rect 5316 1884 5322 1896
rect 15378 1884 15384 1896
rect 5316 1856 15384 1884
rect 5316 1844 5322 1856
rect 15378 1844 15384 1856
rect 15436 1844 15442 1896
rect 3418 1776 3424 1828
rect 3476 1816 3482 1828
rect 4338 1816 4344 1828
rect 3476 1788 4344 1816
rect 3476 1776 3482 1788
rect 4338 1776 4344 1788
rect 4396 1776 4402 1828
rect 5994 1776 6000 1828
rect 6052 1816 6058 1828
rect 9490 1816 9496 1828
rect 6052 1788 9496 1816
rect 6052 1776 6058 1788
rect 9490 1776 9496 1788
rect 9548 1776 9554 1828
rect 9585 1819 9643 1825
rect 9585 1785 9597 1819
rect 9631 1816 9643 1819
rect 17954 1816 17960 1828
rect 9631 1788 17960 1816
rect 9631 1785 9643 1788
rect 9585 1779 9643 1785
rect 17954 1776 17960 1788
rect 18012 1776 18018 1828
rect 2866 1708 2872 1760
rect 2924 1748 2930 1760
rect 3878 1748 3884 1760
rect 2924 1720 3884 1748
rect 2924 1708 2930 1720
rect 3878 1708 3884 1720
rect 3936 1708 3942 1760
rect 5718 1708 5724 1760
rect 5776 1748 5782 1760
rect 17862 1748 17868 1760
rect 5776 1720 17868 1748
rect 5776 1708 5782 1720
rect 17862 1708 17868 1720
rect 17920 1708 17926 1760
rect 3142 1640 3148 1692
rect 3200 1680 3206 1692
rect 10226 1680 10232 1692
rect 3200 1652 10232 1680
rect 3200 1640 3206 1652
rect 10226 1640 10232 1652
rect 10284 1640 10290 1692
rect 14274 1612 14280 1624
rect 2746 1584 14280 1612
rect 14274 1572 14280 1584
rect 14332 1572 14338 1624
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 18972 20519 19024 20528
rect 18972 20485 18981 20519
rect 18981 20485 19015 20519
rect 19015 20485 19024 20519
rect 18972 20476 19024 20485
rect 19524 20519 19576 20528
rect 19524 20485 19533 20519
rect 19533 20485 19567 20519
rect 19567 20485 19576 20519
rect 19524 20476 19576 20485
rect 20628 20408 20680 20460
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 17592 20340 17644 20392
rect 18788 20315 18840 20324
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 20076 20272 20128 20324
rect 20812 20315 20864 20324
rect 5908 20247 5960 20256
rect 5908 20213 5917 20247
rect 5917 20213 5951 20247
rect 5951 20213 5960 20247
rect 5908 20204 5960 20213
rect 17408 20247 17460 20256
rect 17408 20213 17417 20247
rect 17417 20213 17451 20247
rect 17451 20213 17460 20247
rect 17408 20204 17460 20213
rect 17960 20204 18012 20256
rect 20812 20281 20821 20315
rect 20821 20281 20855 20315
rect 20855 20281 20864 20315
rect 20812 20272 20864 20281
rect 21088 20315 21140 20324
rect 21088 20281 21097 20315
rect 21097 20281 21131 20315
rect 21131 20281 21140 20315
rect 21088 20272 21140 20281
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 17224 20000 17276 20052
rect 17592 20043 17644 20052
rect 17592 20009 17601 20043
rect 17601 20009 17635 20043
rect 17635 20009 17644 20043
rect 17592 20000 17644 20009
rect 18788 20000 18840 20052
rect 18604 19932 18656 19984
rect 19708 19864 19760 19916
rect 20260 19907 20312 19916
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 20628 19907 20680 19916
rect 20628 19873 20637 19907
rect 20637 19873 20671 19907
rect 20671 19873 20680 19907
rect 20628 19864 20680 19873
rect 20812 19907 20864 19916
rect 20812 19873 20821 19907
rect 20821 19873 20855 19907
rect 20855 19873 20864 19907
rect 20812 19864 20864 19873
rect 21180 19907 21232 19916
rect 21180 19873 21189 19907
rect 21189 19873 21223 19907
rect 21223 19873 21232 19907
rect 21180 19864 21232 19873
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 19708 19499 19760 19508
rect 19708 19465 19717 19499
rect 19717 19465 19751 19499
rect 19751 19465 19760 19499
rect 19708 19456 19760 19465
rect 20076 19456 20128 19508
rect 20628 19499 20680 19508
rect 20628 19465 20637 19499
rect 20637 19465 20671 19499
rect 20671 19465 20680 19499
rect 20628 19456 20680 19465
rect 5908 19252 5960 19304
rect 11980 19252 12032 19304
rect 18696 19252 18748 19304
rect 20076 19252 20128 19304
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 7288 19184 7340 19236
rect 16764 19184 16816 19236
rect 21364 19227 21416 19236
rect 21364 19193 21373 19227
rect 21373 19193 21407 19227
rect 21407 19193 21416 19227
rect 21364 19184 21416 19193
rect 17960 19116 18012 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 11980 18955 12032 18964
rect 11980 18921 11989 18955
rect 11989 18921 12023 18955
rect 12023 18921 12032 18955
rect 11980 18912 12032 18921
rect 18696 18955 18748 18964
rect 18696 18921 18705 18955
rect 18705 18921 18739 18955
rect 18739 18921 18748 18955
rect 18696 18912 18748 18921
rect 20076 18955 20128 18964
rect 20076 18921 20085 18955
rect 20085 18921 20119 18955
rect 20119 18921 20128 18955
rect 20076 18912 20128 18921
rect 21180 18912 21232 18964
rect 11980 18776 12032 18828
rect 18604 18776 18656 18828
rect 19616 18776 19668 18828
rect 20628 18819 20680 18828
rect 20628 18785 20637 18819
rect 20637 18785 20671 18819
rect 20671 18785 20680 18819
rect 20628 18776 20680 18785
rect 21180 18819 21232 18828
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 21364 18683 21416 18692
rect 21364 18649 21373 18683
rect 21373 18649 21407 18683
rect 21407 18649 21416 18683
rect 21364 18640 21416 18649
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 20260 18368 20312 18420
rect 16764 18300 16816 18352
rect 9496 18164 9548 18216
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 19984 18164 20036 18216
rect 20812 18164 20864 18216
rect 20260 18096 20312 18148
rect 21364 18139 21416 18148
rect 21364 18105 21373 18139
rect 21373 18105 21407 18139
rect 21407 18105 21416 18139
rect 21364 18096 21416 18105
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 21180 17824 21232 17876
rect 8300 17688 8352 17740
rect 19800 17688 19852 17740
rect 20352 17620 20404 17672
rect 21364 17595 21416 17604
rect 21364 17561 21373 17595
rect 21373 17561 21407 17595
rect 21407 17561 21416 17595
rect 21364 17552 21416 17561
rect 20628 17484 20680 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 12164 17280 12216 17332
rect 19800 17323 19852 17332
rect 19800 17289 19809 17323
rect 19809 17289 19843 17323
rect 19843 17289 19852 17323
rect 19800 17280 19852 17289
rect 20260 17323 20312 17332
rect 20260 17289 20269 17323
rect 20269 17289 20303 17323
rect 20303 17289 20312 17323
rect 20260 17280 20312 17289
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 11796 17076 11848 17128
rect 13820 17076 13872 17128
rect 20076 17119 20128 17128
rect 20076 17085 20085 17119
rect 20085 17085 20119 17119
rect 20119 17085 20128 17119
rect 20076 17076 20128 17085
rect 20628 17051 20680 17060
rect 20628 17017 20637 17051
rect 20637 17017 20671 17051
rect 20671 17017 20680 17051
rect 20628 17008 20680 17017
rect 21180 17051 21232 17060
rect 21180 17017 21189 17051
rect 21189 17017 21223 17051
rect 21223 17017 21232 17051
rect 21180 17008 21232 17017
rect 21456 17008 21508 17060
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 20076 16736 20128 16788
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 20628 16779 20680 16788
rect 20628 16745 20637 16779
rect 20637 16745 20671 16779
rect 20671 16745 20680 16779
rect 20628 16736 20680 16745
rect 20260 16668 20312 16720
rect 17684 16600 17736 16652
rect 17960 16600 18012 16652
rect 20168 16643 20220 16652
rect 20168 16609 20177 16643
rect 20177 16609 20211 16643
rect 20211 16609 20220 16643
rect 20168 16600 20220 16609
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 20168 16192 20220 16244
rect 21180 16192 21232 16244
rect 16580 15988 16632 16040
rect 16028 15920 16080 15972
rect 21364 15963 21416 15972
rect 20444 15852 20496 15904
rect 21364 15929 21373 15963
rect 21373 15929 21407 15963
rect 21407 15929 21416 15963
rect 21364 15920 21416 15929
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 17960 15648 18012 15700
rect 20260 15691 20312 15700
rect 20260 15657 20269 15691
rect 20269 15657 20303 15691
rect 20303 15657 20312 15691
rect 20260 15648 20312 15657
rect 20812 15623 20864 15632
rect 20812 15589 20821 15623
rect 20821 15589 20855 15623
rect 20855 15589 20864 15623
rect 20812 15580 20864 15589
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 20628 15555 20680 15564
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 16028 15104 16080 15156
rect 20628 15147 20680 15156
rect 20628 15113 20637 15147
rect 20637 15113 20671 15147
rect 20671 15113 20680 15147
rect 20628 15104 20680 15113
rect 11888 14943 11940 14952
rect 11888 14909 11897 14943
rect 11897 14909 11931 14943
rect 11931 14909 11940 14943
rect 11888 14900 11940 14909
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 20352 14832 20404 14884
rect 21456 14832 21508 14884
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 20076 14560 20128 14612
rect 20444 14560 20496 14612
rect 21180 14560 21232 14612
rect 8852 14424 8904 14476
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 16304 14424 16356 14476
rect 21180 14467 21232 14476
rect 17960 14356 18012 14408
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 20812 14288 20864 14340
rect 21364 14331 21416 14340
rect 21364 14297 21373 14331
rect 21373 14297 21407 14331
rect 21407 14297 21416 14331
rect 21364 14288 21416 14297
rect 18880 14220 18932 14272
rect 19248 14220 19300 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 20536 14016 20588 14068
rect 16304 13948 16356 14000
rect 20996 13948 21048 14000
rect 17132 13880 17184 13932
rect 12164 13812 12216 13864
rect 17776 13812 17828 13864
rect 18696 13812 18748 13864
rect 18880 13812 18932 13864
rect 19340 13812 19392 13864
rect 20904 13812 20956 13864
rect 21548 13812 21600 13864
rect 8576 13744 8628 13796
rect 18512 13787 18564 13796
rect 18512 13753 18521 13787
rect 18521 13753 18555 13787
rect 18555 13753 18564 13787
rect 18512 13744 18564 13753
rect 19064 13676 19116 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 17960 13472 18012 13524
rect 20352 13515 20404 13524
rect 20352 13481 20361 13515
rect 20361 13481 20395 13515
rect 20395 13481 20404 13515
rect 20352 13472 20404 13481
rect 21180 13472 21232 13524
rect 17408 13404 17460 13456
rect 13268 13336 13320 13388
rect 18696 13404 18748 13456
rect 21364 13447 21416 13456
rect 21364 13413 21373 13447
rect 21373 13413 21407 13447
rect 21407 13413 21416 13447
rect 21364 13404 21416 13413
rect 18512 13336 18564 13388
rect 19064 13379 19116 13388
rect 19064 13345 19073 13379
rect 19073 13345 19107 13379
rect 19107 13345 19116 13379
rect 19064 13336 19116 13345
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 20628 13379 20680 13388
rect 20628 13345 20637 13379
rect 20637 13345 20671 13379
rect 20671 13345 20680 13379
rect 20628 13336 20680 13345
rect 17868 13200 17920 13252
rect 16028 13132 16080 13184
rect 20812 13268 20864 13320
rect 21088 13268 21140 13320
rect 19156 13200 19208 13252
rect 20260 13132 20312 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 18788 12928 18840 12980
rect 20628 12928 20680 12980
rect 21088 12928 21140 12980
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 16948 12724 17000 12776
rect 18420 12724 18472 12776
rect 18972 12724 19024 12776
rect 19156 12767 19208 12776
rect 19156 12733 19165 12767
rect 19165 12733 19199 12767
rect 19199 12733 19208 12767
rect 19156 12724 19208 12733
rect 19708 12724 19760 12776
rect 19892 12724 19944 12776
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 16856 12656 16908 12708
rect 17040 12656 17092 12708
rect 18052 12656 18104 12708
rect 18512 12631 18564 12640
rect 18512 12597 18521 12631
rect 18521 12597 18555 12631
rect 18555 12597 18564 12631
rect 18512 12588 18564 12597
rect 20628 12588 20680 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 20168 12384 20220 12436
rect 21088 12384 21140 12436
rect 14648 12248 14700 12300
rect 17960 12316 18012 12368
rect 18512 12316 18564 12368
rect 20904 12316 20956 12368
rect 15936 12291 15988 12300
rect 15936 12257 15970 12291
rect 15970 12257 15988 12291
rect 15936 12248 15988 12257
rect 16948 12248 17000 12300
rect 17316 12248 17368 12300
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 19616 12248 19668 12300
rect 20536 12291 20588 12300
rect 20536 12257 20545 12291
rect 20545 12257 20579 12291
rect 20579 12257 20588 12291
rect 20536 12248 20588 12257
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 18880 12180 18932 12232
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 15292 12087 15344 12096
rect 15292 12053 15301 12087
rect 15301 12053 15335 12087
rect 15335 12053 15344 12087
rect 15292 12044 15344 12053
rect 16948 12044 17000 12096
rect 17868 12044 17920 12096
rect 18052 12044 18104 12096
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 20352 12087 20404 12096
rect 20352 12053 20361 12087
rect 20361 12053 20395 12087
rect 20395 12053 20404 12087
rect 20352 12044 20404 12053
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 13544 11840 13596 11892
rect 18052 11840 18104 11892
rect 18604 11840 18656 11892
rect 13728 11772 13780 11824
rect 18880 11772 18932 11824
rect 15844 11704 15896 11756
rect 15292 11636 15344 11688
rect 16120 11636 16172 11688
rect 16488 11636 16540 11688
rect 17776 11704 17828 11756
rect 17960 11704 18012 11756
rect 17592 11636 17644 11688
rect 19248 11636 19300 11688
rect 20076 11679 20128 11688
rect 20076 11645 20094 11679
rect 20094 11645 20128 11679
rect 20076 11636 20128 11645
rect 20996 11679 21048 11688
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 9312 11568 9364 11620
rect 17040 11568 17092 11620
rect 8668 11500 8720 11552
rect 14004 11500 14056 11552
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 19984 11568 20036 11620
rect 20168 11568 20220 11620
rect 20996 11645 21005 11679
rect 21005 11645 21039 11679
rect 21039 11645 21048 11679
rect 20996 11636 21048 11645
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 17500 11500 17552 11552
rect 19340 11500 19392 11552
rect 20996 11500 21048 11552
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 15752 11296 15804 11348
rect 17040 11296 17092 11348
rect 17500 11339 17552 11348
rect 17500 11305 17509 11339
rect 17509 11305 17543 11339
rect 17543 11305 17552 11339
rect 17500 11296 17552 11305
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 14648 11203 14700 11212
rect 14648 11169 14657 11203
rect 14657 11169 14691 11203
rect 14691 11169 14700 11203
rect 14648 11160 14700 11169
rect 15476 11160 15528 11212
rect 16856 11160 16908 11212
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 17040 11135 17092 11144
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17408 11228 17460 11280
rect 17868 11160 17920 11212
rect 19248 11160 19300 11212
rect 19984 11160 20036 11212
rect 20720 11160 20772 11212
rect 17040 11092 17092 11101
rect 13912 11024 13964 11076
rect 15844 11024 15896 11076
rect 16304 11024 16356 11076
rect 19064 11092 19116 11144
rect 19340 11092 19392 11144
rect 19800 11092 19852 11144
rect 20076 11092 20128 11144
rect 19524 11024 19576 11076
rect 19248 10956 19300 11008
rect 20720 10956 20772 11008
rect 21272 10999 21324 11008
rect 21272 10965 21281 10999
rect 21281 10965 21315 10999
rect 21315 10965 21324 10999
rect 21272 10956 21324 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 13912 10752 13964 10804
rect 11704 10616 11756 10668
rect 15476 10752 15528 10804
rect 19524 10752 19576 10804
rect 17408 10684 17460 10736
rect 15936 10591 15988 10600
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 12900 10523 12952 10532
rect 12900 10489 12934 10523
rect 12934 10489 12952 10523
rect 12900 10480 12952 10489
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 17040 10548 17092 10600
rect 17859 10591 17911 10600
rect 17859 10557 17868 10591
rect 17868 10557 17902 10591
rect 17902 10557 17911 10591
rect 17859 10548 17911 10557
rect 18972 10548 19024 10600
rect 14648 10480 14700 10532
rect 16304 10480 16356 10532
rect 19800 10548 19852 10600
rect 16672 10412 16724 10464
rect 18696 10412 18748 10464
rect 19340 10412 19392 10464
rect 19432 10455 19484 10464
rect 19432 10421 19441 10455
rect 19441 10421 19475 10455
rect 19475 10421 19484 10455
rect 20076 10480 20128 10532
rect 19432 10412 19484 10421
rect 20904 10412 20956 10464
rect 21088 10455 21140 10464
rect 21088 10421 21097 10455
rect 21097 10421 21131 10455
rect 21131 10421 21140 10455
rect 21088 10412 21140 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 13544 10208 13596 10260
rect 13636 10208 13688 10260
rect 14648 10140 14700 10192
rect 15660 10208 15712 10260
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 18604 10208 18656 10260
rect 20076 10208 20128 10260
rect 20812 10251 20864 10260
rect 20812 10217 20821 10251
rect 20821 10217 20855 10251
rect 20855 10217 20864 10251
rect 20812 10208 20864 10217
rect 16764 10140 16816 10192
rect 17408 10140 17460 10192
rect 14188 10072 14240 10124
rect 14740 10072 14792 10124
rect 17592 10072 17644 10124
rect 14648 9936 14700 9988
rect 14280 9868 14332 9920
rect 15292 10004 15344 10056
rect 15936 10047 15988 10056
rect 15476 9936 15528 9988
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 18328 10072 18380 10124
rect 19248 10115 19300 10124
rect 19248 10081 19257 10115
rect 19257 10081 19291 10115
rect 19291 10081 19300 10115
rect 19248 10072 19300 10081
rect 19800 10072 19852 10124
rect 20720 10115 20772 10124
rect 20720 10081 20729 10115
rect 20729 10081 20763 10115
rect 20763 10081 20772 10115
rect 20720 10072 20772 10081
rect 21088 10004 21140 10056
rect 15844 9936 15896 9988
rect 17224 9936 17276 9988
rect 18788 9936 18840 9988
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 20536 9868 20588 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 13544 9664 13596 9716
rect 15292 9664 15344 9716
rect 15936 9664 15988 9716
rect 16396 9707 16448 9716
rect 16396 9673 16405 9707
rect 16405 9673 16439 9707
rect 16439 9673 16448 9707
rect 16396 9664 16448 9673
rect 18788 9664 18840 9716
rect 11704 9596 11756 9648
rect 11888 9639 11940 9648
rect 11888 9605 11897 9639
rect 11897 9605 11931 9639
rect 11931 9605 11940 9639
rect 11888 9596 11940 9605
rect 17040 9639 17092 9648
rect 17040 9605 17049 9639
rect 17049 9605 17083 9639
rect 17083 9605 17092 9639
rect 17040 9596 17092 9605
rect 17960 9596 18012 9648
rect 12256 9528 12308 9580
rect 10048 9460 10100 9512
rect 14004 9460 14056 9512
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 16856 9528 16908 9580
rect 17868 9528 17920 9580
rect 12348 9367 12400 9376
rect 12348 9333 12357 9367
rect 12357 9333 12391 9367
rect 12391 9333 12400 9367
rect 12348 9324 12400 9333
rect 12992 9324 13044 9376
rect 14372 9324 14424 9376
rect 15936 9392 15988 9444
rect 16304 9324 16356 9376
rect 18880 9460 18932 9512
rect 19340 9460 19392 9512
rect 20076 9460 20128 9512
rect 20628 9460 20680 9512
rect 18144 9392 18196 9444
rect 18880 9324 18932 9376
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 20260 9324 20312 9376
rect 21088 9324 21140 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 9772 9120 9824 9172
rect 15936 9163 15988 9172
rect 8668 9052 8720 9104
rect 15936 9129 15945 9163
rect 15945 9129 15979 9163
rect 15979 9129 15988 9163
rect 15936 9120 15988 9129
rect 16764 9120 16816 9172
rect 17592 9120 17644 9172
rect 12256 9095 12308 9104
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 10968 8984 11020 9036
rect 12256 9061 12290 9095
rect 12290 9061 12308 9095
rect 12256 9052 12308 9061
rect 14096 8984 14148 9036
rect 15200 8984 15252 9036
rect 16396 9052 16448 9104
rect 18972 9052 19024 9104
rect 19340 9052 19392 9104
rect 20076 9052 20128 9104
rect 18696 9027 18748 9036
rect 8116 8916 8168 8968
rect 9588 8959 9640 8968
rect 9588 8925 9597 8959
rect 9597 8925 9631 8959
rect 9631 8925 9640 8959
rect 9588 8916 9640 8925
rect 9772 8780 9824 8832
rect 11704 8916 11756 8968
rect 14464 8916 14516 8968
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 18696 8993 18705 9027
rect 18705 8993 18739 9027
rect 18739 8993 18748 9027
rect 18696 8984 18748 8993
rect 17776 8916 17828 8968
rect 20260 8984 20312 9036
rect 20628 8984 20680 9036
rect 20720 8984 20772 9036
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 20076 8848 20128 8900
rect 15200 8780 15252 8832
rect 17592 8823 17644 8832
rect 17592 8789 17601 8823
rect 17601 8789 17635 8823
rect 17635 8789 17644 8823
rect 17592 8780 17644 8789
rect 18052 8780 18104 8832
rect 18604 8780 18656 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 10968 8576 11020 8628
rect 14740 8576 14792 8628
rect 17316 8508 17368 8560
rect 17684 8576 17736 8628
rect 20720 8619 20772 8628
rect 20720 8585 20729 8619
rect 20729 8585 20763 8619
rect 20763 8585 20772 8619
rect 20720 8576 20772 8585
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 16764 8440 16816 8492
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 11888 8372 11940 8424
rect 12072 8372 12124 8424
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 13360 8372 13412 8424
rect 15200 8372 15252 8424
rect 18972 8372 19024 8424
rect 19340 8415 19392 8424
rect 19340 8381 19349 8415
rect 19349 8381 19383 8415
rect 19383 8381 19392 8415
rect 19340 8372 19392 8381
rect 9220 8347 9272 8356
rect 9220 8313 9238 8347
rect 9238 8313 9272 8347
rect 9220 8304 9272 8313
rect 10140 8304 10192 8356
rect 17132 8304 17184 8356
rect 18144 8304 18196 8356
rect 20168 8304 20220 8356
rect 20260 8304 20312 8356
rect 12072 8279 12124 8288
rect 12072 8245 12081 8279
rect 12081 8245 12115 8279
rect 12115 8245 12124 8279
rect 12072 8236 12124 8245
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 14096 8279 14148 8288
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 14096 8236 14148 8245
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 9680 8032 9732 8084
rect 8484 7964 8536 8016
rect 12348 8032 12400 8084
rect 16120 8032 16172 8084
rect 16396 8032 16448 8084
rect 10140 7896 10192 7948
rect 10968 7964 11020 8016
rect 14464 7964 14516 8016
rect 15752 7964 15804 8016
rect 17592 7964 17644 8016
rect 11704 7896 11756 7948
rect 12164 7896 12216 7948
rect 12348 7896 12400 7948
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 15660 7896 15712 7948
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 10876 7828 10928 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14096 7828 14148 7880
rect 14556 7803 14608 7812
rect 14556 7769 14565 7803
rect 14565 7769 14599 7803
rect 14599 7769 14608 7803
rect 14556 7760 14608 7769
rect 15936 7760 15988 7812
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 12900 7692 12952 7744
rect 17868 7896 17920 7948
rect 18236 7896 18288 7948
rect 18512 7896 18564 7948
rect 16764 7692 16816 7744
rect 16948 7692 17000 7744
rect 18512 7760 18564 7812
rect 18788 7828 18840 7880
rect 20628 7964 20680 8016
rect 19984 7896 20036 7948
rect 20720 7760 20772 7812
rect 18788 7692 18840 7744
rect 20076 7692 20128 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 9496 7531 9548 7540
rect 9496 7497 9505 7531
rect 9505 7497 9539 7531
rect 9539 7497 9548 7531
rect 9496 7488 9548 7497
rect 11152 7488 11204 7540
rect 11980 7488 12032 7540
rect 12348 7488 12400 7540
rect 12716 7488 12768 7540
rect 16488 7531 16540 7540
rect 9404 7352 9456 7404
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 12164 7352 12216 7404
rect 12072 7284 12124 7336
rect 16488 7497 16497 7531
rect 16497 7497 16531 7531
rect 16531 7497 16540 7531
rect 16488 7488 16540 7497
rect 17408 7488 17460 7540
rect 19892 7488 19944 7540
rect 20720 7488 20772 7540
rect 18512 7420 18564 7472
rect 19524 7420 19576 7472
rect 14832 7284 14884 7336
rect 16580 7352 16632 7404
rect 17592 7352 17644 7404
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 20168 7395 20220 7404
rect 20168 7361 20177 7395
rect 20177 7361 20211 7395
rect 20211 7361 20220 7395
rect 20168 7352 20220 7361
rect 19248 7284 19300 7336
rect 19800 7284 19852 7336
rect 20260 7284 20312 7336
rect 10232 7216 10284 7268
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 10876 7191 10928 7200
rect 9128 7148 9180 7157
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 12624 7216 12676 7268
rect 13544 7216 13596 7268
rect 16764 7216 16816 7268
rect 12808 7148 12860 7200
rect 13084 7148 13136 7200
rect 14556 7148 14608 7200
rect 15660 7148 15712 7200
rect 15844 7148 15896 7200
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 16304 7148 16356 7200
rect 18144 7216 18196 7268
rect 19156 7216 19208 7268
rect 17040 7148 17092 7200
rect 17408 7191 17460 7200
rect 17408 7157 17417 7191
rect 17417 7157 17451 7191
rect 17451 7157 17460 7191
rect 17408 7148 17460 7157
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 18880 7191 18932 7200
rect 17500 7148 17552 7157
rect 18880 7157 18889 7191
rect 18889 7157 18923 7191
rect 18923 7157 18932 7191
rect 18880 7148 18932 7157
rect 19248 7148 19300 7200
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 9128 6944 9180 6996
rect 10692 6987 10744 6996
rect 5172 6876 5224 6928
rect 10692 6953 10701 6987
rect 10701 6953 10735 6987
rect 10735 6953 10744 6987
rect 10692 6944 10744 6953
rect 12164 6944 12216 6996
rect 12808 6944 12860 6996
rect 17960 6944 18012 6996
rect 9404 6808 9456 6860
rect 17500 6876 17552 6928
rect 17592 6876 17644 6928
rect 10692 6808 10744 6860
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 14280 6808 14332 6860
rect 15384 6808 15436 6860
rect 16028 6808 16080 6860
rect 16764 6808 16816 6860
rect 17868 6851 17920 6860
rect 13176 6783 13228 6792
rect 8208 6604 8260 6656
rect 9496 6604 9548 6656
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 14740 6740 14792 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 16304 6740 16356 6792
rect 13820 6715 13872 6724
rect 13820 6681 13829 6715
rect 13829 6681 13863 6715
rect 13863 6681 13872 6715
rect 13820 6672 13872 6681
rect 16580 6672 16632 6724
rect 17132 6672 17184 6724
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 18144 6851 18196 6860
rect 18144 6817 18178 6851
rect 18178 6817 18196 6851
rect 18144 6808 18196 6817
rect 19524 6808 19576 6860
rect 19800 6808 19852 6860
rect 12348 6604 12400 6656
rect 12440 6604 12492 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 16304 6604 16356 6656
rect 19340 6604 19392 6656
rect 21272 6647 21324 6656
rect 21272 6613 21281 6647
rect 21281 6613 21315 6647
rect 21315 6613 21324 6647
rect 21272 6604 21324 6613
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 9404 6400 9456 6452
rect 11704 6400 11756 6452
rect 13452 6443 13504 6452
rect 13452 6409 13461 6443
rect 13461 6409 13495 6443
rect 13495 6409 13504 6443
rect 13452 6400 13504 6409
rect 15384 6400 15436 6452
rect 18144 6400 18196 6452
rect 14740 6332 14792 6384
rect 19800 6400 19852 6452
rect 20628 6332 20680 6384
rect 12624 6264 12676 6316
rect 13084 6264 13136 6316
rect 16580 6264 16632 6316
rect 8668 6196 8720 6248
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 11152 6239 11204 6248
rect 11152 6205 11161 6239
rect 11161 6205 11195 6239
rect 11195 6205 11204 6239
rect 11152 6196 11204 6205
rect 11704 6196 11756 6248
rect 12440 6196 12492 6248
rect 13728 6239 13780 6248
rect 13728 6205 13737 6239
rect 13737 6205 13771 6239
rect 13771 6205 13780 6239
rect 13728 6196 13780 6205
rect 14004 6196 14056 6248
rect 14372 6239 14424 6248
rect 7656 6171 7708 6180
rect 7656 6137 7690 6171
rect 7690 6137 7708 6171
rect 7656 6128 7708 6137
rect 9772 6128 9824 6180
rect 14096 6128 14148 6180
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 15292 6196 15344 6248
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 16488 6196 16540 6248
rect 17132 6239 17184 6248
rect 7104 6060 7156 6112
rect 8576 6060 8628 6112
rect 8760 6103 8812 6112
rect 8760 6069 8769 6103
rect 8769 6069 8803 6103
rect 8803 6069 8812 6103
rect 8760 6060 8812 6069
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 12072 6060 12124 6112
rect 12716 6060 12768 6112
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 15568 6060 15620 6112
rect 16212 6128 16264 6180
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 17868 6196 17920 6248
rect 18696 6128 18748 6180
rect 19340 6128 19392 6180
rect 16488 6060 16540 6112
rect 17224 6060 17276 6112
rect 17592 6060 17644 6112
rect 19524 6128 19576 6180
rect 20168 6060 20220 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 10048 5856 10100 5908
rect 13176 5856 13228 5908
rect 16488 5856 16540 5908
rect 10692 5788 10744 5840
rect 11244 5788 11296 5840
rect 15200 5788 15252 5840
rect 18604 5856 18656 5908
rect 17684 5788 17736 5840
rect 17868 5788 17920 5840
rect 19524 5856 19576 5908
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 8300 5652 8352 5704
rect 9496 5720 9548 5772
rect 12072 5720 12124 5772
rect 12624 5763 12676 5772
rect 12624 5729 12658 5763
rect 12658 5729 12676 5763
rect 12624 5720 12676 5729
rect 15568 5720 15620 5772
rect 16488 5763 16540 5772
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 17500 5763 17552 5772
rect 10140 5652 10192 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 15384 5652 15436 5704
rect 17500 5729 17509 5763
rect 17509 5729 17543 5763
rect 17543 5729 17552 5763
rect 17500 5720 17552 5729
rect 8392 5584 8444 5636
rect 14464 5584 14516 5636
rect 16764 5695 16816 5704
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 20352 5720 20404 5772
rect 15844 5627 15896 5636
rect 15844 5593 15853 5627
rect 15853 5593 15887 5627
rect 15887 5593 15896 5627
rect 15844 5584 15896 5593
rect 17040 5584 17092 5636
rect 20076 5652 20128 5704
rect 7748 5516 7800 5568
rect 9772 5559 9824 5568
rect 9772 5525 9781 5559
rect 9781 5525 9815 5559
rect 9815 5525 9824 5559
rect 9772 5516 9824 5525
rect 10692 5516 10744 5568
rect 17960 5516 18012 5568
rect 19340 5584 19392 5636
rect 20260 5584 20312 5636
rect 18788 5516 18840 5568
rect 19248 5559 19300 5568
rect 19248 5525 19257 5559
rect 19257 5525 19291 5559
rect 19291 5525 19300 5559
rect 19248 5516 19300 5525
rect 19892 5516 19944 5568
rect 20076 5559 20128 5568
rect 20076 5525 20085 5559
rect 20085 5525 20119 5559
rect 20119 5525 20128 5559
rect 20076 5516 20128 5525
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 20628 5516 20680 5568
rect 21364 5516 21416 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 7656 5312 7708 5364
rect 7932 5312 7984 5364
rect 7288 5176 7340 5228
rect 8668 5312 8720 5364
rect 8944 5312 8996 5364
rect 9036 5312 9088 5364
rect 9404 5312 9456 5364
rect 9680 5312 9732 5364
rect 9864 5312 9916 5364
rect 5816 5108 5868 5160
rect 9772 5244 9824 5296
rect 11152 5312 11204 5364
rect 17960 5312 18012 5364
rect 18880 5312 18932 5364
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 8944 5176 8996 5228
rect 14740 5244 14792 5296
rect 20076 5244 20128 5296
rect 20352 5312 20404 5364
rect 21548 5244 21600 5296
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 15936 5176 15988 5228
rect 16488 5176 16540 5228
rect 13084 5108 13136 5160
rect 13176 5108 13228 5160
rect 14004 5108 14056 5160
rect 16672 5108 16724 5160
rect 17224 5108 17276 5160
rect 19340 5176 19392 5228
rect 5356 5040 5408 5092
rect 6920 4972 6972 5024
rect 8392 5040 8444 5092
rect 8668 5040 8720 5092
rect 8208 4972 8260 5024
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 9036 4972 9088 5024
rect 9772 4972 9824 5024
rect 10692 5040 10744 5092
rect 15200 5083 15252 5092
rect 15200 5049 15209 5083
rect 15209 5049 15243 5083
rect 15243 5049 15252 5083
rect 15200 5040 15252 5049
rect 16488 5040 16540 5092
rect 18788 5083 18840 5092
rect 11152 4972 11204 5024
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 11980 4972 12032 5024
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 14464 4972 14516 5024
rect 15384 4972 15436 5024
rect 15476 4972 15528 5024
rect 15936 5015 15988 5024
rect 15936 4981 15945 5015
rect 15945 4981 15979 5015
rect 15979 4981 15988 5015
rect 15936 4972 15988 4981
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 16672 4972 16724 5024
rect 18788 5049 18797 5083
rect 18797 5049 18831 5083
rect 18831 5049 18840 5083
rect 18788 5040 18840 5049
rect 19064 5108 19116 5160
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 20260 5108 20312 5160
rect 19340 5040 19392 5092
rect 19432 5040 19484 5092
rect 19800 4972 19852 5024
rect 19984 4972 20036 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 5816 4768 5868 4820
rect 8300 4811 8352 4820
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7380 4632 7432 4684
rect 8300 4777 8309 4811
rect 8309 4777 8343 4811
rect 8343 4777 8352 4811
rect 8300 4768 8352 4777
rect 9588 4768 9640 4820
rect 11796 4768 11848 4820
rect 11980 4811 12032 4820
rect 11980 4777 11989 4811
rect 11989 4777 12023 4811
rect 12023 4777 12032 4811
rect 11980 4768 12032 4777
rect 13360 4768 13412 4820
rect 15476 4811 15528 4820
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 15568 4811 15620 4820
rect 15568 4777 15577 4811
rect 15577 4777 15611 4811
rect 15611 4777 15620 4811
rect 15568 4768 15620 4777
rect 16120 4768 16172 4820
rect 8852 4700 8904 4752
rect 9496 4700 9548 4752
rect 10692 4700 10744 4752
rect 12440 4700 12492 4752
rect 13728 4700 13780 4752
rect 16396 4743 16448 4752
rect 16396 4709 16405 4743
rect 16405 4709 16439 4743
rect 16439 4709 16448 4743
rect 16396 4700 16448 4709
rect 16948 4743 17000 4752
rect 16948 4709 16957 4743
rect 16957 4709 16991 4743
rect 16991 4709 17000 4743
rect 16948 4700 17000 4709
rect 18696 4700 18748 4752
rect 8668 4632 8720 4684
rect 9404 4632 9456 4684
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 7196 4496 7248 4548
rect 10140 4564 10192 4616
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 11336 4632 11388 4684
rect 12992 4675 13044 4684
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 13084 4632 13136 4684
rect 14096 4632 14148 4684
rect 14556 4632 14608 4684
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 19156 4768 19208 4820
rect 19708 4768 19760 4820
rect 19248 4700 19300 4752
rect 20996 4768 21048 4820
rect 18972 4632 19024 4684
rect 15292 4607 15344 4616
rect 8392 4496 8444 4548
rect 6828 4471 6880 4480
rect 6828 4437 6837 4471
rect 6837 4437 6871 4471
rect 6871 4437 6880 4471
rect 6828 4428 6880 4437
rect 9312 4428 9364 4480
rect 12624 4496 12676 4548
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 19340 4564 19392 4616
rect 20168 4675 20220 4684
rect 20168 4641 20177 4675
rect 20177 4641 20211 4675
rect 20211 4641 20220 4675
rect 20168 4632 20220 4641
rect 20536 4632 20588 4684
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 14372 4496 14424 4548
rect 15476 4496 15528 4548
rect 16764 4539 16816 4548
rect 16764 4505 16773 4539
rect 16773 4505 16807 4539
rect 16807 4505 16816 4539
rect 16764 4496 16816 4505
rect 12532 4428 12584 4480
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 13544 4428 13596 4480
rect 17960 4496 18012 4548
rect 17684 4471 17736 4480
rect 17684 4437 17693 4471
rect 17693 4437 17727 4471
rect 17727 4437 17736 4471
rect 17684 4428 17736 4437
rect 20628 4428 20680 4480
rect 21272 4428 21324 4480
rect 21456 4428 21508 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 5356 4224 5408 4276
rect 6828 4224 6880 4276
rect 8944 4224 8996 4276
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 14740 4224 14792 4276
rect 9496 4156 9548 4208
rect 13728 4156 13780 4208
rect 19708 4156 19760 4208
rect 20628 4156 20680 4208
rect 6920 4063 6972 4072
rect 6920 4029 6929 4063
rect 6929 4029 6963 4063
rect 6963 4029 6972 4063
rect 6920 4020 6972 4029
rect 7196 4020 7248 4072
rect 7564 4020 7616 4072
rect 7656 4020 7708 4072
rect 10048 4088 10100 4140
rect 11060 4088 11112 4140
rect 12348 4088 12400 4140
rect 13820 4088 13872 4140
rect 16028 4088 16080 4140
rect 16304 4088 16356 4140
rect 17132 4088 17184 4140
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 9772 4020 9824 4072
rect 10140 4020 10192 4072
rect 11612 4020 11664 4072
rect 11980 4020 12032 4072
rect 13728 4020 13780 4072
rect 15200 4020 15252 4072
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 18052 4088 18104 4140
rect 18696 4020 18748 4072
rect 19156 4020 19208 4072
rect 20536 4063 20588 4072
rect 7288 3952 7340 4004
rect 7472 3952 7524 4004
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 6000 3927 6052 3936
rect 6000 3893 6009 3927
rect 6009 3893 6043 3927
rect 6043 3893 6052 3927
rect 6000 3884 6052 3893
rect 6736 3884 6788 3936
rect 10600 3952 10652 4004
rect 10048 3884 10100 3936
rect 11704 3952 11756 4004
rect 11888 3884 11940 3936
rect 12624 3884 12676 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 13268 3927 13320 3936
rect 12900 3884 12952 3893
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 15292 3952 15344 4004
rect 16856 3952 16908 4004
rect 18144 3952 18196 4004
rect 14096 3884 14148 3936
rect 14556 3927 14608 3936
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 14648 3884 14700 3936
rect 18604 3884 18656 3936
rect 19248 3952 19300 4004
rect 20536 4029 20545 4063
rect 20545 4029 20579 4063
rect 20579 4029 20588 4063
rect 20536 4020 20588 4029
rect 21272 4156 21324 4208
rect 20904 4020 20956 4072
rect 20996 3952 21048 4004
rect 20076 3884 20128 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 7012 3680 7064 3732
rect 8760 3680 8812 3732
rect 11612 3723 11664 3732
rect 11612 3689 11621 3723
rect 11621 3689 11655 3723
rect 11655 3689 11664 3723
rect 11612 3680 11664 3689
rect 12440 3680 12492 3732
rect 14464 3680 14516 3732
rect 16028 3680 16080 3732
rect 16764 3680 16816 3732
rect 7472 3612 7524 3664
rect 9220 3612 9272 3664
rect 10048 3612 10100 3664
rect 8484 3587 8536 3596
rect 8484 3553 8502 3587
rect 8502 3553 8536 3587
rect 8484 3544 8536 3553
rect 7748 3476 7800 3528
rect 8760 3519 8812 3528
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 1216 3340 1268 3392
rect 4344 3383 4396 3392
rect 4344 3349 4353 3383
rect 4353 3349 4387 3383
rect 4387 3349 4396 3383
rect 4344 3340 4396 3349
rect 5080 3340 5132 3392
rect 5540 3340 5592 3392
rect 7012 3340 7064 3392
rect 7472 3340 7524 3392
rect 8852 3340 8904 3392
rect 9772 3544 9824 3596
rect 10600 3544 10652 3596
rect 11244 3544 11296 3596
rect 13820 3612 13872 3664
rect 14188 3612 14240 3664
rect 16212 3612 16264 3664
rect 17684 3655 17736 3664
rect 17684 3621 17702 3655
rect 17702 3621 17736 3655
rect 20168 3680 20220 3732
rect 20720 3680 20772 3732
rect 17684 3612 17736 3621
rect 19432 3612 19484 3664
rect 19892 3612 19944 3664
rect 15108 3544 15160 3596
rect 16856 3544 16908 3596
rect 14004 3476 14056 3528
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 11888 3340 11940 3392
rect 12072 3383 12124 3392
rect 12072 3349 12081 3383
rect 12081 3349 12115 3383
rect 12115 3349 12124 3383
rect 12072 3340 12124 3349
rect 12164 3340 12216 3392
rect 13820 3383 13872 3392
rect 13820 3349 13829 3383
rect 13829 3349 13863 3383
rect 13863 3349 13872 3383
rect 13820 3340 13872 3349
rect 15292 3340 15344 3392
rect 16120 3340 16172 3392
rect 16580 3383 16632 3392
rect 16580 3349 16589 3383
rect 16589 3349 16623 3383
rect 16623 3349 16632 3383
rect 16580 3340 16632 3349
rect 20076 3544 20128 3596
rect 20352 3544 20404 3596
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 19064 3476 19116 3528
rect 20812 3544 20864 3596
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 21456 3476 21508 3528
rect 21272 3408 21324 3460
rect 18972 3340 19024 3392
rect 19892 3340 19944 3392
rect 20444 3340 20496 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 4804 3136 4856 3188
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 6092 3179 6144 3188
rect 6092 3145 6101 3179
rect 6101 3145 6135 3179
rect 6135 3145 6144 3179
rect 6092 3136 6144 3145
rect 8484 3136 8536 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 10048 3136 10100 3188
rect 10508 3136 10560 3188
rect 10876 3136 10928 3188
rect 12164 3136 12216 3188
rect 13912 3136 13964 3188
rect 16120 3136 16172 3188
rect 19064 3179 19116 3188
rect 5632 3111 5684 3120
rect 5632 3077 5641 3111
rect 5641 3077 5675 3111
rect 5675 3077 5684 3111
rect 5632 3068 5684 3077
rect 1216 2932 1268 2984
rect 3976 2932 4028 2984
rect 4896 2932 4948 2984
rect 5080 2932 5132 2984
rect 5356 2932 5408 2984
rect 5724 2932 5776 2984
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 7288 2932 7340 2984
rect 7656 2932 7708 2984
rect 8760 2932 8812 2984
rect 9220 3000 9272 3052
rect 18696 3068 18748 3120
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 20260 3179 20312 3188
rect 20260 3145 20269 3179
rect 20269 3145 20303 3179
rect 20303 3145 20312 3179
rect 20260 3136 20312 3145
rect 20628 3179 20680 3188
rect 20628 3145 20637 3179
rect 20637 3145 20671 3179
rect 20671 3145 20680 3179
rect 20628 3136 20680 3145
rect 19524 3068 19576 3120
rect 9312 2932 9364 2984
rect 10048 2932 10100 2984
rect 11244 2932 11296 2984
rect 12808 2932 12860 2984
rect 204 2864 256 2916
rect 1676 2864 1728 2916
rect 2320 2864 2372 2916
rect 3056 2864 3108 2916
rect 8208 2864 8260 2916
rect 9956 2864 10008 2916
rect 12072 2864 12124 2916
rect 12716 2864 12768 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 2596 2839 2648 2848
rect 2596 2805 2605 2839
rect 2605 2805 2639 2839
rect 2639 2805 2648 2839
rect 2596 2796 2648 2805
rect 3884 2839 3936 2848
rect 3884 2805 3893 2839
rect 3893 2805 3927 2839
rect 3927 2805 3936 2839
rect 3884 2796 3936 2805
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 8668 2796 8720 2848
rect 10048 2796 10100 2848
rect 10140 2796 10192 2848
rect 14004 3000 14056 3052
rect 15292 3000 15344 3052
rect 16304 3000 16356 3052
rect 16580 3000 16632 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 18604 3000 18656 3052
rect 19800 3043 19852 3052
rect 19800 3009 19809 3043
rect 19809 3009 19843 3043
rect 19843 3009 19852 3043
rect 19800 3000 19852 3009
rect 20444 3000 20496 3052
rect 21364 3000 21416 3052
rect 14556 2932 14608 2984
rect 15936 2932 15988 2984
rect 16120 2932 16172 2984
rect 13268 2796 13320 2848
rect 14740 2796 14792 2848
rect 15108 2864 15160 2916
rect 16212 2907 16264 2916
rect 16212 2873 16221 2907
rect 16221 2873 16255 2907
rect 16255 2873 16264 2907
rect 16212 2864 16264 2873
rect 17408 2932 17460 2984
rect 17592 2975 17644 2984
rect 17592 2941 17601 2975
rect 17601 2941 17635 2975
rect 17635 2941 17644 2975
rect 17592 2932 17644 2941
rect 18420 2932 18472 2984
rect 16488 2864 16540 2916
rect 18972 2864 19024 2916
rect 15568 2796 15620 2848
rect 15844 2839 15896 2848
rect 15844 2805 15853 2839
rect 15853 2805 15887 2839
rect 15887 2805 15896 2839
rect 15844 2796 15896 2805
rect 17132 2839 17184 2848
rect 17132 2805 17141 2839
rect 17141 2805 17175 2839
rect 17175 2805 17184 2839
rect 17132 2796 17184 2805
rect 18512 2796 18564 2848
rect 19708 2932 19760 2984
rect 19892 2975 19944 2984
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 20628 2932 20680 2984
rect 22652 2932 22704 2984
rect 19156 2864 19208 2916
rect 21272 2907 21324 2916
rect 21272 2873 21281 2907
rect 21281 2873 21315 2907
rect 21315 2873 21324 2907
rect 21272 2864 21324 2873
rect 19432 2796 19484 2848
rect 20536 2796 20588 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 1676 2567 1728 2576
rect 1676 2533 1685 2567
rect 1685 2533 1719 2567
rect 1719 2533 1728 2567
rect 1676 2524 1728 2533
rect 2228 2456 2280 2508
rect 2596 2499 2648 2508
rect 2596 2465 2605 2499
rect 2605 2465 2639 2499
rect 2639 2465 2648 2499
rect 2596 2456 2648 2465
rect 3056 2499 3108 2508
rect 3056 2465 3065 2499
rect 3065 2465 3099 2499
rect 3099 2465 3108 2499
rect 3056 2456 3108 2465
rect 3884 2456 3936 2508
rect 4344 2456 4396 2508
rect 5172 2456 5224 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6552 2456 6604 2508
rect 6920 2456 6972 2508
rect 7748 2592 7800 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 9404 2592 9456 2644
rect 9680 2524 9732 2576
rect 9864 2524 9916 2576
rect 10876 2592 10928 2644
rect 11060 2592 11112 2644
rect 11888 2592 11940 2644
rect 12900 2592 12952 2644
rect 14740 2592 14792 2644
rect 15844 2592 15896 2644
rect 16488 2592 16540 2644
rect 12624 2524 12676 2576
rect 17132 2524 17184 2576
rect 18420 2592 18472 2644
rect 20076 2635 20128 2644
rect 18604 2524 18656 2576
rect 20076 2601 20085 2635
rect 20085 2601 20119 2635
rect 20119 2601 20128 2635
rect 20076 2592 20128 2601
rect 7380 2388 7432 2440
rect 7840 2456 7892 2508
rect 16396 2456 16448 2508
rect 19064 2456 19116 2508
rect 20720 2456 20772 2508
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 2504 2252 2556 2304
rect 3148 2252 3200 2304
rect 5264 2295 5316 2304
rect 5264 2261 5273 2295
rect 5273 2261 5307 2295
rect 5307 2261 5316 2295
rect 5264 2252 5316 2261
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 6184 2295 6236 2304
rect 6184 2261 6193 2295
rect 6193 2261 6227 2295
rect 6227 2261 6236 2295
rect 6184 2252 6236 2261
rect 8392 2320 8444 2372
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 10600 2431 10652 2440
rect 8576 2388 8628 2397
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 13912 2388 13964 2440
rect 14556 2388 14608 2440
rect 9036 2252 9088 2304
rect 12164 2320 12216 2372
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 10968 2252 11020 2304
rect 11704 2252 11756 2304
rect 15568 2252 15620 2304
rect 15844 2320 15896 2372
rect 16488 2320 16540 2372
rect 17132 2320 17184 2372
rect 17684 2320 17736 2372
rect 20628 2320 20680 2372
rect 19064 2252 19116 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 1768 2048 1820 2100
rect 7564 2048 7616 2100
rect 15568 2048 15620 2100
rect 19616 2048 19668 2100
rect 17592 1980 17644 2032
rect 6184 1912 6236 1964
rect 18972 1912 19024 1964
rect 2504 1844 2556 1896
rect 1768 1776 1820 1828
rect 2596 1776 2648 1828
rect 664 1708 716 1760
rect 2228 1708 2280 1760
rect 5264 1844 5316 1896
rect 15384 1844 15436 1896
rect 3424 1776 3476 1828
rect 4344 1776 4396 1828
rect 6000 1776 6052 1828
rect 9496 1776 9548 1828
rect 17960 1776 18012 1828
rect 2872 1708 2924 1760
rect 3884 1708 3936 1760
rect 5724 1708 5776 1760
rect 17868 1708 17920 1760
rect 3148 1640 3200 1692
rect 10232 1640 10284 1692
rect 14280 1572 14332 1624
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 20626 22672 20682 22681
rect 20626 22607 20682 22616
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 5736 20398 5764 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 5920 19310 5948 20198
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 17236 20058 17264 22200
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 7300 12434 7328 19178
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 11992 18970 12020 19246
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7024 12406 7328 12434
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 1676 11552 1728 11558
rect 1674 11520 1676 11529
rect 1728 11520 1730 11529
rect 1674 11455 1730 11464
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4802 3496 4858 3505
rect 4802 3431 4858 3440
rect 1216 3392 1268 3398
rect 1216 3334 1268 3340
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 1228 2990 1256 3334
rect 1216 2984 1268 2990
rect 3976 2984 4028 2990
rect 1216 2926 1268 2932
rect 1582 2952 1638 2961
rect 204 2916 256 2922
rect 204 2858 256 2864
rect 216 800 244 2858
rect 664 1760 716 1766
rect 664 1702 716 1708
rect 676 800 704 1702
rect 1228 800 1256 2926
rect 3976 2926 4028 2932
rect 1582 2887 1638 2896
rect 1676 2916 1728 2922
rect 1596 2854 1624 2887
rect 1676 2858 1728 2864
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1688 2582 1716 2858
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 2240 2514 2268 2790
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 2106 1808 2246
rect 1768 2100 1820 2106
rect 1768 2042 1820 2048
rect 1768 1828 1820 1834
rect 1768 1770 1820 1776
rect 1780 800 1808 1770
rect 2240 1766 2268 2450
rect 2228 1760 2280 1766
rect 2228 1702 2280 1708
rect 2332 800 2360 2858
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 2514 2636 2790
rect 3068 2514 3096 2858
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3896 2514 3924 2790
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 1902 2544 2246
rect 2504 1896 2556 1902
rect 2504 1838 2556 1844
rect 2608 1834 2636 2450
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 2596 1828 2648 1834
rect 2596 1770 2648 1776
rect 2872 1760 2924 1766
rect 2872 1702 2924 1708
rect 2884 800 2912 1702
rect 3160 1698 3188 2246
rect 3424 1828 3476 1834
rect 3424 1770 3476 1776
rect 3148 1692 3200 1698
rect 3148 1634 3200 1640
rect 3436 800 3464 1770
rect 3896 1766 3924 2450
rect 3884 1760 3936 1766
rect 3884 1702 3936 1708
rect 3988 800 4016 2926
rect 4356 2514 4384 3334
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4816 3194 4844 3431
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4908 2990 4936 3878
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 3074 5120 3334
rect 5184 3194 5212 6870
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5368 4826 5396 5034
rect 5828 4826 5856 5102
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5368 4282 5396 4762
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4282 6868 4422
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6932 4078 6960 4966
rect 6920 4072 6972 4078
rect 7024 4049 7052 12406
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8128 8634 8156 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7116 4690 7144 6054
rect 7668 5710 7696 6122
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7668 5370 7696 5646
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7760 5352 7788 5510
rect 8220 5409 8248 6598
rect 8312 5914 8340 17682
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8206 5400 8262 5409
rect 7932 5364 7984 5370
rect 7760 5324 7932 5352
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7300 5137 7328 5170
rect 7286 5128 7342 5137
rect 7286 5063 7342 5072
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7208 4078 7236 4490
rect 7196 4072 7248 4078
rect 6920 4014 6972 4020
rect 7010 4040 7066 4049
rect 7196 4014 7248 4020
rect 7010 3975 7066 3984
rect 7288 4004 7340 4010
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5092 3046 5212 3074
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4908 2774 4936 2926
rect 4816 2746 4936 2774
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4356 1834 4384 2450
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4344 1828 4396 1834
rect 4344 1770 4396 1776
rect 4816 1442 4844 2746
rect 4540 1414 4844 1442
rect 4540 800 4568 1414
rect 5092 800 5120 2926
rect 5184 2514 5212 3046
rect 5368 2990 5396 3878
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5552 2553 5580 3334
rect 5632 3120 5684 3126
rect 5630 3088 5632 3097
rect 5684 3088 5686 3097
rect 5630 3023 5686 3032
rect 5736 2990 5764 3878
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5736 2774 5764 2926
rect 5644 2746 5764 2774
rect 5538 2544 5594 2553
rect 5172 2508 5224 2514
rect 5538 2479 5540 2488
rect 5172 2450 5224 2456
rect 5592 2479 5594 2488
rect 5540 2450 5592 2456
rect 5184 2417 5212 2450
rect 5170 2408 5226 2417
rect 5170 2343 5226 2352
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5276 1902 5304 2246
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 5644 800 5672 2746
rect 6012 2514 6040 3878
rect 6090 3632 6146 3641
rect 6090 3567 6146 3576
rect 6104 3194 6132 3567
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2514 6592 2790
rect 6748 2774 6776 3878
rect 7024 3738 7052 3975
rect 7288 3946 7340 3952
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 2990 7052 3334
rect 7300 3233 7328 3946
rect 7286 3224 7342 3233
rect 7286 3159 7342 3168
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6748 2746 6960 2774
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5736 1766 5764 2246
rect 6012 1834 6040 2450
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 6196 1970 6224 2246
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 6000 1828 6052 1834
rect 6564 1816 6592 2450
rect 6000 1770 6052 1776
rect 6196 1788 6592 1816
rect 5724 1760 5776 1766
rect 5724 1702 5776 1708
rect 6196 800 6224 1788
rect 6748 800 6776 2746
rect 6932 2514 6960 2746
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7300 800 7328 2926
rect 7392 2446 7420 4626
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7656 4072 7708 4078
rect 7760 4060 7788 5324
rect 8206 5335 8262 5344
rect 7932 5306 7984 5312
rect 8220 5030 8248 5335
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8312 4826 8340 5646
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8404 5098 8432 5578
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8404 4554 8432 5034
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8496 4434 8524 7958
rect 8588 6118 8616 13738
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 9110 8708 11494
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8680 8090 8708 9046
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5914 8616 6054
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8680 5370 8708 6190
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8772 5234 8800 6054
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8864 5114 8892 14418
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9048 5370 9076 7142
rect 9140 7002 9168 7142
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8956 5234 8984 5306
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8772 5086 8892 5114
rect 8680 4690 8708 5034
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 7708 4032 7788 4060
rect 8404 4406 8524 4434
rect 7656 4014 7708 4020
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7484 3670 7512 3946
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7484 3398 7512 3606
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7576 2106 7604 4014
rect 7668 2990 7696 4014
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7760 2650 7788 3470
rect 8208 2916 8260 2922
rect 8260 2876 8340 2904
rect 8208 2858 8260 2864
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8312 2650 8340 2876
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7852 800 7880 2450
rect 8404 2378 8432 4406
rect 8772 3738 8800 5086
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8864 4758 8892 4966
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8496 3194 8524 3538
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8496 2774 8524 3130
rect 8772 2990 8800 3470
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8496 2746 8616 2774
rect 8588 2446 8616 2746
rect 8680 2553 8708 2790
rect 8666 2544 8722 2553
rect 8666 2479 8722 2488
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8864 1442 8892 3334
rect 8404 1414 8892 1442
rect 8404 800 8432 1414
rect 8956 800 8984 4218
rect 9048 2310 9076 4966
rect 9232 4593 9260 8298
rect 9218 4584 9274 4593
rect 9218 4519 9274 4528
rect 9232 4282 9260 4519
rect 9324 4486 9352 11562
rect 9508 7546 9536 18158
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 9178 9812 14418
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11716 9654 11744 10610
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9416 6866 9444 7346
rect 9494 6896 9550 6905
rect 9404 6860 9456 6866
rect 9494 6831 9550 6840
rect 9404 6802 9456 6808
rect 9416 6458 9444 6802
rect 9508 6662 9536 6831
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9508 5778 9536 6598
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 4690 9444 5306
rect 9600 4826 9628 8910
rect 9692 8090 9720 8978
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8430 9812 8774
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 10060 7750 10088 9454
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 8634 11008 8978
rect 11716 8974 11744 9590
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 7954 10180 8298
rect 10980 8022 11008 8570
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11716 7954 11744 8910
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 9692 5370 9720 5607
rect 9784 5574 9812 6122
rect 10060 5914 10088 7686
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10152 5710 10180 7890
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9784 5302 9812 5510
rect 9862 5400 9918 5409
rect 9862 5335 9864 5344
rect 9916 5335 9918 5344
rect 9864 5306 9916 5312
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9862 5264 9918 5273
rect 9862 5199 9918 5208
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9496 4752 9548 4758
rect 9494 4720 9496 4729
rect 9548 4720 9550 4729
rect 9404 4684 9456 4690
rect 9494 4655 9550 4664
rect 9680 4684 9732 4690
rect 9404 4626 9456 4632
rect 9680 4626 9732 4632
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9232 3058 9260 3606
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9324 2417 9352 2926
rect 9416 2650 9444 4626
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9508 4078 9536 4150
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9692 2582 9720 4626
rect 9784 4078 9812 4966
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 3194 9812 3538
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 2582 9904 5199
rect 10140 4616 10192 4622
rect 10138 4584 10140 4593
rect 10192 4584 10194 4593
rect 10138 4519 10194 4528
rect 10138 4176 10194 4185
rect 10048 4140 10100 4146
rect 10138 4111 10194 4120
rect 10048 4082 10100 4088
rect 10060 4026 10088 4082
rect 10152 4078 10180 4111
rect 9968 3998 10088 4026
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 9968 3398 9996 3998
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3670 10088 3878
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 2922 9996 3334
rect 10138 3224 10194 3233
rect 10048 3188 10100 3194
rect 10138 3159 10194 3168
rect 10048 3130 10100 3136
rect 10060 2990 10088 3130
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 10152 2854 10180 3159
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9310 2408 9366 2417
rect 9310 2343 9366 2352
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9496 1828 9548 1834
rect 9496 1770 9548 1776
rect 9508 800 9536 1770
rect 10060 800 10088 2790
rect 10244 1698 10272 7210
rect 10704 7002 10732 7346
rect 10888 7206 10916 7822
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10704 6866 10732 6938
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10888 6361 10916 7142
rect 10874 6352 10930 6361
rect 10874 6287 10930 6296
rect 11164 6254 11192 7482
rect 11702 6760 11758 6769
rect 11702 6695 11758 6704
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11716 6458 11744 6695
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 10692 6248 10744 6254
rect 11152 6248 11204 6254
rect 10692 6190 10744 6196
rect 10874 6216 10930 6225
rect 10704 5846 10732 6190
rect 11152 6190 11204 6196
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 10874 6151 10930 6160
rect 10888 6118 10916 6151
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10704 5574 10732 5782
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 11164 5370 11192 6190
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 4758 10732 5034
rect 11152 5024 11204 5030
rect 11256 5012 11284 5782
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11336 5024 11388 5030
rect 11256 4984 11336 5012
rect 11152 4966 11204 4972
rect 11336 4966 11388 4972
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10598 4040 10654 4049
rect 10598 3975 10600 3984
rect 10652 3975 10654 3984
rect 10600 3946 10652 3952
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10232 1692 10284 1698
rect 10232 1634 10284 1640
rect 10520 1442 10548 3130
rect 10612 2446 10640 3538
rect 10888 3194 10916 4558
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10888 2650 10916 3130
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10980 2310 11008 4626
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11072 2650 11100 4082
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10520 1414 10640 1442
rect 10612 800 10640 1414
rect 11164 800 11192 4966
rect 11348 4690 11376 4966
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11624 3738 11652 4014
rect 11716 4010 11744 6190
rect 11808 4826 11836 17070
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11900 9654 11928 14894
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11900 3942 11928 8366
rect 11992 7546 12020 18770
rect 16776 18358 16804 19178
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12176 17338 12204 18158
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12176 12434 12204 13806
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 12084 12406 12204 12434
rect 12084 8430 12112 12406
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12084 7342 12112 8230
rect 12176 8106 12204 10406
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12268 9110 12296 9522
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12176 8078 12296 8106
rect 12360 8090 12388 9318
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12176 7410 12204 7890
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12176 7002 12204 7346
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5778 12112 6054
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4826 12020 4966
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 12084 4593 12112 5714
rect 12070 4584 12126 4593
rect 12070 4519 12126 4528
rect 12268 4298 12296 8078
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12360 7546 12388 7890
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12360 6662 12388 7482
rect 12452 6662 12480 8230
rect 12728 7546 12756 8366
rect 12912 7750 12940 10474
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12636 6866 12664 7210
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 7002 12848 7142
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 6254 12480 6598
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12636 5778 12664 6258
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12360 4604 12388 5646
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4758 12480 4966
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12360 4576 12480 4604
rect 11992 4270 12296 4298
rect 11992 4078 12020 4270
rect 12084 4146 12388 4162
rect 12084 4140 12400 4146
rect 12084 4134 12348 4140
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11256 2990 11284 3538
rect 12084 3398 12112 4134
rect 12348 4082 12400 4088
rect 12452 3738 12480 4576
rect 12636 4554 12664 5714
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4321 12572 4422
rect 12530 4312 12586 4321
rect 12530 4247 12586 4256
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11900 2650 11928 3334
rect 12084 2922 12112 3334
rect 12176 3194 12204 3334
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12636 2582 12664 3878
rect 12728 3505 12756 6054
rect 13004 4690 13032 9318
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 6322 13124 7142
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13188 5914 13216 6734
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13188 5166 13216 5850
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13096 4690 13124 5102
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12714 3496 12770 3505
rect 12714 3431 12770 3440
rect 12820 2990 12848 4422
rect 13280 3942 13308 13330
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13556 11354 13584 11834
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 10266 13676 11154
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13556 9722 13584 10202
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8430 13400 8774
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13372 7886 13400 8366
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13360 7880 13412 7886
rect 13544 7880 13596 7886
rect 13360 7822 13412 7828
rect 13542 7848 13544 7857
rect 13596 7848 13598 7857
rect 13542 7783 13598 7792
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 4826 13400 6734
rect 13464 6458 13492 6802
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13556 4486 13584 7210
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 800 11744 2246
rect 12176 800 12204 2314
rect 12728 800 12756 2858
rect 12912 2650 12940 3878
rect 13648 3641 13676 7890
rect 13740 6254 13768 11766
rect 13832 6730 13860 17070
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13924 10810 13952 11018
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14016 9518 14044 11494
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 14016 6254 14044 9454
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 8294 14136 8978
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14108 7886 14136 8230
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14200 6746 14228 10066
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 6866 14320 9862
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14200 6718 14320 6746
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14108 5234 14136 6122
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13740 4214 13768 4694
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13740 4078 13768 4150
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13832 3670 13860 4082
rect 13820 3664 13872 3670
rect 13634 3632 13690 3641
rect 13820 3606 13872 3612
rect 13634 3567 13690 3576
rect 13832 3482 13860 3606
rect 14016 3534 14044 5102
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 14108 3942 14136 4626
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14200 3670 14228 6054
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14004 3528 14056 3534
rect 13832 3454 13952 3482
rect 14004 3470 14056 3476
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13280 800 13308 2790
rect 13832 800 13860 3334
rect 13924 3194 13952 3454
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13924 2446 13952 3130
rect 14016 3058 14044 3470
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14292 1630 14320 6718
rect 14384 6254 14412 9318
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14476 8022 14504 8910
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14568 7818 14596 15506
rect 16040 15162 16068 15914
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16316 14006 16344 14418
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14648 12300 14700 12306
rect 15936 12300 15988 12306
rect 14648 12242 14700 12248
rect 15856 12260 15936 12288
rect 14660 11218 14688 12242
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14660 10538 14688 11154
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14648 10192 14700 10198
rect 14646 10160 14648 10169
rect 14700 10160 14702 10169
rect 14752 10130 14780 12038
rect 15304 11694 15332 12038
rect 15856 11762 15884 12260
rect 15936 12242 15988 12248
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15488 10810 15516 11154
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14646 10095 14702 10104
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14660 7993 14688 9930
rect 15304 9722 15332 9998
rect 15488 9994 15516 10746
rect 15672 10266 15700 11494
rect 15764 11354 15792 11494
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15856 11082 15884 11698
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15948 10169 15976 10542
rect 15934 10160 15990 10169
rect 15934 10095 15990 10104
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14752 8634 14780 9454
rect 15028 9364 15056 9454
rect 15028 9336 15240 9364
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15212 9042 15240 9336
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15212 8838 15240 8978
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14646 7984 14702 7993
rect 14646 7919 14702 7928
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14832 7336 14884 7342
rect 14752 7296 14832 7324
rect 14556 7200 14608 7206
rect 14476 7160 14556 7188
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14476 5642 14504 7160
rect 14556 7142 14608 7148
rect 14752 6798 14780 7296
rect 14832 7278 14884 7284
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14556 6656 14608 6662
rect 14554 6624 14556 6633
rect 14608 6624 14610 6633
rect 14554 6559 14610 6568
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14554 5808 14610 5817
rect 14554 5743 14610 5752
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14476 5030 14504 5578
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14280 1624 14332 1630
rect 14280 1566 14332 1572
rect 14384 800 14412 4490
rect 14476 4049 14504 4966
rect 14568 4690 14596 5743
rect 14752 5302 14780 6326
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 15212 5846 15240 8366
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15672 7206 15700 7890
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6497 15332 6734
rect 15290 6488 15346 6497
rect 15396 6458 15424 6802
rect 15290 6423 15346 6432
rect 15384 6452 15436 6458
rect 15304 6254 15332 6423
rect 15384 6394 15436 6400
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15396 5710 15424 6394
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5930 15608 6054
rect 15580 5902 15700 5930
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15384 5704 15436 5710
rect 15304 5652 15384 5658
rect 15304 5646 15436 5652
rect 15304 5630 15424 5646
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14752 4282 14780 4626
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 15212 4078 15240 5034
rect 15304 4622 15332 5630
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15200 4072 15252 4078
rect 14462 4040 14518 4049
rect 15200 4014 15252 4020
rect 14462 3975 14518 3984
rect 15292 4004 15344 4010
rect 14476 3738 14504 3975
rect 15292 3946 15344 3952
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14568 2990 14596 3878
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14568 2446 14596 2926
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14660 1442 14688 3878
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 2922 15148 3538
rect 15304 3398 15332 3946
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15304 3058 15332 3334
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14752 2650 14780 2790
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 15396 1902 15424 4966
rect 15488 4826 15516 4966
rect 15580 4826 15608 5714
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 14660 1414 14964 1442
rect 14936 800 14964 1414
rect 15488 800 15516 4490
rect 15568 2848 15620 2854
rect 15566 2816 15568 2825
rect 15620 2816 15622 2825
rect 15566 2751 15622 2760
rect 15672 2774 15700 5902
rect 15764 5250 15792 7958
rect 15856 7954 15884 9930
rect 15948 9722 15976 9998
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15948 9178 15976 9386
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15948 7818 15976 9114
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 5642 15884 7142
rect 16040 6866 16068 13126
rect 16120 11688 16172 11694
rect 16488 11688 16540 11694
rect 16172 11636 16252 11642
rect 16120 11630 16252 11636
rect 16488 11630 16540 11636
rect 16132 11614 16252 11630
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16132 8090 16160 9998
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16224 7970 16252 11614
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16316 10538 16344 11018
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8072 16344 9318
rect 16408 9110 16436 9658
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16396 8084 16448 8090
rect 16316 8044 16396 8072
rect 16396 8026 16448 8032
rect 16394 7984 16450 7993
rect 16224 7942 16344 7970
rect 16316 7206 16344 7942
rect 16394 7919 16450 7928
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16040 6610 16068 6802
rect 15948 6582 16068 6610
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15764 5222 15884 5250
rect 15948 5234 15976 6582
rect 15856 3097 15884 5222
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15842 3088 15898 3097
rect 15842 3023 15898 3032
rect 15948 2990 15976 4966
rect 16132 4826 16160 7142
rect 16304 6792 16356 6798
rect 16224 6752 16304 6780
rect 16224 6186 16252 6752
rect 16304 6734 16356 6740
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16210 4720 16266 4729
rect 16210 4655 16266 4664
rect 16026 4312 16082 4321
rect 16026 4247 16082 4256
rect 16040 4146 16068 4247
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15672 2746 15792 2774
rect 15764 2530 15792 2746
rect 15856 2650 15884 2790
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15764 2502 15884 2530
rect 15856 2378 15884 2502
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15580 2106 15608 2246
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 16040 800 16068 3674
rect 16224 3670 16252 4655
rect 16316 4570 16344 6598
rect 16408 6254 16436 7919
rect 16500 7546 16528 11630
rect 16592 10266 16620 15982
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16868 11218 16896 12650
rect 16960 12306 16988 12718
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17052 12186 17080 12650
rect 16960 12158 17080 12186
rect 16960 12102 16988 12158
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16960 11150 16988 12038
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 17052 11354 17080 11562
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17052 10690 17080 11086
rect 16960 10662 17080 10690
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16592 6730 16620 7346
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16592 6322 16620 6666
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16500 6118 16528 6190
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16486 5944 16542 5953
rect 16486 5879 16488 5888
rect 16540 5879 16542 5888
rect 16488 5850 16540 5856
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16500 5681 16528 5714
rect 16486 5672 16542 5681
rect 16486 5607 16542 5616
rect 16500 5234 16528 5607
rect 16578 5264 16634 5273
rect 16488 5228 16540 5234
rect 16578 5199 16634 5208
rect 16488 5170 16540 5176
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4758 16436 4966
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16316 4542 16436 4570
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16132 3194 16160 3334
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16132 2990 16160 3130
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16224 2922 16252 3606
rect 16316 3534 16344 4082
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16316 2446 16344 2994
rect 16408 2514 16436 4542
rect 16500 2922 16528 5034
rect 16592 5001 16620 5199
rect 16684 5166 16712 10406
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16776 9178 16804 10134
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 9586 16896 9862
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16776 7750 16804 8434
rect 16960 7834 16988 10662
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17052 9654 17080 10542
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17144 8362 17172 13874
rect 17420 13462 17448 20198
rect 17604 20058 17632 20334
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17972 19174 18000 20198
rect 18616 19990 18644 21655
rect 18970 21312 19026 21321
rect 18970 21247 19026 21256
rect 18984 20534 19012 21247
rect 19522 20904 19578 20913
rect 19522 20839 19578 20848
rect 19536 20534 19564 20839
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 20640 20466 20668 22607
rect 21546 22264 21602 22273
rect 21546 22199 21602 22208
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20810 20360 20866 20369
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 20076 20324 20128 20330
rect 20810 20295 20812 20304
rect 20076 20266 20128 20272
rect 20864 20295 20866 20304
rect 21088 20324 21140 20330
rect 20812 20266 20864 20272
rect 21088 20266 21140 20272
rect 18800 20058 18828 20266
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18604 19984 18656 19990
rect 18604 19926 18656 19932
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 19720 19514 19748 19858
rect 20088 19514 20116 20266
rect 20810 19952 20866 19961
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20628 19916 20680 19922
rect 20810 19887 20812 19896
rect 20628 19858 20680 19864
rect 20864 19887 20866 19896
rect 20812 19858 20864 19864
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 18708 18970 18736 19246
rect 20088 18970 20116 19246
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 11098 17356 12242
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17604 11694 17632 12174
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17420 11286 17448 11494
rect 17512 11354 17540 11494
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17328 11070 17448 11098
rect 17420 10742 17448 11070
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17420 10198 17448 10678
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17236 7993 17264 9930
rect 17604 9178 17632 10066
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17222 7984 17278 7993
rect 17222 7919 17278 7928
rect 16960 7806 17080 7834
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16776 7274 16804 7686
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16776 5710 16804 6802
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16672 5024 16724 5030
rect 16578 4992 16634 5001
rect 16672 4966 16724 4972
rect 16578 4927 16634 4936
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16592 3058 16620 3334
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16684 2774 16712 4966
rect 16960 4758 16988 7686
rect 17052 7206 17080 7806
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 17144 6497 17172 6666
rect 17130 6488 17186 6497
rect 17130 6423 17186 6432
rect 17144 6254 17172 6423
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16776 3738 16804 4490
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16868 3602 16896 3946
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 17052 2961 17080 5578
rect 17144 4146 17172 6190
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5166 17264 6054
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17328 4078 17356 8502
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7546 17448 8230
rect 17604 8022 17632 8774
rect 17696 8634 17724 16594
rect 17972 15706 18000 16594
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17788 11762 17816 13806
rect 17972 13530 18000 14350
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18524 13394 18552 13738
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17880 12306 17908 13194
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17788 9353 17816 11698
rect 17880 11218 17908 12038
rect 17972 11762 18000 12310
rect 18064 12102 18092 12650
rect 18432 12186 18460 12718
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18524 12374 18552 12582
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18156 12158 18460 12186
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 11212 17920 11218
rect 17920 11172 18000 11200
rect 17868 11154 17920 11160
rect 17859 10600 17911 10606
rect 17859 10542 17911 10548
rect 17880 9586 17908 10542
rect 17972 9761 18000 11172
rect 17958 9752 18014 9761
rect 17958 9687 18014 9696
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17774 9344 17830 9353
rect 17774 9279 17830 9288
rect 17776 8968 17828 8974
rect 17972 8945 18000 9590
rect 17776 8910 17828 8916
rect 17958 8936 18014 8945
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17604 7410 17632 7958
rect 17682 7848 17738 7857
rect 17682 7783 17738 7792
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17420 6780 17448 7142
rect 17512 6934 17540 7142
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17604 6780 17632 6870
rect 17420 6752 17632 6780
rect 17420 6633 17448 6752
rect 17406 6624 17462 6633
rect 17406 6559 17462 6568
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17420 2990 17448 6559
rect 17696 6440 17724 7783
rect 17604 6412 17724 6440
rect 17604 6118 17632 6412
rect 17682 6352 17738 6361
rect 17682 6287 17738 6296
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 5137 17540 5714
rect 17498 5128 17554 5137
rect 17498 5063 17554 5072
rect 17604 2990 17632 6054
rect 17696 5846 17724 6287
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 3670 17724 4422
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17408 2984 17460 2990
rect 17038 2952 17094 2961
rect 17408 2926 17460 2932
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17038 2887 17094 2896
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 16592 2746 16712 2774
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16500 2378 16528 2586
rect 16488 2372 16540 2378
rect 16488 2314 16540 2320
rect 16592 800 16620 2746
rect 17144 2582 17172 2790
rect 17788 2774 17816 8910
rect 18064 8922 18092 11834
rect 18156 10305 18184 12158
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18616 11898 18644 18770
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 18892 13870 18920 14214
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 19260 13852 19288 14214
rect 19340 13864 19392 13870
rect 19260 13824 19340 13852
rect 18708 13462 18736 13806
rect 18696 13456 18748 13462
rect 18696 13398 18748 13404
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18708 11257 18736 13398
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18694 11248 18750 11257
rect 18694 11183 18750 11192
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18800 10690 18828 12922
rect 18892 12617 18920 13806
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 19076 13394 19104 13670
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18878 12608 18934 12617
rect 18878 12543 18934 12552
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11830 18920 12174
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18984 10713 19012 12718
rect 19076 12073 19104 13330
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19168 12782 19196 13194
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19260 12434 19288 13824
rect 19340 13806 19392 13812
rect 19628 12434 19656 18770
rect 20272 18426 20300 19858
rect 20640 19514 20668 19858
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19812 17338 19840 17682
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19168 12406 19288 12434
rect 19536 12406 19656 12434
rect 19062 12064 19118 12073
rect 19062 11999 19118 12008
rect 19168 11665 19196 12406
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11694 19288 12038
rect 19248 11688 19300 11694
rect 19154 11656 19210 11665
rect 19248 11630 19300 11636
rect 19154 11591 19210 11600
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 18970 10704 19026 10713
rect 18800 10662 18920 10690
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18142 10296 18198 10305
rect 18142 10231 18198 10240
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18340 10033 18368 10066
rect 18326 10024 18382 10033
rect 18326 9959 18382 9968
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18142 9752 18198 9761
rect 18282 9744 18578 9764
rect 18142 9687 18198 9696
rect 18156 9450 18184 9687
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18616 8922 18644 10202
rect 18708 9897 18736 10406
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18694 9888 18750 9897
rect 18694 9823 18750 9832
rect 18694 9752 18750 9761
rect 18800 9722 18828 9930
rect 18694 9687 18750 9696
rect 18788 9716 18840 9722
rect 18708 9042 18736 9687
rect 18788 9658 18840 9664
rect 18786 9616 18842 9625
rect 18786 9551 18842 9560
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18064 8894 18184 8922
rect 18616 8894 18736 8922
rect 17958 8871 18014 8880
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17880 6866 17908 7890
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6254 17908 6802
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17972 6089 18000 6938
rect 17958 6080 18014 6089
rect 17958 6015 18014 6024
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17604 2746 17816 2774
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17144 800 17172 2314
rect 17604 2038 17632 2746
rect 17684 2372 17736 2378
rect 17684 2314 17736 2320
rect 17592 2032 17644 2038
rect 17592 1974 17644 1980
rect 17696 800 17724 2314
rect 17880 1766 17908 5782
rect 17958 5672 18014 5681
rect 17958 5607 18014 5616
rect 17972 5574 18000 5607
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 5273 18000 5306
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17958 4720 18014 4729
rect 17958 4655 18014 4664
rect 17972 4554 18000 4655
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 18064 4146 18092 8774
rect 18156 8514 18184 8894
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18156 8486 18276 8514
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18156 7410 18184 8298
rect 18248 7954 18276 8486
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18524 7818 18552 7890
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18156 7041 18184 7210
rect 18142 7032 18198 7041
rect 18142 6967 18198 6976
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18156 6458 18184 6802
rect 18524 6644 18552 7414
rect 18616 6769 18644 8774
rect 18708 7585 18736 8894
rect 18800 8401 18828 9551
rect 18892 9518 18920 10662
rect 18970 10639 19026 10648
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18892 8498 18920 9318
rect 18984 9110 19012 10542
rect 19076 10010 19104 11086
rect 19260 11014 19288 11154
rect 19352 11150 19380 11494
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19536 11082 19564 12406
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19076 9982 19196 10010
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18984 8430 19012 8910
rect 18972 8424 19024 8430
rect 18786 8392 18842 8401
rect 18972 8366 19024 8372
rect 18786 8327 18842 8336
rect 18788 7880 18840 7886
rect 18786 7848 18788 7857
rect 18840 7848 18842 7857
rect 18786 7783 18842 7792
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18694 7576 18750 7585
rect 18694 7511 18750 7520
rect 18602 6760 18658 6769
rect 18602 6695 18658 6704
rect 18524 6616 18644 6644
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18616 5914 18644 6616
rect 18694 6624 18750 6633
rect 18694 6559 18750 6568
rect 18708 6186 18736 6559
rect 18696 6180 18748 6186
rect 18696 6122 18748 6128
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18800 5574 18828 7686
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18892 5370 18920 7142
rect 19076 6168 19104 9862
rect 19168 7274 19196 9982
rect 19260 7342 19288 10066
rect 19352 9518 19380 10406
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19352 8430 19380 9046
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 18984 6140 19104 6168
rect 18984 5624 19012 6140
rect 19260 5828 19288 7142
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6186 19380 6598
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19168 5800 19288 5828
rect 19168 5658 19196 5800
rect 19168 5630 19288 5658
rect 19352 5642 19380 6122
rect 18984 5596 19095 5624
rect 19067 5556 19095 5596
rect 19260 5574 19288 5630
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19248 5568 19300 5574
rect 19067 5528 19104 5556
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 19076 5166 19104 5528
rect 19248 5510 19300 5516
rect 19338 5400 19394 5409
rect 19338 5335 19394 5344
rect 19352 5234 19380 5335
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19444 5098 19472 10406
rect 19536 7478 19564 10746
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19536 6186 19564 6802
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 18602 4856 18658 4865
rect 18602 4791 18658 4800
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18616 4264 18644 4791
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18524 4236 18644 4264
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 17958 3632 18014 3641
rect 17958 3567 18014 3576
rect 17972 2961 18000 3567
rect 17958 2952 18014 2961
rect 17958 2887 18014 2896
rect 17958 2408 18014 2417
rect 17958 2343 18014 2352
rect 17972 1834 18000 2343
rect 17960 1828 18012 1834
rect 17960 1770 18012 1776
rect 17868 1760 17920 1766
rect 17868 1702 17920 1708
rect 18156 1442 18184 3946
rect 18524 3924 18552 4236
rect 18708 4078 18736 4694
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18604 3936 18656 3942
rect 18524 3896 18604 3924
rect 18604 3878 18656 3884
rect 18616 3534 18644 3878
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 3058 18644 3470
rect 18694 3360 18750 3369
rect 18694 3295 18750 3304
rect 18708 3126 18736 3295
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18432 2650 18460 2926
rect 18524 2854 18552 2994
rect 18602 2952 18658 2961
rect 18602 2887 18658 2896
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 18616 2582 18644 2887
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1414 18276 1442
rect 18248 800 18276 1414
rect 18800 800 18828 5034
rect 19246 4992 19302 5001
rect 19246 4927 19302 4936
rect 19154 4856 19210 4865
rect 19154 4791 19156 4800
rect 19208 4791 19210 4800
rect 19156 4762 19208 4768
rect 19260 4758 19288 4927
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19352 4706 19380 5034
rect 18972 4684 19024 4690
rect 19352 4678 19472 4706
rect 18972 4626 19024 4632
rect 18984 4162 19012 4626
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 18984 4134 19288 4162
rect 18984 3398 19012 4134
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 19076 3194 19104 3470
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19168 2922 19196 4014
rect 19260 4010 19288 4134
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 18972 2916 19024 2922
rect 18972 2858 19024 2864
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 18984 1970 19012 2858
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 19076 2310 19104 2450
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19076 2009 19104 2246
rect 19062 2000 19118 2009
rect 18972 1964 19024 1970
rect 19062 1935 19118 1944
rect 18972 1906 19024 1912
rect 19168 1601 19196 2858
rect 19154 1592 19210 1601
rect 19154 1527 19210 1536
rect 19352 800 19380 4558
rect 19444 4185 19472 4678
rect 19430 4176 19486 4185
rect 19430 4111 19486 4120
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19444 2854 19472 3606
rect 19536 3126 19564 5850
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19628 2106 19656 12242
rect 19720 4826 19748 12718
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19812 10606 19840 11086
rect 19800 10600 19852 10606
rect 19800 10542 19852 10548
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19812 7426 19840 10066
rect 19904 7546 19932 12718
rect 19996 11626 20024 18158
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 20272 17338 20300 18090
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20088 16794 20116 17070
rect 20364 16794 20392 17614
rect 20640 17542 20668 18770
rect 20824 18222 20852 19246
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20810 17232 20866 17241
rect 20810 17167 20812 17176
rect 20864 17167 20866 17176
rect 20812 17138 20864 17144
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20640 16794 20668 17002
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20260 16720 20312 16726
rect 20260 16662 20312 16668
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20180 16250 20208 16594
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20272 15706 20300 16662
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20088 14618 20116 15506
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20364 13530 20392 14826
rect 20456 14618 20484 15846
rect 20810 15736 20866 15745
rect 20810 15671 20866 15680
rect 20824 15638 20852 15671
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 15162 20668 15506
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20824 14346 20852 14894
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20180 12442 20208 13330
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19996 7954 20024 11154
rect 20088 11150 20116 11630
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20180 10962 20208 11562
rect 20272 11354 20300 13126
rect 20548 12306 20576 14010
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20640 12986 20668 13330
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20088 10934 20208 10962
rect 20088 10538 20116 10934
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 20088 10266 20116 10474
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20088 9518 20116 10202
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20088 9110 20116 9454
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 19984 7948 20036 7954
rect 20088 7936 20116 8842
rect 20180 8362 20208 9318
rect 20272 9042 20300 9318
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20088 7908 20208 7936
rect 19984 7890 20036 7896
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19812 7398 19932 7426
rect 20088 7410 20116 7686
rect 20180 7410 20208 7908
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19812 6866 19840 7278
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19812 6458 19840 6802
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19904 6225 19932 7398
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20272 7342 20300 8298
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20364 6746 20392 12038
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 19996 6718 20392 6746
rect 19890 6216 19946 6225
rect 19890 6151 19946 6160
rect 19996 5794 20024 6718
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 19812 5766 20024 5794
rect 20074 5808 20130 5817
rect 19812 5030 19840 5766
rect 20074 5743 20130 5752
rect 20088 5710 20116 5743
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19800 5024 19852 5030
rect 19800 4966 19852 4972
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19708 4208 19760 4214
rect 19708 4150 19760 4156
rect 19720 2990 19748 4150
rect 19798 3768 19854 3777
rect 19798 3703 19854 3712
rect 19812 3058 19840 3703
rect 19904 3670 19932 5510
rect 20088 5302 20116 5510
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 19984 5160 20036 5166
rect 20180 5148 20208 6054
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20272 5166 20300 5578
rect 20364 5370 20392 5714
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20036 5120 20208 5148
rect 20260 5160 20312 5166
rect 19984 5102 20036 5108
rect 20260 5102 20312 5108
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19904 2990 19932 3334
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19996 2774 20024 4966
rect 20548 4690 20576 9862
rect 20640 9518 20668 12582
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20732 11014 20760 11154
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10130 20760 10950
rect 20824 10266 20852 13262
rect 20916 12374 20944 13806
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 21008 11694 21036 13942
rect 21100 13410 21128 20266
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21192 18970 21220 19858
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 21376 19417 21404 19722
rect 21362 19408 21418 19417
rect 21362 19343 21418 19352
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21376 19009 21404 19178
rect 21362 19000 21418 19009
rect 21180 18964 21232 18970
rect 21362 18935 21418 18944
rect 21180 18906 21232 18912
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21192 17882 21220 18770
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21376 18601 21404 18634
rect 21362 18592 21418 18601
rect 21362 18527 21418 18536
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 18057 21404 18090
rect 21362 18048 21418 18057
rect 21362 17983 21418 17992
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21362 17640 21418 17649
rect 21362 17575 21364 17584
rect 21416 17575 21418 17584
rect 21364 17546 21416 17552
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21192 16250 21220 17002
rect 21468 16697 21496 17002
rect 21454 16688 21510 16697
rect 21364 16652 21416 16658
rect 21454 16623 21510 16632
rect 21364 16594 21416 16600
rect 21376 16289 21404 16594
rect 21362 16280 21418 16289
rect 21180 16244 21232 16250
rect 21362 16215 21418 16224
rect 21180 16186 21232 16192
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21192 14618 21220 15506
rect 21272 15360 21324 15366
rect 21376 15337 21404 15914
rect 21272 15302 21324 15308
rect 21362 15328 21418 15337
rect 21284 14929 21312 15302
rect 21362 15263 21418 15272
rect 21270 14920 21326 14929
rect 21270 14855 21326 14864
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21192 13530 21220 14418
rect 21468 14385 21496 14826
rect 21454 14376 21510 14385
rect 21364 14340 21416 14346
rect 21454 14311 21510 14320
rect 21364 14282 21416 14288
rect 21376 13977 21404 14282
rect 21362 13968 21418 13977
rect 21362 13903 21418 13912
rect 21560 13870 21588 22199
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21362 13560 21418 13569
rect 21180 13524 21232 13530
rect 21362 13495 21418 13504
rect 21180 13466 21232 13472
rect 21376 13462 21404 13495
rect 21364 13456 21416 13462
rect 21100 13382 21220 13410
rect 21364 13398 21416 13404
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21100 12986 21128 13262
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21100 12442 21128 12718
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20732 9364 20760 10066
rect 20640 9336 20760 9364
rect 20640 9042 20668 9336
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20640 8022 20668 8978
rect 20732 8634 20760 8978
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20640 7528 20668 7958
rect 20732 7818 20760 8570
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20720 7540 20772 7546
rect 20640 7500 20720 7528
rect 20720 7482 20772 7488
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20640 5710 20668 6326
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20088 3777 20116 3878
rect 20074 3768 20130 3777
rect 20180 3738 20208 4626
rect 20260 4616 20312 4622
rect 20640 4570 20668 5510
rect 20718 5128 20774 5137
rect 20718 5063 20774 5072
rect 20260 4558 20312 4564
rect 20272 4049 20300 4558
rect 20456 4542 20668 4570
rect 20258 4040 20314 4049
rect 20258 3975 20314 3984
rect 20074 3703 20130 3712
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 19904 2746 20024 2774
rect 19616 2100 19668 2106
rect 19616 2042 19668 2048
rect 19904 800 19932 2746
rect 20088 2650 20116 3538
rect 20258 3224 20314 3233
rect 20258 3159 20260 3168
rect 20312 3159 20314 3168
rect 20260 3130 20312 3136
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20364 1057 20392 3538
rect 20456 3398 20484 4542
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4214 20668 4422
rect 20628 4208 20680 4214
rect 20534 4176 20590 4185
rect 20628 4150 20680 4156
rect 20534 4111 20590 4120
rect 20548 4078 20576 4111
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20548 3890 20576 4014
rect 20548 3862 20668 3890
rect 20534 3768 20590 3777
rect 20534 3703 20590 3712
rect 20548 3534 20576 3703
rect 20640 3584 20668 3862
rect 20732 3738 20760 5063
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20824 3602 20852 7142
rect 20916 4078 20944 10406
rect 21008 4826 21036 11494
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21100 10062 21128 10406
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 20812 3596 20864 3602
rect 20640 3556 20760 3584
rect 20536 3528 20588 3534
rect 20588 3488 20668 3516
rect 20536 3470 20588 3476
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20456 3210 20484 3334
rect 20456 3182 20576 3210
rect 20640 3194 20668 3488
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20350 1048 20406 1057
rect 20350 983 20406 992
rect 20456 800 20484 2994
rect 20548 2854 20576 3182
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12714 0 12770 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19890 0 19946 800
rect 20442 0 20498 800
rect 20548 649 20576 2382
rect 20640 2378 20668 2926
rect 20732 2514 20760 3556
rect 20812 3538 20864 3544
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 21008 800 21036 3946
rect 21100 2825 21128 9318
rect 21192 5953 21220 13382
rect 21270 13016 21326 13025
rect 21270 12951 21272 12960
rect 21324 12951 21326 12960
rect 21272 12922 21324 12928
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21284 11014 21312 11494
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21178 5944 21234 5953
rect 21178 5879 21234 5888
rect 21192 4298 21220 5879
rect 21284 4486 21312 6598
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21192 4270 21312 4298
rect 21284 4214 21312 4270
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 21284 2922 21312 3402
rect 21376 3058 21404 5510
rect 22006 5400 22062 5409
rect 22062 5358 22140 5386
rect 22006 5335 22062 5344
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21468 3534 21496 4422
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21086 2816 21142 2825
rect 21086 2751 21142 2760
rect 20534 640 20590 649
rect 20534 575 20590 584
rect 20994 0 21050 800
rect 21284 241 21312 2858
rect 21560 800 21588 5238
rect 22112 800 22140 5358
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22664 800 22692 2926
rect 21270 232 21326 241
rect 21270 167 21326 176
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
<< via2 >>
rect 20626 22616 20682 22672
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 18602 21664 18658 21720
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 1674 11500 1676 11520
rect 1676 11500 1728 11520
rect 1728 11500 1730 11520
rect 1674 11464 1730 11500
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4802 3440 4858 3496
rect 1582 2896 1638 2952
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7286 5072 7342 5128
rect 7010 3984 7066 4040
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5630 3068 5632 3088
rect 5632 3068 5684 3088
rect 5684 3068 5686 3088
rect 5630 3032 5686 3068
rect 5538 2508 5594 2544
rect 5538 2488 5540 2508
rect 5540 2488 5592 2508
rect 5592 2488 5594 2508
rect 5170 2352 5226 2408
rect 6090 3576 6146 3632
rect 7286 3168 7342 3224
rect 8206 5344 8262 5400
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8666 2488 8722 2544
rect 9218 4528 9274 4584
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 9494 6840 9550 6896
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 9678 5616 9734 5672
rect 9862 5364 9918 5400
rect 9862 5344 9864 5364
rect 9864 5344 9916 5364
rect 9916 5344 9918 5364
rect 9862 5208 9918 5264
rect 9494 4700 9496 4720
rect 9496 4700 9548 4720
rect 9548 4700 9550 4720
rect 9494 4664 9550 4700
rect 10138 4564 10140 4584
rect 10140 4564 10192 4584
rect 10192 4564 10194 4584
rect 10138 4528 10194 4564
rect 10138 4120 10194 4176
rect 10138 3168 10194 3224
rect 9310 2352 9366 2408
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 10874 6296 10930 6352
rect 11702 6704 11758 6760
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 10874 6160 10930 6216
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 10598 4004 10654 4040
rect 10598 3984 10600 4004
rect 10600 3984 10652 4004
rect 10652 3984 10654 4004
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 12070 4528 12126 4584
rect 12530 4256 12586 4312
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12714 3440 12770 3496
rect 13542 7828 13544 7848
rect 13544 7828 13596 7848
rect 13596 7828 13598 7848
rect 13542 7792 13598 7828
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 13634 3576 13690 3632
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14646 10140 14648 10160
rect 14648 10140 14700 10160
rect 14700 10140 14702 10160
rect 14646 10104 14702 10140
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 15934 10104 15990 10160
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14646 7928 14702 7984
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14554 6604 14556 6624
rect 14556 6604 14608 6624
rect 14608 6604 14610 6624
rect 14554 6568 14610 6604
rect 14554 5752 14610 5808
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 15290 6432 15346 6488
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14462 3984 14518 4040
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 15566 2796 15568 2816
rect 15568 2796 15620 2816
rect 15620 2796 15622 2816
rect 15566 2760 15622 2796
rect 16394 7928 16450 7984
rect 15842 3032 15898 3088
rect 16210 4664 16266 4720
rect 16026 4256 16082 4312
rect 16486 5908 16542 5944
rect 16486 5888 16488 5908
rect 16488 5888 16540 5908
rect 16540 5888 16542 5908
rect 16486 5616 16542 5672
rect 16578 5208 16634 5264
rect 18970 21256 19026 21312
rect 19522 20848 19578 20904
rect 21546 22208 21602 22264
rect 20810 20324 20866 20360
rect 20810 20304 20812 20324
rect 20812 20304 20864 20324
rect 20864 20304 20866 20324
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 20810 19916 20866 19952
rect 20810 19896 20812 19916
rect 20812 19896 20864 19916
rect 20864 19896 20866 19916
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 17222 7928 17278 7984
rect 16578 4936 16634 4992
rect 17130 6432 17186 6488
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 17958 9696 18014 9752
rect 17774 9288 17830 9344
rect 17682 7792 17738 7848
rect 17406 6568 17462 6624
rect 17682 6296 17738 6352
rect 17498 5072 17554 5128
rect 17038 2896 17094 2952
rect 17958 8880 18014 8936
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18694 11192 18750 11248
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18878 12552 18934 12608
rect 19062 12008 19118 12064
rect 19154 11600 19210 11656
rect 18142 10240 18198 10296
rect 18326 9968 18382 10024
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18142 9696 18198 9752
rect 18694 9832 18750 9888
rect 18694 9696 18750 9752
rect 18786 9560 18842 9616
rect 17958 6024 18014 6080
rect 17958 5616 18014 5672
rect 17958 5208 18014 5264
rect 17958 4664 18014 4720
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18142 6976 18198 7032
rect 18970 10648 19026 10704
rect 18786 8336 18842 8392
rect 18786 7828 18788 7848
rect 18788 7828 18840 7848
rect 18840 7828 18842 7848
rect 18786 7792 18842 7828
rect 18694 7520 18750 7576
rect 18602 6704 18658 6760
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18694 6568 18750 6624
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 19338 5344 19394 5400
rect 18602 4800 18658 4856
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 17958 3576 18014 3632
rect 17958 2896 18014 2952
rect 17958 2352 18014 2408
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18694 3304 18750 3360
rect 18602 2896 18658 2952
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19246 4936 19302 4992
rect 19154 4820 19210 4856
rect 19154 4800 19156 4820
rect 19156 4800 19208 4820
rect 19208 4800 19210 4820
rect 19062 1944 19118 2000
rect 19154 1536 19210 1592
rect 19430 4120 19486 4176
rect 20810 17196 20866 17232
rect 20810 17176 20812 17196
rect 20812 17176 20864 17196
rect 20864 17176 20866 17196
rect 20810 15680 20866 15736
rect 19890 6160 19946 6216
rect 20074 5752 20130 5808
rect 19798 3712 19854 3768
rect 21362 19352 21418 19408
rect 21362 18944 21418 19000
rect 21362 18536 21418 18592
rect 21362 17992 21418 18048
rect 21362 17604 21418 17640
rect 21362 17584 21364 17604
rect 21364 17584 21416 17604
rect 21416 17584 21418 17604
rect 21454 16632 21510 16688
rect 21362 16224 21418 16280
rect 21362 15272 21418 15328
rect 21270 14864 21326 14920
rect 21454 14320 21510 14376
rect 21362 13912 21418 13968
rect 21362 13504 21418 13560
rect 20074 3712 20130 3768
rect 20718 5072 20774 5128
rect 20258 3984 20314 4040
rect 20258 3188 20314 3224
rect 20258 3168 20260 3188
rect 20260 3168 20312 3188
rect 20312 3168 20314 3188
rect 20534 4120 20590 4176
rect 20534 3712 20590 3768
rect 20350 992 20406 1048
rect 21270 12980 21326 13016
rect 21270 12960 21272 12980
rect 21272 12960 21324 12980
rect 21324 12960 21326 12980
rect 21178 5888 21234 5944
rect 22006 5344 22062 5400
rect 21086 2760 21142 2816
rect 20534 584 20590 640
rect 21270 176 21326 232
<< metal3 >>
rect 20621 22674 20687 22677
rect 22200 22674 23000 22704
rect 20621 22672 23000 22674
rect 20621 22616 20626 22672
rect 20682 22616 23000 22672
rect 20621 22614 23000 22616
rect 20621 22611 20687 22614
rect 22200 22584 23000 22614
rect 21541 22266 21607 22269
rect 22200 22266 23000 22296
rect 21541 22264 23000 22266
rect 21541 22208 21546 22264
rect 21602 22208 23000 22264
rect 21541 22206 23000 22208
rect 21541 22203 21607 22206
rect 22200 22176 23000 22206
rect 18597 21722 18663 21725
rect 22200 21722 23000 21752
rect 18597 21720 23000 21722
rect 18597 21664 18602 21720
rect 18658 21664 23000 21720
rect 18597 21662 23000 21664
rect 18597 21659 18663 21662
rect 22200 21632 23000 21662
rect 18965 21314 19031 21317
rect 22200 21314 23000 21344
rect 18965 21312 23000 21314
rect 18965 21256 18970 21312
rect 19026 21256 23000 21312
rect 18965 21254 23000 21256
rect 18965 21251 19031 21254
rect 22200 21224 23000 21254
rect 19517 20906 19583 20909
rect 22200 20906 23000 20936
rect 19517 20904 23000 20906
rect 19517 20848 19522 20904
rect 19578 20848 23000 20904
rect 19517 20846 23000 20848
rect 19517 20843 19583 20846
rect 22200 20816 23000 20846
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 20805 20362 20871 20365
rect 22200 20362 23000 20392
rect 20805 20360 23000 20362
rect 20805 20304 20810 20360
rect 20866 20304 23000 20360
rect 20805 20302 23000 20304
rect 20805 20299 20871 20302
rect 22200 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 20805 19954 20871 19957
rect 22200 19954 23000 19984
rect 20805 19952 23000 19954
rect 20805 19896 20810 19952
rect 20866 19896 23000 19952
rect 20805 19894 23000 19896
rect 20805 19891 20871 19894
rect 22200 19864 23000 19894
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 21357 19410 21423 19413
rect 22200 19410 23000 19440
rect 21357 19408 23000 19410
rect 21357 19352 21362 19408
rect 21418 19352 23000 19408
rect 21357 19350 23000 19352
rect 21357 19347 21423 19350
rect 22200 19320 23000 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 21357 19002 21423 19005
rect 22200 19002 23000 19032
rect 21357 19000 23000 19002
rect 21357 18944 21362 19000
rect 21418 18944 23000 19000
rect 21357 18942 23000 18944
rect 21357 18939 21423 18942
rect 22200 18912 23000 18942
rect 21357 18594 21423 18597
rect 22200 18594 23000 18624
rect 21357 18592 23000 18594
rect 21357 18536 21362 18592
rect 21418 18536 23000 18592
rect 21357 18534 23000 18536
rect 21357 18531 21423 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 22200 18504 23000 18534
rect 18270 18463 18590 18464
rect 21357 18050 21423 18053
rect 22200 18050 23000 18080
rect 21357 18048 23000 18050
rect 21357 17992 21362 18048
rect 21418 17992 23000 18048
rect 21357 17990 23000 17992
rect 21357 17987 21423 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 21357 17642 21423 17645
rect 22200 17642 23000 17672
rect 21357 17640 23000 17642
rect 21357 17584 21362 17640
rect 21418 17584 23000 17640
rect 21357 17582 23000 17584
rect 21357 17579 21423 17582
rect 22200 17552 23000 17582
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 20805 17234 20871 17237
rect 22200 17234 23000 17264
rect 20805 17232 23000 17234
rect 20805 17176 20810 17232
rect 20866 17176 23000 17232
rect 20805 17174 23000 17176
rect 20805 17171 20871 17174
rect 22200 17144 23000 17174
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 21449 16690 21515 16693
rect 22200 16690 23000 16720
rect 21449 16688 23000 16690
rect 21449 16632 21454 16688
rect 21510 16632 23000 16688
rect 21449 16630 23000 16632
rect 21449 16627 21515 16630
rect 22200 16600 23000 16630
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 21357 16282 21423 16285
rect 22200 16282 23000 16312
rect 21357 16280 23000 16282
rect 21357 16224 21362 16280
rect 21418 16224 23000 16280
rect 21357 16222 23000 16224
rect 21357 16219 21423 16222
rect 22200 16192 23000 16222
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 20805 15738 20871 15741
rect 22200 15738 23000 15768
rect 20805 15736 23000 15738
rect 20805 15680 20810 15736
rect 20866 15680 23000 15736
rect 20805 15678 23000 15680
rect 20805 15675 20871 15678
rect 22200 15648 23000 15678
rect 21357 15330 21423 15333
rect 22200 15330 23000 15360
rect 21357 15328 23000 15330
rect 21357 15272 21362 15328
rect 21418 15272 23000 15328
rect 21357 15270 23000 15272
rect 21357 15267 21423 15270
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 22200 15240 23000 15270
rect 18270 15199 18590 15200
rect 21265 14922 21331 14925
rect 22200 14922 23000 14952
rect 21265 14920 23000 14922
rect 21265 14864 21270 14920
rect 21326 14864 23000 14920
rect 21265 14862 23000 14864
rect 21265 14859 21331 14862
rect 22200 14832 23000 14862
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 21449 14378 21515 14381
rect 22200 14378 23000 14408
rect 21449 14376 23000 14378
rect 21449 14320 21454 14376
rect 21510 14320 23000 14376
rect 21449 14318 23000 14320
rect 21449 14315 21515 14318
rect 22200 14288 23000 14318
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 21357 13970 21423 13973
rect 22200 13970 23000 14000
rect 21357 13968 23000 13970
rect 21357 13912 21362 13968
rect 21418 13912 23000 13968
rect 21357 13910 23000 13912
rect 21357 13907 21423 13910
rect 22200 13880 23000 13910
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 21357 13562 21423 13565
rect 22200 13562 23000 13592
rect 21357 13560 23000 13562
rect 21357 13504 21362 13560
rect 21418 13504 23000 13560
rect 21357 13502 23000 13504
rect 21357 13499 21423 13502
rect 22200 13472 23000 13502
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 21265 13018 21331 13021
rect 22200 13018 23000 13048
rect 21265 13016 23000 13018
rect 21265 12960 21270 13016
rect 21326 12960 23000 13016
rect 21265 12958 23000 12960
rect 21265 12955 21331 12958
rect 22200 12928 23000 12958
rect 18873 12610 18939 12613
rect 22200 12610 23000 12640
rect 18873 12608 23000 12610
rect 18873 12552 18878 12608
rect 18934 12552 23000 12608
rect 18873 12550 23000 12552
rect 18873 12547 18939 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 22200 12520 23000 12550
rect 14805 12479 15125 12480
rect 19057 12066 19123 12069
rect 22200 12066 23000 12096
rect 19057 12064 23000 12066
rect 19057 12008 19062 12064
rect 19118 12008 23000 12064
rect 19057 12006 23000 12008
rect 19057 12003 19123 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 22200 11976 23000 12006
rect 18270 11935 18590 11936
rect 19149 11658 19215 11661
rect 22200 11658 23000 11688
rect 19149 11656 23000 11658
rect 19149 11600 19154 11656
rect 19210 11600 23000 11656
rect 19149 11598 23000 11600
rect 19149 11595 19215 11598
rect 22200 11568 23000 11598
rect 0 11522 800 11552
rect 1669 11522 1735 11525
rect 0 11520 1735 11522
rect 0 11464 1674 11520
rect 1730 11464 1735 11520
rect 0 11462 1735 11464
rect 0 11432 800 11462
rect 1669 11459 1735 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 18689 11250 18755 11253
rect 22200 11250 23000 11280
rect 18689 11248 23000 11250
rect 18689 11192 18694 11248
rect 18750 11192 23000 11248
rect 18689 11190 23000 11192
rect 18689 11187 18755 11190
rect 22200 11160 23000 11190
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 18965 10706 19031 10709
rect 22200 10706 23000 10736
rect 18965 10704 23000 10706
rect 18965 10648 18970 10704
rect 19026 10648 23000 10704
rect 18965 10646 23000 10648
rect 18965 10643 19031 10646
rect 22200 10616 23000 10646
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 18137 10298 18203 10301
rect 22200 10298 23000 10328
rect 18137 10296 23000 10298
rect 18137 10240 18142 10296
rect 18198 10240 23000 10296
rect 18137 10238 23000 10240
rect 18137 10235 18203 10238
rect 22200 10208 23000 10238
rect 14641 10162 14707 10165
rect 15929 10162 15995 10165
rect 14641 10160 19350 10162
rect 14641 10104 14646 10160
rect 14702 10104 15934 10160
rect 15990 10104 19350 10160
rect 14641 10102 19350 10104
rect 14641 10099 14707 10102
rect 15929 10099 15995 10102
rect 18321 10026 18387 10029
rect 18140 10024 18387 10026
rect 18140 9968 18326 10024
rect 18382 9968 18387 10024
rect 18140 9966 18387 9968
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18140 9757 18200 9966
rect 18321 9963 18387 9966
rect 18689 9888 18755 9893
rect 18689 9832 18694 9888
rect 18750 9832 18755 9888
rect 18689 9827 18755 9832
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 18692 9757 18752 9827
rect 17953 9752 18019 9757
rect 17953 9696 17958 9752
rect 18014 9696 18019 9752
rect 17953 9691 18019 9696
rect 18137 9752 18203 9757
rect 18137 9696 18142 9752
rect 18198 9696 18203 9752
rect 18137 9691 18203 9696
rect 18689 9752 18755 9757
rect 18689 9696 18694 9752
rect 18750 9696 18755 9752
rect 18689 9691 18755 9696
rect 19290 9754 19350 10102
rect 22200 9754 23000 9784
rect 19290 9694 23000 9754
rect 17956 9618 18016 9691
rect 22200 9664 23000 9694
rect 18781 9618 18847 9621
rect 17956 9616 18847 9618
rect 17956 9560 18786 9616
rect 18842 9560 18847 9616
rect 17956 9558 18847 9560
rect 18781 9555 18847 9558
rect 17769 9346 17835 9349
rect 22200 9346 23000 9376
rect 17769 9344 23000 9346
rect 17769 9288 17774 9344
rect 17830 9288 23000 9344
rect 17769 9286 23000 9288
rect 17769 9283 17835 9286
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 22200 9256 23000 9286
rect 14805 9215 15125 9216
rect 17953 8938 18019 8941
rect 22200 8938 23000 8968
rect 17953 8936 23000 8938
rect 17953 8880 17958 8936
rect 18014 8880 23000 8936
rect 17953 8878 23000 8880
rect 17953 8875 18019 8878
rect 22200 8848 23000 8878
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 18781 8394 18847 8397
rect 22200 8394 23000 8424
rect 18781 8392 23000 8394
rect 18781 8336 18786 8392
rect 18842 8336 23000 8392
rect 18781 8334 23000 8336
rect 18781 8331 18847 8334
rect 22200 8304 23000 8334
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 14641 7986 14707 7989
rect 16389 7986 16455 7989
rect 14641 7984 16455 7986
rect 14641 7928 14646 7984
rect 14702 7928 16394 7984
rect 16450 7928 16455 7984
rect 14641 7926 16455 7928
rect 14641 7923 14707 7926
rect 16389 7923 16455 7926
rect 17217 7986 17283 7989
rect 22200 7986 23000 8016
rect 17217 7984 23000 7986
rect 17217 7928 17222 7984
rect 17278 7928 23000 7984
rect 17217 7926 23000 7928
rect 17217 7923 17283 7926
rect 22200 7896 23000 7926
rect 13537 7850 13603 7853
rect 17677 7850 17743 7853
rect 18781 7850 18847 7853
rect 13537 7848 18847 7850
rect 13537 7792 13542 7848
rect 13598 7792 17682 7848
rect 17738 7792 18786 7848
rect 18842 7792 18847 7848
rect 13537 7790 18847 7792
rect 13537 7787 13603 7790
rect 17677 7787 17743 7790
rect 18781 7787 18847 7790
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 18689 7578 18755 7581
rect 22200 7578 23000 7608
rect 18689 7576 23000 7578
rect 18689 7520 18694 7576
rect 18750 7520 23000 7576
rect 18689 7518 23000 7520
rect 18689 7515 18755 7518
rect 22200 7488 23000 7518
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 18137 7034 18203 7037
rect 22200 7034 23000 7064
rect 18137 7032 23000 7034
rect 18137 6976 18142 7032
rect 18198 6976 23000 7032
rect 18137 6974 23000 6976
rect 18137 6971 18203 6974
rect 22200 6944 23000 6974
rect 9489 6898 9555 6901
rect 18822 6898 18828 6900
rect 9489 6896 18828 6898
rect 9489 6840 9494 6896
rect 9550 6840 18828 6896
rect 9489 6838 18828 6840
rect 9489 6835 9555 6838
rect 18822 6836 18828 6838
rect 18892 6836 18898 6900
rect 11697 6762 11763 6765
rect 18597 6762 18663 6765
rect 11697 6760 18663 6762
rect 11697 6704 11702 6760
rect 11758 6704 18602 6760
rect 18658 6704 18663 6760
rect 11697 6702 18663 6704
rect 11697 6699 11763 6702
rect 18597 6699 18663 6702
rect 14549 6626 14615 6629
rect 17401 6626 17467 6629
rect 14549 6624 17467 6626
rect 14549 6568 14554 6624
rect 14610 6568 17406 6624
rect 17462 6568 17467 6624
rect 14549 6566 17467 6568
rect 14549 6563 14615 6566
rect 17401 6563 17467 6566
rect 18689 6626 18755 6629
rect 22200 6626 23000 6656
rect 18689 6624 23000 6626
rect 18689 6568 18694 6624
rect 18750 6568 23000 6624
rect 18689 6566 23000 6568
rect 18689 6563 18755 6566
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 22200 6536 23000 6566
rect 18270 6495 18590 6496
rect 15285 6490 15351 6493
rect 17125 6490 17191 6493
rect 15285 6488 17191 6490
rect 15285 6432 15290 6488
rect 15346 6432 17130 6488
rect 17186 6432 17191 6488
rect 15285 6430 17191 6432
rect 15285 6427 15351 6430
rect 17125 6427 17191 6430
rect 10869 6354 10935 6357
rect 17677 6354 17743 6357
rect 10869 6352 17743 6354
rect 10869 6296 10874 6352
rect 10930 6296 17682 6352
rect 17738 6296 17743 6352
rect 10869 6294 17743 6296
rect 10869 6291 10935 6294
rect 17677 6291 17743 6294
rect 10869 6218 10935 6221
rect 19885 6218 19951 6221
rect 10869 6216 19951 6218
rect 10869 6160 10874 6216
rect 10930 6160 19890 6216
rect 19946 6160 19951 6216
rect 10869 6158 19951 6160
rect 10869 6155 10935 6158
rect 19885 6155 19951 6158
rect 17953 6082 18019 6085
rect 22200 6082 23000 6112
rect 17953 6080 23000 6082
rect 17953 6024 17958 6080
rect 18014 6024 23000 6080
rect 17953 6022 23000 6024
rect 17953 6019 18019 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 22200 5992 23000 6022
rect 14805 5951 15125 5952
rect 16481 5946 16547 5949
rect 21173 5946 21239 5949
rect 15702 5944 21239 5946
rect 15702 5888 16486 5944
rect 16542 5888 21178 5944
rect 21234 5888 21239 5944
rect 15702 5886 21239 5888
rect 14549 5810 14615 5813
rect 15702 5810 15762 5886
rect 16481 5883 16547 5886
rect 21173 5883 21239 5886
rect 14549 5808 15762 5810
rect 14549 5752 14554 5808
rect 14610 5752 15762 5808
rect 14549 5750 15762 5752
rect 20069 5810 20135 5813
rect 20478 5810 20484 5812
rect 20069 5808 20484 5810
rect 20069 5752 20074 5808
rect 20130 5752 20484 5808
rect 20069 5750 20484 5752
rect 14549 5747 14615 5750
rect 20069 5747 20135 5750
rect 20478 5748 20484 5750
rect 20548 5748 20554 5812
rect 9673 5674 9739 5677
rect 16481 5674 16547 5677
rect 9673 5672 16547 5674
rect 9673 5616 9678 5672
rect 9734 5616 16486 5672
rect 16542 5616 16547 5672
rect 9673 5614 16547 5616
rect 9673 5611 9739 5614
rect 16481 5611 16547 5614
rect 17953 5674 18019 5677
rect 22200 5674 23000 5704
rect 17953 5672 23000 5674
rect 17953 5616 17958 5672
rect 18014 5616 23000 5672
rect 17953 5614 23000 5616
rect 17953 5611 18019 5614
rect 22200 5584 23000 5614
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 8201 5402 8267 5405
rect 9857 5402 9923 5405
rect 8201 5400 9923 5402
rect 8201 5344 8206 5400
rect 8262 5344 9862 5400
rect 9918 5344 9923 5400
rect 8201 5342 9923 5344
rect 8201 5339 8267 5342
rect 9857 5339 9923 5342
rect 19333 5402 19399 5405
rect 22001 5402 22067 5405
rect 19333 5400 22067 5402
rect 19333 5344 19338 5400
rect 19394 5344 22006 5400
rect 22062 5344 22067 5400
rect 19333 5342 22067 5344
rect 19333 5339 19399 5342
rect 22001 5339 22067 5342
rect 9857 5266 9923 5269
rect 16573 5266 16639 5269
rect 9630 5264 16639 5266
rect 9630 5208 9862 5264
rect 9918 5208 16578 5264
rect 16634 5208 16639 5264
rect 9630 5206 16639 5208
rect 7281 5130 7347 5133
rect 9630 5130 9690 5206
rect 9857 5203 9923 5206
rect 16573 5203 16639 5206
rect 17953 5266 18019 5269
rect 22200 5266 23000 5296
rect 17953 5264 23000 5266
rect 17953 5208 17958 5264
rect 18014 5208 23000 5264
rect 17953 5206 23000 5208
rect 17953 5203 18019 5206
rect 22200 5176 23000 5206
rect 7281 5128 9690 5130
rect 7281 5072 7286 5128
rect 7342 5072 9690 5128
rect 7281 5070 9690 5072
rect 17493 5130 17559 5133
rect 20713 5130 20779 5133
rect 17493 5128 20779 5130
rect 17493 5072 17498 5128
rect 17554 5072 20718 5128
rect 20774 5072 20779 5128
rect 17493 5070 20779 5072
rect 7281 5067 7347 5070
rect 17493 5067 17559 5070
rect 20713 5067 20779 5070
rect 16573 4994 16639 4997
rect 19241 4994 19307 4997
rect 16573 4992 19307 4994
rect 16573 4936 16578 4992
rect 16634 4936 19246 4992
rect 19302 4936 19307 4992
rect 16573 4934 19307 4936
rect 16573 4931 16639 4934
rect 19241 4931 19307 4934
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 18597 4858 18663 4861
rect 19149 4858 19215 4861
rect 18597 4856 19215 4858
rect 18597 4800 18602 4856
rect 18658 4800 19154 4856
rect 19210 4800 19215 4856
rect 18597 4798 19215 4800
rect 18597 4795 18663 4798
rect 19149 4795 19215 4798
rect 9489 4722 9555 4725
rect 16205 4722 16271 4725
rect 9489 4720 16271 4722
rect 9489 4664 9494 4720
rect 9550 4664 16210 4720
rect 16266 4664 16271 4720
rect 9489 4662 16271 4664
rect 9489 4659 9555 4662
rect 16205 4659 16271 4662
rect 17953 4722 18019 4725
rect 22200 4722 23000 4752
rect 17953 4720 23000 4722
rect 17953 4664 17958 4720
rect 18014 4664 23000 4720
rect 17953 4662 23000 4664
rect 17953 4659 18019 4662
rect 22200 4632 23000 4662
rect 9213 4586 9279 4589
rect 10133 4586 10199 4589
rect 9213 4584 10199 4586
rect 9213 4528 9218 4584
rect 9274 4528 10138 4584
rect 10194 4528 10199 4584
rect 9213 4526 10199 4528
rect 9213 4523 9279 4526
rect 10133 4523 10199 4526
rect 12065 4586 12131 4589
rect 12065 4584 19350 4586
rect 12065 4528 12070 4584
rect 12126 4528 19350 4584
rect 12065 4526 19350 4528
rect 12065 4523 12131 4526
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 12525 4314 12591 4317
rect 16021 4314 16087 4317
rect 12525 4312 16087 4314
rect 12525 4256 12530 4312
rect 12586 4256 16026 4312
rect 16082 4256 16087 4312
rect 12525 4254 16087 4256
rect 19290 4314 19350 4526
rect 22200 4314 23000 4344
rect 19290 4254 23000 4314
rect 12525 4251 12591 4254
rect 16021 4251 16087 4254
rect 22200 4224 23000 4254
rect 10133 4178 10199 4181
rect 19425 4178 19491 4181
rect 20529 4178 20595 4181
rect 10133 4176 19350 4178
rect 10133 4120 10138 4176
rect 10194 4120 19350 4176
rect 10133 4118 19350 4120
rect 10133 4115 10199 4118
rect 7005 4042 7071 4045
rect 10593 4042 10659 4045
rect 14457 4042 14523 4045
rect 7005 4040 8402 4042
rect 7005 3984 7010 4040
rect 7066 3984 8402 4040
rect 7005 3982 8402 3984
rect 7005 3979 7071 3982
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 8342 3770 8402 3982
rect 10593 4040 14523 4042
rect 10593 3984 10598 4040
rect 10654 3984 14462 4040
rect 14518 3984 14523 4040
rect 10593 3982 14523 3984
rect 10593 3979 10659 3982
rect 14457 3979 14523 3982
rect 19290 3906 19350 4118
rect 19425 4176 20595 4178
rect 19425 4120 19430 4176
rect 19486 4120 20534 4176
rect 20590 4120 20595 4176
rect 19425 4118 20595 4120
rect 19425 4115 19491 4118
rect 20529 4115 20595 4118
rect 20253 4044 20319 4045
rect 20253 4040 20300 4044
rect 20364 4042 20370 4044
rect 20253 3984 20258 4040
rect 20253 3980 20300 3984
rect 20364 3982 20410 4042
rect 20364 3980 20370 3982
rect 20253 3979 20319 3980
rect 22200 3906 23000 3936
rect 19290 3846 23000 3906
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 19793 3770 19859 3773
rect 20069 3770 20135 3773
rect 20529 3772 20595 3773
rect 8342 3710 14658 3770
rect 6085 3634 6151 3637
rect 13629 3634 13695 3637
rect 6085 3632 13695 3634
rect 6085 3576 6090 3632
rect 6146 3576 13634 3632
rect 13690 3576 13695 3632
rect 6085 3574 13695 3576
rect 14598 3634 14658 3710
rect 19793 3768 20135 3770
rect 19793 3712 19798 3768
rect 19854 3712 20074 3768
rect 20130 3712 20135 3768
rect 19793 3710 20135 3712
rect 19793 3707 19859 3710
rect 20069 3707 20135 3710
rect 20478 3708 20484 3772
rect 20548 3770 20595 3772
rect 20548 3768 20640 3770
rect 20590 3712 20640 3768
rect 20548 3710 20640 3712
rect 20548 3708 20595 3710
rect 20529 3707 20595 3708
rect 17953 3634 18019 3637
rect 14598 3632 18019 3634
rect 14598 3576 17958 3632
rect 18014 3576 18019 3632
rect 14598 3574 18019 3576
rect 6085 3571 6151 3574
rect 13629 3571 13695 3574
rect 17953 3571 18019 3574
rect 4797 3498 4863 3501
rect 12709 3498 12775 3501
rect 4797 3496 12775 3498
rect 4797 3440 4802 3496
rect 4858 3440 12714 3496
rect 12770 3440 12775 3496
rect 4797 3438 12775 3440
rect 4797 3435 4863 3438
rect 12709 3435 12775 3438
rect 18689 3362 18755 3365
rect 22200 3362 23000 3392
rect 18689 3360 23000 3362
rect 18689 3304 18694 3360
rect 18750 3304 23000 3360
rect 18689 3302 23000 3304
rect 18689 3299 18755 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 22200 3272 23000 3302
rect 18270 3231 18590 3232
rect 7281 3226 7347 3229
rect 10133 3226 10199 3229
rect 20253 3228 20319 3229
rect 20253 3226 20300 3228
rect 7281 3224 10199 3226
rect 7281 3168 7286 3224
rect 7342 3168 10138 3224
rect 10194 3168 10199 3224
rect 7281 3166 10199 3168
rect 20208 3224 20300 3226
rect 20208 3168 20258 3224
rect 20208 3166 20300 3168
rect 7281 3163 7347 3166
rect 10133 3163 10199 3166
rect 20253 3164 20300 3166
rect 20364 3164 20370 3228
rect 20253 3163 20319 3164
rect 5625 3090 5691 3093
rect 15837 3090 15903 3093
rect 5625 3088 15903 3090
rect 5625 3032 5630 3088
rect 5686 3032 15842 3088
rect 15898 3032 15903 3088
rect 5625 3030 15903 3032
rect 5625 3027 5691 3030
rect 15837 3027 15903 3030
rect 1577 2954 1643 2957
rect 17033 2954 17099 2957
rect 1577 2952 17099 2954
rect 1577 2896 1582 2952
rect 1638 2896 17038 2952
rect 17094 2896 17099 2952
rect 1577 2894 17099 2896
rect 1577 2891 1643 2894
rect 17033 2891 17099 2894
rect 17953 2954 18019 2957
rect 18597 2954 18663 2957
rect 17953 2952 18663 2954
rect 17953 2896 17958 2952
rect 18014 2896 18602 2952
rect 18658 2896 18663 2952
rect 17953 2894 18663 2896
rect 17953 2891 18019 2894
rect 18597 2891 18663 2894
rect 18822 2892 18828 2956
rect 18892 2954 18898 2956
rect 22200 2954 23000 2984
rect 18892 2894 23000 2954
rect 18892 2892 18898 2894
rect 22200 2864 23000 2894
rect 15561 2818 15627 2821
rect 21081 2818 21147 2821
rect 15561 2816 21147 2818
rect 15561 2760 15566 2816
rect 15622 2760 21086 2816
rect 21142 2760 21147 2816
rect 15561 2758 21147 2760
rect 15561 2755 15627 2758
rect 21081 2755 21147 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 5533 2546 5599 2549
rect 8661 2546 8727 2549
rect 5533 2544 8727 2546
rect 5533 2488 5538 2544
rect 5594 2488 8666 2544
rect 8722 2488 8727 2544
rect 5533 2486 8727 2488
rect 5533 2483 5599 2486
rect 8661 2483 8727 2486
rect 5165 2410 5231 2413
rect 9305 2410 9371 2413
rect 5165 2408 9371 2410
rect 5165 2352 5170 2408
rect 5226 2352 9310 2408
rect 9366 2352 9371 2408
rect 5165 2350 9371 2352
rect 5165 2347 5231 2350
rect 9305 2347 9371 2350
rect 17953 2410 18019 2413
rect 22200 2410 23000 2440
rect 17953 2408 23000 2410
rect 17953 2352 17958 2408
rect 18014 2352 23000 2408
rect 17953 2350 23000 2352
rect 17953 2347 18019 2350
rect 22200 2320 23000 2350
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 19057 2002 19123 2005
rect 22200 2002 23000 2032
rect 19057 2000 23000 2002
rect 19057 1944 19062 2000
rect 19118 1944 23000 2000
rect 19057 1942 23000 1944
rect 19057 1939 19123 1942
rect 22200 1912 23000 1942
rect 19149 1594 19215 1597
rect 22200 1594 23000 1624
rect 19149 1592 23000 1594
rect 19149 1536 19154 1592
rect 19210 1536 23000 1592
rect 19149 1534 23000 1536
rect 19149 1531 19215 1534
rect 22200 1504 23000 1534
rect 20345 1050 20411 1053
rect 22200 1050 23000 1080
rect 20345 1048 23000 1050
rect 20345 992 20350 1048
rect 20406 992 23000 1048
rect 20345 990 23000 992
rect 20345 987 20411 990
rect 22200 960 23000 990
rect 20529 642 20595 645
rect 22200 642 23000 672
rect 20529 640 23000 642
rect 20529 584 20534 640
rect 20590 584 23000 640
rect 20529 582 23000 584
rect 20529 579 20595 582
rect 22200 552 23000 582
rect 21265 234 21331 237
rect 22200 234 23000 264
rect 21265 232 23000 234
rect 21265 176 21270 232
rect 21326 176 23000 232
rect 21265 174 23000 176
rect 21265 171 21331 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 18828 6836 18892 6900
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 20484 5748 20548 5812
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 20300 4040 20364 4044
rect 20300 3984 20314 4040
rect 20314 3984 20364 4040
rect 20300 3980 20364 3984
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 20484 3768 20548 3772
rect 20484 3712 20534 3768
rect 20534 3712 20548 3768
rect 20484 3708 20548 3712
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 20300 3224 20364 3228
rect 20300 3168 20314 3224
rect 20314 3168 20364 3224
rect 20300 3164 20364 3168
rect 18828 2892 18892 2956
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18827 6900 18893 6901
rect 18827 6836 18828 6900
rect 18892 6836 18893 6900
rect 18827 6835 18893 6836
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18830 2957 18890 6835
rect 20483 5812 20549 5813
rect 20483 5748 20484 5812
rect 20548 5748 20549 5812
rect 20483 5747 20549 5748
rect 20299 4044 20365 4045
rect 20299 3980 20300 4044
rect 20364 3980 20365 4044
rect 20299 3979 20365 3980
rect 20302 3229 20362 3979
rect 20486 3773 20546 5747
rect 20483 3772 20549 3773
rect 20483 3708 20484 3772
rect 20548 3708 20549 3772
rect 20483 3707 20549 3708
rect 20299 3228 20365 3229
rect 20299 3164 20300 3228
rect 20364 3164 20365 3228
rect 20299 3163 20365 3164
rect 18827 2956 18893 2957
rect 18827 2892 18828 2956
rect 18892 2892 18893 2956
rect 18827 2891 18893 2892
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_6
timestamp 1624635492
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_14
timestamp 1624635492
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_10
timestamp 1624635492
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14
timestamp 1624635492
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1624635492
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18
timestamp 1624635492
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1624635492
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1624635492
transform 1 0 2576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 3128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1624635492
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3312 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_28
timestamp 1624635492
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1624635492
transform 1 0 4048 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1624635492
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1624635492
transform -1 0 4324 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1624635492
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_36
timestamp 1624635492
transform 1 0 4416 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40
timestamp 1624635492
transform 1 0 4784 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1624635492
transform 1 0 4508 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1624635492
transform -1 0 4784 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1624635492
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1624635492
transform -1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46
timestamp 1624635492
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1624635492
transform 1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1624635492
transform 1 0 5520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_50
timestamp 1624635492
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51
timestamp 1624635492
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1624635492
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1624635492
transform -1 0 6256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55
timestamp 1624635492
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1624635492
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 6716 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_61
timestamp 1624635492
transform 1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1624635492
transform -1 0 6992 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8924 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1624635492
transform -1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1624635492
transform -1 0 7268 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64
timestamp 1624635492
transform 1 0 6992 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1624635492
transform 1 0 7452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73
timestamp 1624635492
transform 1 0 7820 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1624635492
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_67
timestamp 1624635492
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1624635492
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1624635492
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93
timestamp 1624635492
transform 1 0 9660 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624635492
transform -1 0 9660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _42_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 9108 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1624635492
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11224 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11224 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1624635492
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1624635492
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1624635492
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp 1624635492
transform 1 0 12236 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1624635492
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13340 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1624635492
transform -1 0 12328 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13892 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform -1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 14444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp 1624635492
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_139
timestamp 1624635492
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1624635492
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1624635492
transform 1 0 14444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1624635492
transform 1 0 15824 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1624635492
transform 1 0 15732 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1624635492
transform 1 0 14812 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15548 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_146
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1624635492
transform 1 0 15548 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp 1624635492
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1624635492
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1624635492
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_168
timestamp 1624635492
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_183
timestamp 1624635492
transform 1 0 17940 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 1624635492
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1624635492
transform -1 0 19136 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1624635492
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 20332 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1624635492
transform -1 0 19596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_195
timestamp 1624635492
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1624635492
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1624635492
transform 1 0 19136 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_215
timestamp 1624635492
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1624635492
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1624635492
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1624635492
transform -1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform -1 0 21436 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1624635492
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1624635492
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 20516 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_17
timestamp 1624635492
transform 1 0 2668 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 4508 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output53_A
timestamp 1624635492
transform -1 0 4140 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_33
timestamp 1624635492
transform 1 0 4140 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1624635492
transform 1 0 4508 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7176 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 6164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 5428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 1624635492
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_47
timestamp 1624635492
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1624635492
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1624635492
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8832 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1624635492
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11408 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1624635492
transform -1 0 9568 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1624635492
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1624635492
transform 1 0 9568 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1624635492
transform 1 0 11592 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 13524 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1624635492
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_117
timestamp 1624635492
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_135
timestamp 1624635492
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1624635492
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 16376 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_148
timestamp 1624635492
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1624635492
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18032 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1624635492
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 20056 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1624635492
transform -1 0 19228 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1624635492
transform 1 0 19228 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1624635492
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1624635492
transform -1 0 21436 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1624635492
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1624635492
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1624635492
transform 1 0 4324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_38
timestamp 1624635492
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp 1624635492
transform 1 0 4968 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1624635492
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp 1624635492
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1624635492
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 6716 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_61
timestamp 1624635492
transform 1 0 6716 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1624635492
transform 1 0 7360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1624635492
transform 1 0 6900 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1624635492
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1624635492
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11224 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1624635492
transform -1 0 10212 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1624635492
transform -1 0 9752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1624635492
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1624635492
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1624635492
transform -1 0 12144 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13340 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1624635492
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_120
timestamp 1624635492
transform 1 0 12144 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1624635492
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1624635492
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 16008 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 16560 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1624635492
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 19780 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform 1 0 17756 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform 1 0 17204 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_168
timestamp 1624635492
transform 1 0 16560 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1624635492
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_185
timestamp 1624635492
transform 1 0 18124 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20148 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_203
timestamp 1624635492
transform 1 0 19780 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1624635492
transform 1 0 21160 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_216
timestamp 1624635492
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1624635492
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_mem_bottom_track_1.prog_clk_A
timestamp 1624635492
transform -1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp 1624635492
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1624635492
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_47
timestamp 1624635492
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_51
timestamp 1624635492
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_55
timestamp 1624635492
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1624635492
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1624635492
transform -1 0 8372 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1624635492
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 7360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1624635492
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1624635492
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1624635492
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11408 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1624635492
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1624635492
transform 1 0 10120 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1624635492
transform 1 0 10488 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11592 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1624635492
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_123
timestamp 1624635492
transform 1 0 12420 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1624635492
transform 1 0 12788 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 1624635492
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1624635492
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1624635492
transform -1 0 16008 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 14904 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 16560 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1624635492
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_162
timestamp 1624635492
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 17112 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_168
timestamp 1624635492
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1624635492
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 1624635492
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1624635492
transform 1 0 19780 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_196
timestamp 1624635492
transform 1 0 19136 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 21160 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1624635492
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1624635492
transform 1 0 21160 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_222
timestamp 1624635492
transform 1 0 21528 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1624635492
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1624635492
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1624635492
transform 1 0 4692 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 6716 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1624635492
transform -1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47
timestamp 1624635492
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 1624635492
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1624635492
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_61
timestamp 1624635492
transform 1 0 6716 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8372 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9384 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_79
timestamp 1624635492
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9936 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1624635492
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1624635492
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1624635492
transform -1 0 12144 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13892 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1624635492
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_120
timestamp 1624635492
transform 1 0 12144 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1624635492
transform 1 0 14076 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1624635492
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1624635492
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1624635492
transform 1 0 15916 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1624635492
transform 1 0 16376 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1624635492
transform -1 0 15732 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1624635492
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_159
timestamp 1624635492
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1624635492
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform 1 0 17664 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform -1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1624635492
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1624635492
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1624635492
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 19136 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_190
timestamp 1624635492
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_196
timestamp 1624635492
transform 1 0 19136 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_200
timestamp 1624635492
transform 1 0 19504 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1624635492
transform 1 0 21160 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1624635492
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1624635492
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1624635492
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1624635492
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624635492
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1624635492
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 6900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1624635492
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6072 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1624635492
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1624635492
transform -1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7360 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1624635492
transform -1 0 8372 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1624635492
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_68
timestamp 1624635492
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1624635492
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_66
timestamp 1624635492
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_84
timestamp 1624635492
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1624635492
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1624635492
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1624635492
transform 1 0 9568 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1624635492
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_95
timestamp 1624635492
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1624635492
transform -1 0 10948 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9016 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11500 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1624635492
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1624635492
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 1624635492
transform 1 0 11500 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1624635492
transform -1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_124
timestamp 1624635492
transform 1 0 12512 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_119
timestamp 1624635492
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1624635492
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1624635492
transform -1 0 12144 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp 1624635492
transform -1 0 12512 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12328 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13524 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1624635492
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1624635492
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1624635492
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_138
timestamp 1624635492
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1624635492
transform -1 0 13984 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1624635492
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1624635492
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1624635492
transform -1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1624635492
transform -1 0 16652 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 16100 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15916 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_150
timestamp 1624635492
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1624635492
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_163
timestamp 1624635492
transform 1 0 16100 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17112 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1624635492
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_183
timestamp 1624635492
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_187
timestamp 1624635492
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1624635492
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_190
timestamp 1624635492
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 19320 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1624635492
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_204
timestamp 1624635492
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_198
timestamp 1624635492
transform 1 0 19320 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20056 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 18768 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1624635492
transform 1 0 20424 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 21436 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1624635492
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1624635492
transform 1 0 21436 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1624635492
transform 1 0 21252 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1624635492
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1624635492
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1624635492
transform -1 0 8832 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_66
timestamp 1624635492
transform 1 0 7176 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_72
timestamp 1624635492
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp 1624635492
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1624635492
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9292 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1624635492
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1624635492
transform -1 0 12880 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1624635492
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1624635492
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1624635492
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139
timestamp 1624635492
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1624635492
transform -1 0 15088 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_147
timestamp 1624635492
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_152
timestamp 1624635492
transform 1 0 15088 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17848 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 17572 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1624635492
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_179
timestamp 1624635492
transform 1 0 17572 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19872 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1624635492
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_220
timestamp 1624635492
transform 1 0 21344 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1624635492
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9568 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_70
timestamp 1624635492
transform 1 0 7544 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_78
timestamp 1624635492
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_81
timestamp 1624635492
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11408 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1624635492
transform -1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1624635492
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1624635492
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1624635492
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1624635492
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 14720 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_126
timestamp 1624635492
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_130
timestamp 1624635492
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1624635492
transform -1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 16560 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_148
timestamp 1624635492
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1624635492
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1624635492
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1624635492
transform 1 0 18124 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17940 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_168
timestamp 1624635492
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_183
timestamp 1624635492
transform 1 0 17940 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1624635492
transform -1 0 19412 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1624635492
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_199
timestamp 1624635492
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1624635492
transform 1 0 20792 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_210
timestamp 1624635492
transform 1 0 20424 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1624635492
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1624635492
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1624635492
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1624635492
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1624635492
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1624635492
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_78
timestamp 1624635492
transform 1 0 8280 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1624635492
transform -1 0 9568 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11316 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1624635492
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_92
timestamp 1624635492
transform 1 0 9568 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_96
timestamp 1624635492
transform 1 0 9936 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 1624635492
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11592 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_111
timestamp 1624635492
transform 1 0 11316 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14076 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1624635492
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1624635492
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14536 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16376 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_155
timestamp 1624635492
transform 1 0 15364 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_166
timestamp 1624635492
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18032 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1624635492
transform 1 0 18216 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1624635492
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1624635492
transform 1 0 19872 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_195
timestamp 1624635492
transform 1 0 19044 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_199
timestamp 1624635492
transform 1 0 19412 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1624635492
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20332 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1624635492
transform 1 0 21160 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1624635492
transform 1 0 21528 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1624635492
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1624635492
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1624635492
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1624635492
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9568 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_70
timestamp 1624635492
transform 1 0 7544 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9752 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1624635492
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1624635492
transform -1 0 12144 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12328 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_110
timestamp 1624635492
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1624635492
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_124
timestamp 1624635492
transform 1 0 12512 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12696 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 16192 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1624635492
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1624635492
transform -1 0 16652 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_164
timestamp 1624635492
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18308 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1624635492
transform -1 0 17940 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1624635492
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_183
timestamp 1624635492
transform 1 0 17940 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19320 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1624635492
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1624635492
transform 1 0 20976 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_214
timestamp 1624635492
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1624635492
transform 1 0 21252 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1624635492
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1624635492
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1624635492
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1624635492
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1624635492
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10304 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10120 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_98
timestamp 1624635492
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11960 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_116
timestamp 1624635492
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1624635492
transform -1 0 14076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_134
timestamp 1624635492
transform 1 0 13432 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1624635492
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14536 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 16192 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_162
timestamp 1624635492
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1624635492
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_180
timestamp 1624635492
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1624635492
transform 1 0 18124 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1624635492
transform 1 0 18952 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1624635492
transform 1 0 18492 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 21436 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_192
timestamp 1624635492
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1624635492
transform 1 0 19228 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1624635492
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1624635492
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1624635492
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1624635492
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1624635492
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1624635492
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1624635492
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1624635492
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1624635492
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1624635492
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1624635492
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1624635492
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1624635492
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 1624635492
transform 1 0 11316 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1624635492
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_106
timestamp 1624635492
transform 1 0 10856 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 11408 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1624635492
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1624635492
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1624635492
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1624635492
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1624635492
transform -1 0 13064 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1624635492
transform 1 0 12880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1624635492
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_131
timestamp 1624635492
transform 1 0 13156 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1624635492
transform -1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_135
timestamp 1624635492
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1624635492
transform 1 0 13708 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1624635492
transform 1 0 13708 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_140
timestamp 1624635492
transform 1 0 13984 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1624635492
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1624635492
transform -1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14996 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14536 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16652 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15640 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_149
timestamp 1624635492
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1624635492
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_158
timestamp 1624635492
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18308 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17480 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_167
timestamp 1624635492
transform 1 0 16468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1624635492
transform 1 0 17112 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_187
timestamp 1624635492
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1624635492
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1624635492
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_192
timestamp 1624635492
transform 1 0 18768 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1624635492
transform 1 0 19044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1624635492
transform 1 0 18492 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_207
timestamp 1624635492
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_201
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_198
timestamp 1624635492
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1624635492
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20148 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1624635492
transform -1 0 20148 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 19964 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _72_
timestamp 1624635492
transform -1 0 21436 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20332 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1624635492
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1624635492
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1624635492
transform 1 0 21160 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1624635492
transform 1 0 21528 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624635492
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1624635492
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1624635492
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1624635492
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1624635492
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1624635492
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12604 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 12144 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1624635492
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1624635492
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1624635492
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14260 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1624635492
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1624635492
transform -1 0 16652 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1624635492
transform -1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1624635492
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1624635492
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17572 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17388 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1624635492
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1624635492
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1624635492
transform -1 0 19504 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19688 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1624635492
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1624635492
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_218
timestamp 1624635492
transform 1 0 21160 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_222
timestamp 1624635492
transform 1 0 21528 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1624635492
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624635492
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1624635492
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1624635492
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1624635492
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1624635492
transform 1 0 10212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1624635492
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_123
timestamp 1624635492
transform 1 0 12420 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14076 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_131
timestamp 1624635492
transform 1 0 13156 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1624635492
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1624635492
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14628 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1624635492
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1624635492
transform -1 0 18308 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1624635492
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1624635492
transform 1 0 17572 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1624635492
transform 1 0 17940 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1624635492
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19780 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18492 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1624635492
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1624635492
transform 1 0 20792 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1624635492
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1624635492
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1624635492
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform -1 0 1932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1624635492
transform -1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1624635492
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_13
timestamp 1624635492
transform 1 0 2300 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1624635492
transform 1 0 3404 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1624635492
transform 1 0 4508 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_49
timestamp 1624635492
transform 1 0 5612 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1624635492
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1624635492
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1624635492
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1624635492
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1624635492
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1624635492
transform 1 0 13892 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_143
timestamp 1624635492
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16652 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16192 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1624635492
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1624635492
transform 1 0 14536 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_153
timestamp 1624635492
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_164
timestamp 1624635492
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18492 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1624635492
transform -1 0 17480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1624635492
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_172
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_178
timestamp 1624635492
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 20424 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1624635492
transform 1 0 18492 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_193
timestamp 1624635492
transform 1 0 18860 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _70_
timestamp 1624635492
transform -1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1624635492
transform 1 0 20424 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1624635492
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1624635492
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624635492
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1624635492
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1624635492
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1624635492
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1624635492
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1624635492
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1624635492
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1624635492
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1624635492
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15640 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 15364 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1624635492
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_155
timestamp 1624635492
transform 1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1624635492
transform -1 0 17664 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17848 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_174
timestamp 1624635492
transform 1 0 17112 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1624635492
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20148 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1624635492
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_201
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_207
timestamp 1624635492
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1624635492
transform -1 0 21068 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _88_
timestamp 1624635492
transform -1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1624635492
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1624635492
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1624635492
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1624635492
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1624635492
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1624635492
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1624635492
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1624635492
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1624635492
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1624635492
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1624635492
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1624635492
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1624635492
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1624635492
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1624635492
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1624635492
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1624635492
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1624635492
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1624635492
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1624635492
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1624635492
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1624635492
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_156
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_151
timestamp 1624635492
transform 1 0 14996 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1624635492
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1624635492
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1624635492
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp 1624635492
transform 1 0 15548 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1624635492
transform -1 0 16652 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 17664 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17112 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1624635492
transform -1 0 18124 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1624635492
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1624635492
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1624635492
transform 1 0 18124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1624635492
transform 1 0 18492 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1624635492
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 18952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1624635492
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_194
timestamp 1624635492
transform 1 0 18952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1624635492
transform -1 0 19320 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624635492
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_198
timestamp 1624635492
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1624635492
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 19780 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19872 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_203
timestamp 1624635492
transform 1 0 19780 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_204
timestamp 1624635492
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20332 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1624635492
transform -1 0 20424 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1624635492
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_209
timestamp 1624635492
transform 1 0 20332 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1624635492
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1624635492
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1624635492
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_215
timestamp 1624635492
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform 1 0 21068 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 21068 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1624635492
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1624635492
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1624635492
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1624635492
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1624635492
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1624635492
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1624635492
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1624635492
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1624635492
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11408 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_106
timestamp 1624635492
transform 1 0 10856 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1624635492
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1624635492
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1624635492
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1624635492
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1624635492
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 17664 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 18308 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_172
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1624635492
transform 1 0 17664 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1624635492
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_187
timestamp 1624635492
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21252 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1624635492
transform -1 0 19964 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1624635492
transform -1 0 19504 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_mem_bottom_track_1.prog_clk_A
timestamp 1624635492
transform -1 0 18676 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1624635492
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_195
timestamp 1624635492
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1624635492
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_205
timestamp 1624635492
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1624635492
transform 1 0 21252 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1624635492
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1624635492
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1624635492
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1624635492
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9752 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_92
timestamp 1624635492
transform 1 0 9568 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1624635492
transform 1 0 10028 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1624635492
transform 1 0 11132 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1624635492
transform 1 0 12236 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_133
timestamp 1624635492
transform 1 0 13340 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1624635492
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1624635492
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1624635492
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1624635492
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1624635492
transform -1 0 20424 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 19964 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1624635492
transform 1 0 18768 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1624635492
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_201
timestamp 1624635492
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_205
timestamp 1624635492
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1624635492
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform 1 0 21068 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1624635492
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1624635492
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1624635492
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1624635492
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1624635492
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1624635492
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1624635492
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1624635492
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1624635492
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1624635492
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12144 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1624635492
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_120
timestamp 1624635492
transform 1 0 12144 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_132
timestamp 1624635492
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_144
timestamp 1624635492
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_156
timestamp 1624635492
transform 1 0 15456 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_168
timestamp 1624635492
transform 1 0 16560 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1624635492
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1624635492
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1624635492
transform 1 0 20240 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1624635492
transform 1 0 20608 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform 1 0 21068 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_215
timestamp 1624635492
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1624635492
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1624635492
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1624635492
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1624635492
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1624635492
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1624635492
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1624635492
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1624635492
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1624635492
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1624635492
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1624635492
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_149
timestamp 1624635492
transform 1 0 14812 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_161
timestamp 1624635492
transform 1 0 15916 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_173
timestamp 1624635492
transform 1 0 17020 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_185
timestamp 1624635492
transform 1 0 18124 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1624635492
transform -1 0 20332 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1624635492
transform 1 0 19228 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1624635492
transform 1 0 19596 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_205
timestamp 1624635492
transform 1 0 19964 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform 1 0 21068 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform 1 0 20516 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1624635492
transform 1 0 20332 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1624635492
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1624635492
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1624635492
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1624635492
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1624635492
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1624635492
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1624635492
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1624635492
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1624635492
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1624635492
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1624635492
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1624635492
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1624635492
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1624635492
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1624635492
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20148 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1624635492
transform 1 0 19136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1624635492
transform 1 0 20148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1624635492
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform 1 0 21068 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1624635492
transform 1 0 20516 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1624635492
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1624635492
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1624635492
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1624635492
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1624635492
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1624635492
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1624635492
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1624635492
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1624635492
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1624635492
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1624635492
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1624635492
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1624635492
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1624635492
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1624635492
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1624635492
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12144 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1624635492
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1624635492
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1624635492
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_120
timestamp 1624635492
transform 1 0 12144 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1624635492
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_132
timestamp 1624635492
transform 1 0 13248 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_144
timestamp 1624635492
transform 1 0 14352 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1624635492
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1624635492
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18124 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1624635492
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_180
timestamp 1624635492
transform 1 0 17664 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_185
timestamp 1624635492
transform 1 0 18124 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_168
timestamp 1624635492
transform 1 0 16560 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1624635492
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1624635492
transform -1 0 20424 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1624635492
transform -1 0 20332 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19872 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1624635492
transform 1 0 19228 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_201
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1624635492
transform 1 0 19136 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_200
timestamp 1624635492
transform 1 0 19504 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1624635492
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1624635492
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1624635492
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1624635492
transform 1 0 20608 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1624635492
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1624635492
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform 1 0 21068 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform 1 0 21068 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1624635492
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1624635492
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1624635492
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1624635492
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1624635492
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1624635492
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 8096 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_66
timestamp 1624635492
transform 1 0 7176 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1624635492
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_79
timestamp 1624635492
transform 1 0 8372 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1624635492
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1624635492
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1624635492
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1624635492
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1624635492
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1624635492
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1624635492
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1624635492
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1624635492
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1624635492
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform 1 0 21068 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 1624635492
transform 1 0 20332 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1624635492
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1624635492
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1624635492
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1624635492
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1624635492
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1624635492
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_51
timestamp 1624635492
transform 1 0 5796 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1624635492
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_82
timestamp 1624635492
transform 1 0 8648 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9384 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1624635492
transform 1 0 9660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _62_
timestamp 1624635492
transform 1 0 12144 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_105
timestamp 1624635492
transform 1 0 10764 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1624635492
transform 1 0 11500 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1624635492
transform 1 0 12052 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1624635492
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1624635492
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1624635492
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1624635492
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1624635492
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20148 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_196
timestamp 1624635492
transform 1 0 19136 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_207
timestamp 1624635492
transform 1 0 20148 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1624635492
transform 1 0 21068 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1624635492
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1624635492
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1624635492
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1624635492
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1624635492
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_54
timestamp 1624635492
transform 1 0 6072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1624635492
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1624635492
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1624635492
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1624635492
transform 1 0 11316 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1624635492
transform 1 0 11684 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_119
timestamp 1624635492
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_131
timestamp 1624635492
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1624635492
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1624635492
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_180
timestamp 1624635492
transform 1 0 17664 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20148 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18768 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_188
timestamp 1624635492
transform 1 0 18400 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_192
timestamp 1624635492
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_201
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1624635492
transform 1 0 20148 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1624635492
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1624635492
transform 1 0 21068 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_211
timestamp 1624635492
transform 1 0 20516 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1624635492
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1624635492
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1624635492
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1624635492
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1624635492
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1624635492
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _48_
timestamp 1624635492
transform 1 0 6624 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1624635492
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_64
timestamp 1624635492
transform 1 0 6992 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_76
timestamp 1624635492
transform 1 0 8096 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_88
timestamp 1624635492
transform 1 0 9200 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_100
timestamp 1624635492
transform 1 0 10304 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _65_
timestamp 1624635492
transform 1 0 12604 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_112
timestamp 1624635492
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_115
timestamp 1624635492
transform 1 0 11684 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1624635492
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_128
timestamp 1624635492
transform 1 0 12880 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_140
timestamp 1624635492
transform 1 0 13984 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_152
timestamp 1624635492
transform 1 0 15088 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_164
timestamp 1624635492
transform 1 0 16192 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_170
timestamp 1624635492
transform 1 0 16744 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1624635492
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1624635492
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1624635492
transform 1 0 20148 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1624635492
transform 1 0 19688 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_196
timestamp 1624635492
transform 1 0 19136 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_205
timestamp 1624635492
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1624635492
transform 1 0 20608 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform 1 0 21068 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1624635492
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1624635492
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1624635492
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1624635492
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1624635492
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1624635492
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1624635492
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1624635492
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1624635492
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1624635492
transform 1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1624635492
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1624635492
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1624635492
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1624635492
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1624635492
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1624635492
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1624635492
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1624635492
transform -1 0 17664 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform 1 0 18124 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1624635492
transform 1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 1624635492
transform 1 0 16928 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_175
timestamp 1624635492
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1624635492
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_184
timestamp 1624635492
transform 1 0 18032 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform 1 0 20056 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_189
timestamp 1624635492
transform 1 0 18492 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1624635492
transform 1 0 19228 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_205
timestamp 1624635492
transform 1 0 19964 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform 1 0 21068 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1624635492
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1624635492
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1624635492
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1624635492
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_27
timestamp 1624635492
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_30
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform -1 0 5980 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 6716 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_42
timestamp 1624635492
transform 1 0 4968 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_53
timestamp 1624635492
transform 1 0 5980 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1624635492
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_61
timestamp 1624635492
transform 1 0 6716 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_73
timestamp 1624635492
transform 1 0 7820 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1624635492
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_88
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_100
timestamp 1624635492
transform 1 0 10304 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_112
timestamp 1624635492
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_117
timestamp 1624635492
transform 1 0 11868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_129
timestamp 1624635492
transform 1 0 12972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1624635492
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_146
timestamp 1624635492
transform 1 0 14536 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_158
timestamp 1624635492
transform 1 0 15640 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 18124 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_170
timestamp 1624635492
transform 1 0 16744 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1624635492
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_185
timestamp 1624635492
transform 1 0 18124 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_195
timestamp 1624635492
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1624635492
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_204
timestamp 1624635492
transform 1 0 19872 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1624635492
transform -1 0 21436 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform 1 0 20516 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1624635492
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1624635492
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1624635492
transform 1 0 21436 0 1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 5722 22200 5778 23000 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_1_
port 2 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 ccff_tail
port 4 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 5 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[10]
port 6 nsew signal input
rlabel metal3 s 22200 8848 23000 8968 6 chanx_right_in[11]
port 7 nsew signal input
rlabel metal3 s 22200 9256 23000 9376 6 chanx_right_in[12]
port 8 nsew signal input
rlabel metal3 s 22200 9664 23000 9784 6 chanx_right_in[13]
port 9 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[14]
port 10 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[15]
port 11 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[16]
port 12 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[17]
port 13 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[18]
port 14 nsew signal input
rlabel metal3 s 22200 12520 23000 12640 6 chanx_right_in[19]
port 15 nsew signal input
rlabel metal3 s 22200 4224 23000 4344 6 chanx_right_in[1]
port 16 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[2]
port 17 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 18 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[4]
port 19 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[5]
port 20 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[6]
port 21 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[7]
port 22 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[8]
port 23 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[9]
port 24 nsew signal input
rlabel metal3 s 22200 12928 23000 13048 6 chanx_right_out[0]
port 25 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[10]
port 26 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[11]
port 27 nsew signal tristate
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[12]
port 28 nsew signal tristate
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[13]
port 29 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[14]
port 30 nsew signal tristate
rlabel metal3 s 22200 19864 23000 19984 6 chanx_right_out[15]
port 31 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[16]
port 32 nsew signal tristate
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[17]
port 33 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[18]
port 34 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[19]
port 35 nsew signal tristate
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[1]
port 36 nsew signal tristate
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[2]
port 37 nsew signal tristate
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[3]
port 38 nsew signal tristate
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[4]
port 39 nsew signal tristate
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[5]
port 40 nsew signal tristate
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[6]
port 41 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[7]
port 42 nsew signal tristate
rlabel metal3 s 22200 16600 23000 16720 6 chanx_right_out[8]
port 43 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[9]
port 44 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 chany_bottom_in[0]
port 45 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_in[10]
port 46 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_in[11]
port 47 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[12]
port 48 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[13]
port 49 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 chany_bottom_in[14]
port 50 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[15]
port 51 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[16]
port 52 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[17]
port 53 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[18]
port 54 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 chany_bottom_in[19]
port 55 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 chany_bottom_in[1]
port 56 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_in[2]
port 57 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_in[3]
port 58 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 chany_bottom_in[4]
port 59 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_in[5]
port 60 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_in[6]
port 61 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_in[7]
port 62 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[8]
port 63 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_in[9]
port 64 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_out[0]
port 65 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 chany_bottom_out[10]
port 66 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[11]
port 67 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[12]
port 68 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[13]
port 69 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[14]
port 70 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[15]
port 71 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[16]
port 72 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[17]
port 73 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[18]
port 74 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[19]
port 75 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_out[1]
port 76 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[2]
port 77 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[3]
port 78 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_out[4]
port 79 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[5]
port 80 nsew signal tristate
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_out[6]
port 81 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[7]
port 82 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[8]
port 83 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[9]
port 84 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 prog_clk_0_E_in
port 85 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 86 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 87 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 88 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 89 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 90 nsew signal input
rlabel metal3 s 22200 2320 23000 2440 6 right_bottom_grid_pin_39_
port 91 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 92 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_41_
port 93 nsew signal input
rlabel metal3 s 22200 22584 23000 22704 6 right_top_grid_pin_1_
port 94 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 95 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 96 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 97 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 98 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 99 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
