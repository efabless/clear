magic
tech sky130A
magscale 1 2
timestamp 1625831969
<< obsli1 >>
rect 15690 6671 492482 573567
<< obsm1 >>
rect 5704 6390 502384 573598
<< metal2 >>
rect 13804 575726 13860 576526
rect 32204 575726 32260 576526
rect 50696 575726 50752 576526
rect 69188 575726 69244 576526
rect 87680 575726 87736 576526
rect 106172 575726 106228 576526
rect 124664 575726 124720 576526
rect 143156 575726 143212 576526
rect 161648 575726 161704 576526
rect 180140 575726 180196 576526
rect 198540 575726 198596 576526
rect 217032 575726 217088 576526
rect 235524 575726 235580 576526
rect 254016 575726 254072 576526
rect 272508 575726 272564 576526
rect 291000 575726 291056 576526
rect 309492 575726 309548 576526
rect 327984 575726 328040 576526
rect 346476 575726 346532 576526
rect 364876 575726 364932 576526
rect 383368 575726 383424 576526
rect 401860 575726 401916 576526
rect 420352 575726 420408 576526
rect 438844 575726 438900 576526
rect 457336 575726 457392 576526
rect 475828 575726 475884 576526
rect 494320 575726 494376 576526
rect 5708 3526 5764 4326
rect 8008 3526 8064 4326
rect 10308 3526 10364 4326
rect 12608 3526 12664 4326
rect 14908 3526 14964 4326
rect 17208 3526 17264 4326
rect 19508 3526 19564 4326
rect 21808 3526 21864 4326
rect 24108 3526 24164 4326
rect 26500 3526 26556 4326
rect 28800 3526 28856 4326
rect 31100 3526 31156 4326
rect 33400 3526 33456 4326
rect 35700 3526 35756 4326
rect 38000 3526 38056 4326
rect 40300 3526 40356 4326
rect 42600 3526 42656 4326
rect 44900 3526 44956 4326
rect 47292 3526 47348 4326
rect 49592 3526 49648 4326
rect 51892 3526 51948 4326
rect 54192 3526 54248 4326
rect 56492 3526 56548 4326
rect 58792 3526 58848 4326
rect 61092 3526 61148 4326
rect 63392 3526 63448 4326
rect 65692 3526 65748 4326
rect 68084 3526 68140 4326
rect 70384 3526 70440 4326
rect 72684 3526 72740 4326
rect 74984 3526 75040 4326
rect 77284 3526 77340 4326
rect 79584 3526 79640 4326
rect 81884 3526 81940 4326
rect 84184 3526 84240 4326
rect 86484 3526 86540 4326
rect 88876 3526 88932 4326
rect 91176 3526 91232 4326
rect 93476 3526 93532 4326
rect 95776 3526 95832 4326
rect 98076 3526 98132 4326
rect 100376 3526 100432 4326
rect 102676 3526 102732 4326
rect 104976 3526 105032 4326
rect 107276 3526 107332 4326
rect 109668 3526 109724 4326
rect 111968 3526 112024 4326
rect 114268 3526 114324 4326
rect 116568 3526 116624 4326
rect 118868 3526 118924 4326
rect 121168 3526 121224 4326
rect 123468 3526 123524 4326
rect 125768 3526 125824 4326
rect 128068 3526 128124 4326
rect 130460 3526 130516 4326
rect 132760 3526 132816 4326
rect 135060 3526 135116 4326
rect 137360 3526 137416 4326
rect 139660 3526 139716 4326
rect 141960 3526 142016 4326
rect 144260 3526 144316 4326
rect 146560 3526 146616 4326
rect 148860 3526 148916 4326
rect 151252 3526 151308 4326
rect 153552 3526 153608 4326
rect 155852 3526 155908 4326
rect 158152 3526 158208 4326
rect 160452 3526 160508 4326
rect 162752 3526 162808 4326
rect 165052 3526 165108 4326
rect 167352 3526 167408 4326
rect 169652 3526 169708 4326
rect 172044 3526 172100 4326
rect 174344 3526 174400 4326
rect 176644 3526 176700 4326
rect 178944 3526 179000 4326
rect 181244 3526 181300 4326
rect 183544 3526 183600 4326
rect 185844 3526 185900 4326
rect 188144 3526 188200 4326
rect 190444 3526 190500 4326
rect 192836 3526 192892 4326
rect 195136 3526 195192 4326
rect 197436 3526 197492 4326
rect 199736 3526 199792 4326
rect 202036 3526 202092 4326
rect 204336 3526 204392 4326
rect 206636 3526 206692 4326
rect 208936 3526 208992 4326
rect 211236 3526 211292 4326
rect 213628 3526 213684 4326
rect 215928 3526 215984 4326
rect 218228 3526 218284 4326
rect 220528 3526 220584 4326
rect 222828 3526 222884 4326
rect 225128 3526 225184 4326
rect 227428 3526 227484 4326
rect 229728 3526 229784 4326
rect 232028 3526 232084 4326
rect 234420 3526 234476 4326
rect 236720 3526 236776 4326
rect 239020 3526 239076 4326
rect 241320 3526 241376 4326
rect 243620 3526 243676 4326
rect 245920 3526 245976 4326
rect 248220 3526 248276 4326
rect 250520 3526 250576 4326
rect 252820 3526 252876 4326
rect 255212 3526 255268 4326
rect 257512 3526 257568 4326
rect 259812 3526 259868 4326
rect 262112 3526 262168 4326
rect 264412 3526 264468 4326
rect 266712 3526 266768 4326
rect 269012 3526 269068 4326
rect 271312 3526 271368 4326
rect 273612 3526 273668 4326
rect 276004 3526 276060 4326
rect 278304 3526 278360 4326
rect 280604 3526 280660 4326
rect 282904 3526 282960 4326
rect 285204 3526 285260 4326
rect 287504 3526 287560 4326
rect 289804 3526 289860 4326
rect 292104 3526 292160 4326
rect 294404 3526 294460 4326
rect 296796 3526 296852 4326
rect 299096 3526 299152 4326
rect 301396 3526 301452 4326
rect 303696 3526 303752 4326
rect 305996 3526 306052 4326
rect 308296 3526 308352 4326
rect 310596 3526 310652 4326
rect 312896 3526 312952 4326
rect 315196 3526 315252 4326
rect 317588 3526 317644 4326
rect 319888 3526 319944 4326
rect 322188 3526 322244 4326
rect 324488 3526 324544 4326
rect 326788 3526 326844 4326
rect 329088 3526 329144 4326
rect 331388 3526 331444 4326
rect 333688 3526 333744 4326
rect 335988 3526 336044 4326
rect 338380 3526 338436 4326
rect 340680 3526 340736 4326
rect 342980 3526 343036 4326
rect 345280 3526 345336 4326
rect 347580 3526 347636 4326
rect 349880 3526 349936 4326
rect 352180 3526 352236 4326
rect 354480 3526 354536 4326
rect 356780 3526 356836 4326
rect 359172 3526 359228 4326
rect 361472 3526 361528 4326
rect 363772 3526 363828 4326
rect 366072 3526 366128 4326
rect 368372 3526 368428 4326
rect 370672 3526 370728 4326
rect 372972 3526 373028 4326
rect 375272 3526 375328 4326
rect 377572 3526 377628 4326
rect 379964 3526 380020 4326
rect 382264 3526 382320 4326
rect 384564 3526 384620 4326
rect 386864 3526 386920 4326
rect 389164 3526 389220 4326
rect 391464 3526 391520 4326
rect 393764 3526 393820 4326
rect 396064 3526 396120 4326
rect 398364 3526 398420 4326
rect 400756 3526 400812 4326
rect 403056 3526 403112 4326
rect 405356 3526 405412 4326
rect 407656 3526 407712 4326
rect 409956 3526 410012 4326
rect 412256 3526 412312 4326
rect 414556 3526 414612 4326
rect 416856 3526 416912 4326
rect 419156 3526 419212 4326
rect 421548 3526 421604 4326
rect 423848 3526 423904 4326
rect 426148 3526 426204 4326
rect 428448 3526 428504 4326
rect 430748 3526 430804 4326
rect 433048 3526 433104 4326
rect 435348 3526 435404 4326
rect 437648 3526 437704 4326
rect 439948 3526 440004 4326
rect 442340 3526 442396 4326
rect 444640 3526 444696 4326
rect 446940 3526 446996 4326
rect 449240 3526 449296 4326
rect 451540 3526 451596 4326
rect 453840 3526 453896 4326
rect 456140 3526 456196 4326
rect 458440 3526 458496 4326
rect 460740 3526 460796 4326
rect 463132 3526 463188 4326
rect 465432 3526 465488 4326
rect 467732 3526 467788 4326
rect 470032 3526 470088 4326
rect 472332 3526 472388 4326
rect 474632 3526 474688 4326
rect 476932 3526 476988 4326
rect 479232 3526 479288 4326
rect 481532 3526 481588 4326
rect 483924 3526 483980 4326
rect 486224 3526 486280 4326
rect 488524 3526 488580 4326
rect 490824 3526 490880 4326
rect 493124 3526 493180 4326
rect 495424 3526 495480 4326
rect 497724 3526 497780 4326
rect 500024 3526 500080 4326
rect 502324 3526 502380 4326
<< obsm2 >>
rect 5710 575670 13748 575726
rect 13916 575670 32148 575726
rect 32316 575670 50640 575726
rect 50808 575670 69132 575726
rect 69300 575670 87624 575726
rect 87792 575670 106116 575726
rect 106284 575670 124608 575726
rect 124776 575670 143100 575726
rect 143268 575670 161592 575726
rect 161760 575670 180084 575726
rect 180252 575670 198484 575726
rect 198652 575670 216976 575726
rect 217144 575670 235468 575726
rect 235636 575670 253960 575726
rect 254128 575670 272452 575726
rect 272620 575670 290944 575726
rect 291112 575670 309436 575726
rect 309604 575670 327928 575726
rect 328096 575670 346420 575726
rect 346588 575670 364820 575726
rect 364988 575670 383312 575726
rect 383480 575670 401804 575726
rect 401972 575670 420296 575726
rect 420464 575670 438788 575726
rect 438956 575670 457280 575726
rect 457448 575670 475772 575726
rect 475940 575670 494264 575726
rect 494432 575670 502378 575726
rect 5710 4382 502378 575670
rect 5820 4326 7952 4382
rect 8120 4326 10252 4382
rect 10420 4326 12552 4382
rect 12720 4326 14852 4382
rect 15020 4326 17152 4382
rect 17320 4326 19452 4382
rect 19620 4326 21752 4382
rect 21920 4326 24052 4382
rect 24220 4326 26444 4382
rect 26612 4326 28744 4382
rect 28912 4326 31044 4382
rect 31212 4326 33344 4382
rect 33512 4326 35644 4382
rect 35812 4326 37944 4382
rect 38112 4326 40244 4382
rect 40412 4326 42544 4382
rect 42712 4326 44844 4382
rect 45012 4326 47236 4382
rect 47404 4326 49536 4382
rect 49704 4326 51836 4382
rect 52004 4326 54136 4382
rect 54304 4326 56436 4382
rect 56604 4326 58736 4382
rect 58904 4326 61036 4382
rect 61204 4326 63336 4382
rect 63504 4326 65636 4382
rect 65804 4326 68028 4382
rect 68196 4326 70328 4382
rect 70496 4326 72628 4382
rect 72796 4326 74928 4382
rect 75096 4326 77228 4382
rect 77396 4326 79528 4382
rect 79696 4326 81828 4382
rect 81996 4326 84128 4382
rect 84296 4326 86428 4382
rect 86596 4326 88820 4382
rect 88988 4326 91120 4382
rect 91288 4326 93420 4382
rect 93588 4326 95720 4382
rect 95888 4326 98020 4382
rect 98188 4326 100320 4382
rect 100488 4326 102620 4382
rect 102788 4326 104920 4382
rect 105088 4326 107220 4382
rect 107388 4326 109612 4382
rect 109780 4326 111912 4382
rect 112080 4326 114212 4382
rect 114380 4326 116512 4382
rect 116680 4326 118812 4382
rect 118980 4326 121112 4382
rect 121280 4326 123412 4382
rect 123580 4326 125712 4382
rect 125880 4326 128012 4382
rect 128180 4326 130404 4382
rect 130572 4326 132704 4382
rect 132872 4326 135004 4382
rect 135172 4326 137304 4382
rect 137472 4326 139604 4382
rect 139772 4326 141904 4382
rect 142072 4326 144204 4382
rect 144372 4326 146504 4382
rect 146672 4326 148804 4382
rect 148972 4326 151196 4382
rect 151364 4326 153496 4382
rect 153664 4326 155796 4382
rect 155964 4326 158096 4382
rect 158264 4326 160396 4382
rect 160564 4326 162696 4382
rect 162864 4326 164996 4382
rect 165164 4326 167296 4382
rect 167464 4326 169596 4382
rect 169764 4326 171988 4382
rect 172156 4326 174288 4382
rect 174456 4326 176588 4382
rect 176756 4326 178888 4382
rect 179056 4326 181188 4382
rect 181356 4326 183488 4382
rect 183656 4326 185788 4382
rect 185956 4326 188088 4382
rect 188256 4326 190388 4382
rect 190556 4326 192780 4382
rect 192948 4326 195080 4382
rect 195248 4326 197380 4382
rect 197548 4326 199680 4382
rect 199848 4326 201980 4382
rect 202148 4326 204280 4382
rect 204448 4326 206580 4382
rect 206748 4326 208880 4382
rect 209048 4326 211180 4382
rect 211348 4326 213572 4382
rect 213740 4326 215872 4382
rect 216040 4326 218172 4382
rect 218340 4326 220472 4382
rect 220640 4326 222772 4382
rect 222940 4326 225072 4382
rect 225240 4326 227372 4382
rect 227540 4326 229672 4382
rect 229840 4326 231972 4382
rect 232140 4326 234364 4382
rect 234532 4326 236664 4382
rect 236832 4326 238964 4382
rect 239132 4326 241264 4382
rect 241432 4326 243564 4382
rect 243732 4326 245864 4382
rect 246032 4326 248164 4382
rect 248332 4326 250464 4382
rect 250632 4326 252764 4382
rect 252932 4326 255156 4382
rect 255324 4326 257456 4382
rect 257624 4326 259756 4382
rect 259924 4326 262056 4382
rect 262224 4326 264356 4382
rect 264524 4326 266656 4382
rect 266824 4326 268956 4382
rect 269124 4326 271256 4382
rect 271424 4326 273556 4382
rect 273724 4326 275948 4382
rect 276116 4326 278248 4382
rect 278416 4326 280548 4382
rect 280716 4326 282848 4382
rect 283016 4326 285148 4382
rect 285316 4326 287448 4382
rect 287616 4326 289748 4382
rect 289916 4326 292048 4382
rect 292216 4326 294348 4382
rect 294516 4326 296740 4382
rect 296908 4326 299040 4382
rect 299208 4326 301340 4382
rect 301508 4326 303640 4382
rect 303808 4326 305940 4382
rect 306108 4326 308240 4382
rect 308408 4326 310540 4382
rect 310708 4326 312840 4382
rect 313008 4326 315140 4382
rect 315308 4326 317532 4382
rect 317700 4326 319832 4382
rect 320000 4326 322132 4382
rect 322300 4326 324432 4382
rect 324600 4326 326732 4382
rect 326900 4326 329032 4382
rect 329200 4326 331332 4382
rect 331500 4326 333632 4382
rect 333800 4326 335932 4382
rect 336100 4326 338324 4382
rect 338492 4326 340624 4382
rect 340792 4326 342924 4382
rect 343092 4326 345224 4382
rect 345392 4326 347524 4382
rect 347692 4326 349824 4382
rect 349992 4326 352124 4382
rect 352292 4326 354424 4382
rect 354592 4326 356724 4382
rect 356892 4326 359116 4382
rect 359284 4326 361416 4382
rect 361584 4326 363716 4382
rect 363884 4326 366016 4382
rect 366184 4326 368316 4382
rect 368484 4326 370616 4382
rect 370784 4326 372916 4382
rect 373084 4326 375216 4382
rect 375384 4326 377516 4382
rect 377684 4326 379908 4382
rect 380076 4326 382208 4382
rect 382376 4326 384508 4382
rect 384676 4326 386808 4382
rect 386976 4326 389108 4382
rect 389276 4326 391408 4382
rect 391576 4326 393708 4382
rect 393876 4326 396008 4382
rect 396176 4326 398308 4382
rect 398476 4326 400700 4382
rect 400868 4326 403000 4382
rect 403168 4326 405300 4382
rect 405468 4326 407600 4382
rect 407768 4326 409900 4382
rect 410068 4326 412200 4382
rect 412368 4326 414500 4382
rect 414668 4326 416800 4382
rect 416968 4326 419100 4382
rect 419268 4326 421492 4382
rect 421660 4326 423792 4382
rect 423960 4326 426092 4382
rect 426260 4326 428392 4382
rect 428560 4326 430692 4382
rect 430860 4326 432992 4382
rect 433160 4326 435292 4382
rect 435460 4326 437592 4382
rect 437760 4326 439892 4382
rect 440060 4326 442284 4382
rect 442452 4326 444584 4382
rect 444752 4326 446884 4382
rect 447052 4326 449184 4382
rect 449352 4326 451484 4382
rect 451652 4326 453784 4382
rect 453952 4326 456084 4382
rect 456252 4326 458384 4382
rect 458552 4326 460684 4382
rect 460852 4326 463076 4382
rect 463244 4326 465376 4382
rect 465544 4326 467676 4382
rect 467844 4326 469976 4382
rect 470144 4326 472276 4382
rect 472444 4326 474576 4382
rect 474744 4326 476876 4382
rect 477044 4326 479176 4382
rect 479344 4326 481476 4382
rect 481644 4326 483868 4382
rect 484036 4326 486168 4382
rect 486336 4326 488468 4382
rect 488636 4326 490768 4382
rect 490936 4326 493068 4382
rect 493236 4326 495368 4382
rect 495536 4326 497668 4382
rect 497836 4326 499968 4382
rect 500136 4326 502268 4382
<< metal3 >>
rect 4586 566438 5386 566558
rect 502786 564398 503586 564518
rect 4586 546718 5386 546838
rect 502786 540462 503586 540582
rect 4586 526998 5386 527118
rect 502786 516662 503586 516782
rect 4586 507142 5386 507262
rect 502786 492726 503586 492846
rect 4586 487422 5386 487542
rect 502786 468926 503586 469046
rect 4586 467702 5386 467822
rect 4586 447982 5386 448102
rect 502786 444990 503586 445110
rect 4586 428126 5386 428246
rect 502786 421190 503586 421310
rect 4586 408406 5386 408526
rect 502786 397254 503586 397374
rect 4586 388686 5386 388806
rect 502786 373454 503586 373574
rect 4586 368830 5386 368950
rect 502786 349518 503586 349638
rect 4586 349110 5386 349230
rect 4586 329390 5386 329510
rect 502786 325718 503586 325838
rect 4586 309670 5386 309790
rect 502786 301782 503586 301902
rect 4586 289814 5386 289934
rect 502786 277846 503586 277966
rect 4586 270094 5386 270214
rect 502786 254046 503586 254166
rect 4586 250374 5386 250494
rect 4586 230654 5386 230774
rect 502786 230110 503586 230230
rect 4586 210798 5386 210918
rect 502786 206310 503586 206430
rect 4586 191078 5386 191198
rect 502786 182374 503586 182494
rect 4586 171358 5386 171478
rect 502786 158574 503586 158694
rect 4586 151502 5386 151622
rect 502786 134638 503586 134758
rect 4586 131782 5386 131902
rect 4586 112062 5386 112182
rect 502786 110838 503586 110958
rect 4586 92342 5386 92462
rect 502786 86902 503586 87022
rect 4586 72486 5386 72606
rect 502786 63102 503586 63222
rect 4586 52766 5386 52886
rect 502786 39166 503586 39286
rect 4586 33046 5386 33166
rect 502786 15366 503586 15486
rect 4586 13326 5386 13446
<< obsm3 >>
rect 5386 566638 502786 573583
rect 5466 566358 502786 566638
rect 5386 564598 502786 566358
rect 5386 564318 502706 564598
rect 5386 546918 502786 564318
rect 5466 546638 502786 546918
rect 5386 540662 502786 546638
rect 5386 540382 502706 540662
rect 5386 527198 502786 540382
rect 5466 526918 502786 527198
rect 5386 516862 502786 526918
rect 5386 516582 502706 516862
rect 5386 507342 502786 516582
rect 5466 507062 502786 507342
rect 5386 492926 502786 507062
rect 5386 492646 502706 492926
rect 5386 487622 502786 492646
rect 5466 487342 502786 487622
rect 5386 469126 502786 487342
rect 5386 468846 502706 469126
rect 5386 467902 502786 468846
rect 5466 467622 502786 467902
rect 5386 448182 502786 467622
rect 5466 447902 502786 448182
rect 5386 445190 502786 447902
rect 5386 444910 502706 445190
rect 5386 428326 502786 444910
rect 5466 428046 502786 428326
rect 5386 421390 502786 428046
rect 5386 421110 502706 421390
rect 5386 408606 502786 421110
rect 5466 408326 502786 408606
rect 5386 397454 502786 408326
rect 5386 397174 502706 397454
rect 5386 388886 502786 397174
rect 5466 388606 502786 388886
rect 5386 373654 502786 388606
rect 5386 373374 502706 373654
rect 5386 369030 502786 373374
rect 5466 368750 502786 369030
rect 5386 349718 502786 368750
rect 5386 349438 502706 349718
rect 5386 349310 502786 349438
rect 5466 349030 502786 349310
rect 5386 329590 502786 349030
rect 5466 329310 502786 329590
rect 5386 325918 502786 329310
rect 5386 325638 502706 325918
rect 5386 309870 502786 325638
rect 5466 309590 502786 309870
rect 5386 301982 502786 309590
rect 5386 301702 502706 301982
rect 5386 290014 502786 301702
rect 5466 289734 502786 290014
rect 5386 278046 502786 289734
rect 5386 277766 502706 278046
rect 5386 270294 502786 277766
rect 5466 270014 502786 270294
rect 5386 254246 502786 270014
rect 5386 253966 502706 254246
rect 5386 250574 502786 253966
rect 5466 250294 502786 250574
rect 5386 230854 502786 250294
rect 5466 230574 502786 230854
rect 5386 230310 502786 230574
rect 5386 230030 502706 230310
rect 5386 210998 502786 230030
rect 5466 210718 502786 210998
rect 5386 206510 502786 210718
rect 5386 206230 502706 206510
rect 5386 191278 502786 206230
rect 5466 190998 502786 191278
rect 5386 182574 502786 190998
rect 5386 182294 502706 182574
rect 5386 171558 502786 182294
rect 5466 171278 502786 171558
rect 5386 158774 502786 171278
rect 5386 158494 502706 158774
rect 5386 151702 502786 158494
rect 5466 151422 502786 151702
rect 5386 134838 502786 151422
rect 5386 134558 502706 134838
rect 5386 131982 502786 134558
rect 5466 131702 502786 131982
rect 5386 112262 502786 131702
rect 5466 111982 502786 112262
rect 5386 111038 502786 111982
rect 5386 110758 502706 111038
rect 5386 92542 502786 110758
rect 5466 92262 502786 92542
rect 5386 87102 502786 92262
rect 5386 86822 502706 87102
rect 5386 72686 502786 86822
rect 5466 72406 502786 72686
rect 5386 63302 502786 72406
rect 5386 63022 502706 63302
rect 5386 52966 502786 63022
rect 5466 52686 502786 52966
rect 5386 39366 502786 52686
rect 5386 39086 502706 39366
rect 5386 33246 502786 39086
rect 5466 32966 502786 33246
rect 5386 15566 502786 32966
rect 5386 15286 502706 15566
rect 5386 13526 502786 15286
rect 5466 13353 502786 13526
<< metal4 >>
rect 0 12 900 579872
rect 1240 1252 2140 578632
rect 505948 1252 506848 578632
rect 507188 12 508088 579872
<< obsm4 >>
rect 16973 19745 493047 573598
<< metal5 >>
rect 0 578972 508088 579872
rect 1240 577732 506848 578632
rect 0 572252 508088 573152
rect 0 567752 508088 568652
rect 0 563252 508088 564152
rect 0 558752 508088 559652
rect 0 554252 508088 555152
rect 0 549752 508088 550652
rect 0 545252 508088 546152
rect 0 540752 508088 541652
rect 0 536252 508088 537152
rect 0 531752 508088 532652
rect 0 527252 508088 528152
rect 0 522752 508088 523652
rect 0 518252 508088 519152
rect 0 513752 508088 514652
rect 0 509252 508088 510152
rect 0 504752 508088 505652
rect 0 500252 508088 501152
rect 0 495752 508088 496652
rect 0 491252 508088 492152
rect 0 486752 508088 487652
rect 0 482252 508088 483152
rect 0 477752 508088 478652
rect 0 473252 508088 474152
rect 0 468752 508088 469652
rect 0 464252 508088 465152
rect 0 459752 508088 460652
rect 0 455252 508088 456152
rect 0 450752 508088 451652
rect 0 446252 508088 447152
rect 0 441752 508088 442652
rect 0 437252 508088 438152
rect 0 432752 508088 433652
rect 0 428252 508088 429152
rect 0 423752 508088 424652
rect 0 419252 508088 420152
rect 0 414752 508088 415652
rect 0 410252 508088 411152
rect 0 405752 508088 406652
rect 0 401252 508088 402152
rect 0 396752 508088 397652
rect 0 392252 508088 393152
rect 0 387752 508088 388652
rect 0 383252 508088 384152
rect 0 378752 508088 379652
rect 0 374252 508088 375152
rect 0 369752 508088 370652
rect 0 365252 508088 366152
rect 0 360752 508088 361652
rect 0 356252 508088 357152
rect 0 351752 508088 352652
rect 0 347252 508088 348152
rect 0 342752 508088 343652
rect 0 338252 508088 339152
rect 0 333752 508088 334652
rect 0 329252 508088 330152
rect 0 324752 508088 325652
rect 0 320252 508088 321152
rect 0 315752 508088 316652
rect 0 311252 508088 312152
rect 0 306752 508088 307652
rect 0 302252 508088 303152
rect 0 297752 508088 298652
rect 0 293252 508088 294152
rect 0 288752 508088 289652
rect 0 284252 508088 285152
rect 0 279752 508088 280652
rect 0 275252 508088 276152
rect 0 270752 508088 271652
rect 0 266252 508088 267152
rect 0 261752 508088 262652
rect 0 257252 508088 258152
rect 0 252752 508088 253652
rect 0 248252 508088 249152
rect 0 243752 508088 244652
rect 0 239252 508088 240152
rect 0 234752 508088 235652
rect 0 230252 508088 231152
rect 0 225752 508088 226652
rect 0 221252 508088 222152
rect 0 216752 508088 217652
rect 0 212252 508088 213152
rect 0 207752 508088 208652
rect 0 203252 508088 204152
rect 0 198752 508088 199652
rect 0 194252 508088 195152
rect 0 189752 508088 190652
rect 0 185252 508088 186152
rect 0 180752 508088 181652
rect 0 176252 508088 177152
rect 0 171752 508088 172652
rect 0 167252 508088 168152
rect 0 162752 508088 163652
rect 0 158252 508088 159152
rect 0 153752 508088 154652
rect 0 149252 508088 150152
rect 0 144752 508088 145652
rect 0 140252 508088 141152
rect 0 135752 508088 136652
rect 0 131252 508088 132152
rect 0 126752 508088 127652
rect 0 122252 508088 123152
rect 0 117752 508088 118652
rect 0 113252 508088 114152
rect 0 108752 508088 109652
rect 0 104252 508088 105152
rect 0 99752 508088 100652
rect 0 95252 508088 96152
rect 0 90752 508088 91652
rect 0 86252 508088 87152
rect 0 81752 508088 82652
rect 0 77252 508088 78152
rect 0 72752 508088 73652
rect 0 68252 508088 69152
rect 0 63752 508088 64652
rect 0 59252 508088 60152
rect 0 54752 508088 55652
rect 0 50252 508088 51152
rect 0 45752 508088 46652
rect 0 41252 508088 42152
rect 0 36752 508088 37652
rect 0 32252 508088 33152
rect 0 27752 508088 28652
rect 0 23252 508088 24152
rect 1240 1252 506848 2152
rect 0 12 508088 912
<< obsm5 >>
rect 0 579872 900 579884
rect 0 578960 900 578972
rect 0 577412 920 578652
rect 507168 577412 508088 578652
rect 0 573472 508088 577412
rect 0 568972 508088 571932
rect 0 568652 900 568664
rect 0 567740 900 567752
rect 0 564472 508088 567432
rect 0 559972 508088 562932
rect 0 559652 900 559664
rect 0 558740 900 558752
rect 0 555472 508088 558432
rect 0 550972 508088 553932
rect 0 550652 900 550664
rect 0 549740 900 549752
rect 0 546472 508088 549432
rect 0 541972 508088 544932
rect 0 541652 900 541664
rect 0 540740 900 540752
rect 0 537472 508088 540432
rect 0 532972 508088 535932
rect 0 532652 900 532664
rect 0 531740 900 531752
rect 0 528472 508088 531432
rect 0 523972 508088 526932
rect 0 523652 900 523664
rect 0 522740 900 522752
rect 0 519472 508088 522432
rect 0 514972 508088 517932
rect 0 514652 900 514664
rect 0 513740 900 513752
rect 0 510472 508088 513432
rect 0 505972 508088 508932
rect 0 505652 900 505664
rect 0 504740 900 504752
rect 0 501472 508088 504432
rect 0 496972 508088 499932
rect 0 496652 900 496664
rect 0 495740 900 495752
rect 0 492472 508088 495432
rect 0 487972 508088 490932
rect 0 487652 900 487664
rect 0 486740 900 486752
rect 0 483472 508088 486432
rect 0 478972 508088 481932
rect 0 478652 900 478664
rect 0 477740 900 477752
rect 0 474472 508088 477432
rect 0 469972 508088 472932
rect 0 469652 900 469664
rect 0 468740 900 468752
rect 0 465472 508088 468432
rect 0 460972 508088 463932
rect 0 460652 900 460664
rect 0 459740 900 459752
rect 0 456472 508088 459432
rect 0 451972 508088 454932
rect 0 451652 900 451664
rect 0 450740 900 450752
rect 0 447472 508088 450432
rect 0 442972 508088 445932
rect 0 442652 900 442664
rect 0 441740 900 441752
rect 0 438472 508088 441432
rect 0 433972 508088 436932
rect 0 433652 900 433664
rect 0 432740 900 432752
rect 0 429472 508088 432432
rect 0 424972 508088 427932
rect 0 424652 900 424664
rect 0 423740 900 423752
rect 0 420472 508088 423432
rect 0 415972 508088 418932
rect 0 415652 900 415664
rect 0 414740 900 414752
rect 0 411472 508088 414432
rect 0 406972 508088 409932
rect 0 406652 900 406664
rect 0 405740 900 405752
rect 0 402472 508088 405432
rect 0 397972 508088 400932
rect 0 397652 900 397664
rect 0 396740 900 396752
rect 0 393472 508088 396432
rect 0 388972 508088 391932
rect 0 388652 900 388664
rect 0 387740 900 387752
rect 0 384472 508088 387432
rect 0 379972 508088 382932
rect 0 379652 900 379664
rect 0 378740 900 378752
rect 0 375472 508088 378432
rect 0 370972 508088 373932
rect 0 370652 900 370664
rect 0 369740 900 369752
rect 0 366472 508088 369432
rect 0 361972 508088 364932
rect 0 361652 900 361664
rect 0 360740 900 360752
rect 0 357472 508088 360432
rect 0 352972 508088 355932
rect 0 352652 900 352664
rect 0 351740 900 351752
rect 0 348472 508088 351432
rect 0 343972 508088 346932
rect 0 343652 900 343664
rect 0 342740 900 342752
rect 0 339472 508088 342432
rect 0 334972 508088 337932
rect 0 334652 900 334664
rect 0 333740 900 333752
rect 0 330472 508088 333432
rect 0 325972 508088 328932
rect 0 325652 900 325664
rect 0 324740 900 324752
rect 0 321472 508088 324432
rect 0 316972 508088 319932
rect 0 316652 900 316664
rect 0 315740 900 315752
rect 0 312472 508088 315432
rect 0 307972 508088 310932
rect 0 307652 900 307664
rect 0 306740 900 306752
rect 0 303472 508088 306432
rect 0 298972 508088 301932
rect 0 298652 900 298664
rect 0 297740 900 297752
rect 0 294472 508088 297432
rect 0 289972 508088 292932
rect 0 289652 900 289664
rect 0 288740 900 288752
rect 0 285472 508088 288432
rect 0 280972 508088 283932
rect 0 280652 900 280664
rect 0 279740 900 279752
rect 0 276472 508088 279432
rect 0 271972 508088 274932
rect 0 271652 900 271664
rect 0 270740 900 270752
rect 0 267472 508088 270432
rect 0 262972 508088 265932
rect 0 262652 900 262664
rect 0 261740 900 261752
rect 0 258472 508088 261432
rect 0 253972 508088 256932
rect 0 253652 900 253664
rect 0 252740 900 252752
rect 0 249472 508088 252432
rect 0 244972 508088 247932
rect 0 244652 900 244664
rect 0 243740 900 243752
rect 0 240472 508088 243432
rect 0 235972 508088 238932
rect 0 235652 900 235664
rect 0 234740 900 234752
rect 0 231472 508088 234432
rect 0 226972 508088 229932
rect 0 226652 900 226664
rect 0 225740 900 225752
rect 0 222472 508088 225432
rect 0 217972 508088 220932
rect 0 217652 900 217664
rect 0 216740 900 216752
rect 0 213472 508088 216432
rect 0 208972 508088 211932
rect 0 208652 900 208664
rect 0 207740 900 207752
rect 0 204472 508088 207432
rect 0 199972 508088 202932
rect 0 199652 900 199664
rect 0 198740 900 198752
rect 0 195472 508088 198432
rect 0 190972 508088 193932
rect 0 190652 900 190664
rect 0 189740 900 189752
rect 0 186472 508088 189432
rect 0 181972 508088 184932
rect 0 181652 900 181664
rect 0 180740 900 180752
rect 0 177472 508088 180432
rect 0 172972 508088 175932
rect 0 172652 900 172664
rect 0 171740 900 171752
rect 0 168472 508088 171432
rect 0 163972 508088 166932
rect 0 163652 900 163664
rect 0 162740 900 162752
rect 0 159472 508088 162432
rect 0 154972 508088 157932
rect 0 154652 900 154664
rect 0 153740 900 153752
rect 0 150472 508088 153432
rect 0 145972 508088 148932
rect 0 145652 900 145664
rect 0 144740 900 144752
rect 0 141472 508088 144432
rect 0 136972 508088 139932
rect 0 136652 900 136664
rect 0 135740 900 135752
rect 0 132472 508088 135432
rect 0 127972 508088 130932
rect 0 127652 900 127664
rect 0 126740 900 126752
rect 0 123472 508088 126432
rect 0 118972 508088 121932
rect 0 118652 900 118664
rect 0 117740 900 117752
rect 0 114472 508088 117432
rect 0 109972 508088 112932
rect 0 109652 900 109664
rect 0 108740 900 108752
rect 0 105472 508088 108432
rect 0 100972 508088 103932
rect 0 100652 900 100664
rect 0 99740 900 99752
rect 0 96472 508088 99432
rect 0 91972 508088 94932
rect 0 91652 900 91664
rect 0 90740 900 90752
rect 0 87472 508088 90432
rect 0 82972 508088 85932
rect 0 82652 900 82664
rect 0 81740 900 81752
rect 0 78472 508088 81432
rect 0 73972 508088 76932
rect 0 73652 900 73664
rect 0 72740 900 72752
rect 0 69472 508088 72432
rect 0 64972 508088 67932
rect 0 64652 900 64664
rect 0 63740 900 63752
rect 0 60472 508088 63432
rect 0 55972 508088 58932
rect 0 55652 900 55664
rect 0 54740 900 54752
rect 0 51472 508088 54432
rect 0 46972 508088 49932
rect 0 46652 900 46664
rect 0 45740 900 45752
rect 0 42472 508088 45432
rect 0 37972 508088 40932
rect 0 37652 900 37664
rect 0 36740 900 36752
rect 0 33472 508088 36432
rect 0 28972 508088 31932
rect 0 28652 900 28664
rect 0 27740 900 27752
rect 0 24472 508088 27432
rect 0 2472 508088 22932
rect 0 1232 920 2472
rect 507168 1232 508088 2472
rect 0 912 900 924
rect 0 0 900 12
<< labels >>
rlabel metal3 s 4586 72486 5386 72606 6 IO_ISOL_N
port 1 nsew signal input
rlabel metal3 s 4586 33046 5386 33166 6 Test_en
port 2 nsew signal input
rlabel metal3 s 502786 540462 503586 540582 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 4586 13326 5386 13446 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 4586 52766 5386 52886 6 clk
port 5 nsew signal input
rlabel metal2 s 13804 575726 13860 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 6 nsew signal output
rlabel metal3 s 502786 110838 503586 110958 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
port 7 nsew signal output
rlabel metal3 s 502786 182374 503586 182494 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
port 8 nsew signal output
rlabel metal3 s 502786 254046 503586 254166 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
port 9 nsew signal output
rlabel metal3 s 502786 325718 503586 325838 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
port 10 nsew signal output
rlabel metal3 s 502786 397254 503586 397374 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
port 11 nsew signal output
rlabel metal3 s 502786 468926 503586 469046 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
port 12 nsew signal output
rlabel metal2 s 442340 3526 442396 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
port 13 nsew signal output
rlabel metal2 s 444640 3526 444696 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
port 14 nsew signal output
rlabel metal2 s 446940 3526 446996 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
port 15 nsew signal output
rlabel metal2 s 449240 3526 449296 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
port 16 nsew signal output
rlabel metal2 s 32204 575726 32260 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 17 nsew signal output
rlabel metal2 s 451540 3526 451596 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
port 18 nsew signal output
rlabel metal2 s 453840 3526 453896 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
port 19 nsew signal output
rlabel metal2 s 456140 3526 456196 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
port 20 nsew signal output
rlabel metal2 s 458440 3526 458496 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
port 21 nsew signal output
rlabel metal2 s 460740 3526 460796 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
port 22 nsew signal output
rlabel metal2 s 379964 3526 380020 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
port 23 nsew signal output
rlabel metal2 s 382264 3526 382320 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
port 24 nsew signal output
rlabel metal2 s 384564 3526 384620 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
port 25 nsew signal output
rlabel metal2 s 386864 3526 386920 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
port 26 nsew signal output
rlabel metal2 s 389164 3526 389220 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
port 27 nsew signal output
rlabel metal2 s 50696 575726 50752 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 28 nsew signal output
rlabel metal2 s 391464 3526 391520 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
port 29 nsew signal output
rlabel metal2 s 393764 3526 393820 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
port 30 nsew signal output
rlabel metal2 s 396064 3526 396120 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
port 31 nsew signal output
rlabel metal2 s 398364 3526 398420 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
port 32 nsew signal output
rlabel metal2 s 317588 3526 317644 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
port 33 nsew signal output
rlabel metal2 s 319888 3526 319944 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
port 34 nsew signal output
rlabel metal2 s 322188 3526 322244 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
port 35 nsew signal output
rlabel metal2 s 324488 3526 324544 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
port 36 nsew signal output
rlabel metal2 s 326788 3526 326844 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
port 37 nsew signal output
rlabel metal2 s 329088 3526 329144 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
port 38 nsew signal output
rlabel metal2 s 69188 575726 69244 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 39 nsew signal output
rlabel metal2 s 331388 3526 331444 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
port 40 nsew signal output
rlabel metal2 s 333688 3526 333744 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
port 41 nsew signal output
rlabel metal2 s 335988 3526 336044 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
port 42 nsew signal output
rlabel metal2 s 255212 3526 255268 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
port 43 nsew signal output
rlabel metal2 s 257512 3526 257568 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
port 44 nsew signal output
rlabel metal2 s 259812 3526 259868 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
port 45 nsew signal output
rlabel metal2 s 262112 3526 262168 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
port 46 nsew signal output
rlabel metal2 s 264412 3526 264468 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
port 47 nsew signal output
rlabel metal2 s 266712 3526 266768 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
port 48 nsew signal output
rlabel metal2 s 269012 3526 269068 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
port 49 nsew signal output
rlabel metal2 s 87680 575726 87736 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 50 nsew signal output
rlabel metal2 s 271312 3526 271368 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
port 51 nsew signal output
rlabel metal2 s 273612 3526 273668 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
port 52 nsew signal output
rlabel metal2 s 192836 3526 192892 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
port 53 nsew signal output
rlabel metal2 s 195136 3526 195192 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
port 54 nsew signal output
rlabel metal2 s 197436 3526 197492 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
port 55 nsew signal output
rlabel metal2 s 199736 3526 199792 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
port 56 nsew signal output
rlabel metal2 s 202036 3526 202092 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
port 57 nsew signal output
rlabel metal2 s 204336 3526 204392 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
port 58 nsew signal output
rlabel metal2 s 206636 3526 206692 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
port 59 nsew signal output
rlabel metal2 s 208936 3526 208992 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
port 60 nsew signal output
rlabel metal2 s 106172 575726 106228 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 61 nsew signal output
rlabel metal2 s 211236 3526 211292 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
port 62 nsew signal output
rlabel metal2 s 130460 3526 130516 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
port 63 nsew signal output
rlabel metal2 s 132760 3526 132816 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
port 64 nsew signal output
rlabel metal2 s 135060 3526 135116 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
port 65 nsew signal output
rlabel metal2 s 137360 3526 137416 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
port 66 nsew signal output
rlabel metal2 s 139660 3526 139716 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
port 67 nsew signal output
rlabel metal2 s 141960 3526 142016 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
port 68 nsew signal output
rlabel metal2 s 144260 3526 144316 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
port 69 nsew signal output
rlabel metal2 s 146560 3526 146616 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
port 70 nsew signal output
rlabel metal2 s 148860 3526 148916 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
port 71 nsew signal output
rlabel metal2 s 124664 575726 124720 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 72 nsew signal output
rlabel metal2 s 68084 3526 68140 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
port 73 nsew signal output
rlabel metal2 s 70384 3526 70440 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
port 74 nsew signal output
rlabel metal2 s 72684 3526 72740 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
port 75 nsew signal output
rlabel metal2 s 74984 3526 75040 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
port 76 nsew signal output
rlabel metal2 s 77284 3526 77340 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
port 77 nsew signal output
rlabel metal2 s 79584 3526 79640 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
port 78 nsew signal output
rlabel metal2 s 81884 3526 81940 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
port 79 nsew signal output
rlabel metal2 s 84184 3526 84240 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
port 80 nsew signal output
rlabel metal2 s 86484 3526 86540 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
port 81 nsew signal output
rlabel metal2 s 5708 3526 5764 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
port 82 nsew signal output
rlabel metal2 s 143156 575726 143212 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 83 nsew signal output
rlabel metal2 s 8008 3526 8064 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
port 84 nsew signal output
rlabel metal2 s 10308 3526 10364 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
port 85 nsew signal output
rlabel metal2 s 12608 3526 12664 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
port 86 nsew signal output
rlabel metal2 s 14908 3526 14964 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
port 87 nsew signal output
rlabel metal2 s 17208 3526 17264 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
port 88 nsew signal output
rlabel metal2 s 19508 3526 19564 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
port 89 nsew signal output
rlabel metal2 s 21808 3526 21864 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
port 90 nsew signal output
rlabel metal2 s 24108 3526 24164 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
port 91 nsew signal output
rlabel metal3 s 4586 92342 5386 92462 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
port 92 nsew signal output
rlabel metal3 s 4586 151502 5386 151622 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
port 93 nsew signal output
rlabel metal2 s 161648 575726 161704 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 94 nsew signal output
rlabel metal3 s 4586 210798 5386 210918 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
port 95 nsew signal output
rlabel metal3 s 4586 270094 5386 270214 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
port 96 nsew signal output
rlabel metal3 s 4586 329390 5386 329510 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
port 97 nsew signal output
rlabel metal3 s 4586 388686 5386 388806 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
port 98 nsew signal output
rlabel metal3 s 4586 447982 5386 448102 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
port 99 nsew signal output
rlabel metal3 s 4586 507142 5386 507262 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
port 100 nsew signal output
rlabel metal3 s 502786 39166 503586 39286 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
port 101 nsew signal output
rlabel metal2 s 180140 575726 180196 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 102 nsew signal input
rlabel metal3 s 502786 134638 503586 134758 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
port 103 nsew signal input
rlabel metal3 s 502786 206310 503586 206430 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
port 104 nsew signal input
rlabel metal3 s 502786 277846 503586 277966 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
port 105 nsew signal input
rlabel metal3 s 502786 349518 503586 349638 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
port 106 nsew signal input
rlabel metal3 s 502786 421190 503586 421310 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
port 107 nsew signal input
rlabel metal3 s 502786 492726 503586 492846 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
port 108 nsew signal input
rlabel metal2 s 463132 3526 463188 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
port 109 nsew signal input
rlabel metal2 s 465432 3526 465488 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
port 110 nsew signal input
rlabel metal2 s 467732 3526 467788 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
port 111 nsew signal input
rlabel metal2 s 470032 3526 470088 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
port 112 nsew signal input
rlabel metal2 s 198540 575726 198596 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 113 nsew signal input
rlabel metal2 s 472332 3526 472388 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
port 114 nsew signal input
rlabel metal2 s 474632 3526 474688 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
port 115 nsew signal input
rlabel metal2 s 476932 3526 476988 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
port 116 nsew signal input
rlabel metal2 s 479232 3526 479288 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
port 117 nsew signal input
rlabel metal2 s 481532 3526 481588 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
port 118 nsew signal input
rlabel metal2 s 400756 3526 400812 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
port 119 nsew signal input
rlabel metal2 s 403056 3526 403112 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
port 120 nsew signal input
rlabel metal2 s 405356 3526 405412 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
port 121 nsew signal input
rlabel metal2 s 407656 3526 407712 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
port 122 nsew signal input
rlabel metal2 s 409956 3526 410012 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
port 123 nsew signal input
rlabel metal2 s 217032 575726 217088 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 124 nsew signal input
rlabel metal2 s 412256 3526 412312 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
port 125 nsew signal input
rlabel metal2 s 414556 3526 414612 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
port 126 nsew signal input
rlabel metal2 s 416856 3526 416912 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
port 127 nsew signal input
rlabel metal2 s 419156 3526 419212 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
port 128 nsew signal input
rlabel metal2 s 338380 3526 338436 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
port 129 nsew signal input
rlabel metal2 s 340680 3526 340736 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
port 130 nsew signal input
rlabel metal2 s 342980 3526 343036 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
port 131 nsew signal input
rlabel metal2 s 345280 3526 345336 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
port 132 nsew signal input
rlabel metal2 s 347580 3526 347636 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
port 133 nsew signal input
rlabel metal2 s 349880 3526 349936 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
port 134 nsew signal input
rlabel metal2 s 235524 575726 235580 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 135 nsew signal input
rlabel metal2 s 352180 3526 352236 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
port 136 nsew signal input
rlabel metal2 s 354480 3526 354536 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
port 137 nsew signal input
rlabel metal2 s 356780 3526 356836 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
port 138 nsew signal input
rlabel metal2 s 276004 3526 276060 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
port 139 nsew signal input
rlabel metal2 s 278304 3526 278360 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
port 140 nsew signal input
rlabel metal2 s 280604 3526 280660 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
port 141 nsew signal input
rlabel metal2 s 282904 3526 282960 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
port 142 nsew signal input
rlabel metal2 s 285204 3526 285260 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
port 143 nsew signal input
rlabel metal2 s 287504 3526 287560 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
port 144 nsew signal input
rlabel metal2 s 289804 3526 289860 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
port 145 nsew signal input
rlabel metal2 s 254016 575726 254072 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 146 nsew signal input
rlabel metal2 s 292104 3526 292160 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
port 147 nsew signal input
rlabel metal2 s 294404 3526 294460 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
port 148 nsew signal input
rlabel metal2 s 213628 3526 213684 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
port 149 nsew signal input
rlabel metal2 s 215928 3526 215984 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
port 150 nsew signal input
rlabel metal2 s 218228 3526 218284 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
port 151 nsew signal input
rlabel metal2 s 220528 3526 220584 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
port 152 nsew signal input
rlabel metal2 s 222828 3526 222884 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
port 153 nsew signal input
rlabel metal2 s 225128 3526 225184 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
port 154 nsew signal input
rlabel metal2 s 227428 3526 227484 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
port 155 nsew signal input
rlabel metal2 s 229728 3526 229784 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
port 156 nsew signal input
rlabel metal2 s 272508 575726 272564 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 157 nsew signal input
rlabel metal2 s 232028 3526 232084 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
port 158 nsew signal input
rlabel metal2 s 151252 3526 151308 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
port 159 nsew signal input
rlabel metal2 s 153552 3526 153608 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
port 160 nsew signal input
rlabel metal2 s 155852 3526 155908 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
port 161 nsew signal input
rlabel metal2 s 158152 3526 158208 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
port 162 nsew signal input
rlabel metal2 s 160452 3526 160508 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
port 163 nsew signal input
rlabel metal2 s 162752 3526 162808 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
port 164 nsew signal input
rlabel metal2 s 165052 3526 165108 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
port 165 nsew signal input
rlabel metal2 s 167352 3526 167408 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
port 166 nsew signal input
rlabel metal2 s 169652 3526 169708 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
port 167 nsew signal input
rlabel metal2 s 291000 575726 291056 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 168 nsew signal input
rlabel metal2 s 88876 3526 88932 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
port 169 nsew signal input
rlabel metal2 s 91176 3526 91232 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
port 170 nsew signal input
rlabel metal2 s 93476 3526 93532 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
port 171 nsew signal input
rlabel metal2 s 95776 3526 95832 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
port 172 nsew signal input
rlabel metal2 s 98076 3526 98132 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
port 173 nsew signal input
rlabel metal2 s 100376 3526 100432 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
port 174 nsew signal input
rlabel metal2 s 102676 3526 102732 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
port 175 nsew signal input
rlabel metal2 s 104976 3526 105032 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
port 176 nsew signal input
rlabel metal2 s 107276 3526 107332 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
port 177 nsew signal input
rlabel metal2 s 26500 3526 26556 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
port 178 nsew signal input
rlabel metal2 s 309492 575726 309548 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 179 nsew signal input
rlabel metal2 s 28800 3526 28856 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
port 180 nsew signal input
rlabel metal2 s 31100 3526 31156 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
port 181 nsew signal input
rlabel metal2 s 33400 3526 33456 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
port 182 nsew signal input
rlabel metal2 s 35700 3526 35756 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
port 183 nsew signal input
rlabel metal2 s 38000 3526 38056 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
port 184 nsew signal input
rlabel metal2 s 40300 3526 40356 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
port 185 nsew signal input
rlabel metal2 s 42600 3526 42656 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
port 186 nsew signal input
rlabel metal2 s 44900 3526 44956 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
port 187 nsew signal input
rlabel metal3 s 4586 112062 5386 112182 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
port 188 nsew signal input
rlabel metal3 s 4586 171358 5386 171478 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
port 189 nsew signal input
rlabel metal2 s 327984 575726 328040 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 190 nsew signal input
rlabel metal3 s 4586 230654 5386 230774 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
port 191 nsew signal input
rlabel metal3 s 4586 289814 5386 289934 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
port 192 nsew signal input
rlabel metal3 s 4586 349110 5386 349230 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
port 193 nsew signal input
rlabel metal3 s 4586 408406 5386 408526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
port 194 nsew signal input
rlabel metal3 s 4586 467702 5386 467822 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
port 195 nsew signal input
rlabel metal3 s 4586 526998 5386 527118 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
port 196 nsew signal input
rlabel metal3 s 502786 63102 503586 63222 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
port 197 nsew signal input
rlabel metal2 s 346476 575726 346532 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 198 nsew signal output
rlabel metal3 s 502786 158574 503586 158694 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
port 199 nsew signal output
rlabel metal3 s 502786 230110 503586 230230 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
port 200 nsew signal output
rlabel metal3 s 502786 301782 503586 301902 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
port 201 nsew signal output
rlabel metal3 s 502786 373454 503586 373574 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
port 202 nsew signal output
rlabel metal3 s 502786 444990 503586 445110 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
port 203 nsew signal output
rlabel metal3 s 502786 516662 503586 516782 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
port 204 nsew signal output
rlabel metal2 s 483924 3526 483980 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
port 205 nsew signal output
rlabel metal2 s 486224 3526 486280 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
port 206 nsew signal output
rlabel metal2 s 488524 3526 488580 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
port 207 nsew signal output
rlabel metal2 s 490824 3526 490880 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
port 208 nsew signal output
rlabel metal2 s 364876 575726 364932 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 209 nsew signal output
rlabel metal2 s 493124 3526 493180 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
port 210 nsew signal output
rlabel metal2 s 495424 3526 495480 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
port 211 nsew signal output
rlabel metal2 s 497724 3526 497780 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
port 212 nsew signal output
rlabel metal2 s 500024 3526 500080 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
port 213 nsew signal output
rlabel metal2 s 502324 3526 502380 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
port 214 nsew signal output
rlabel metal2 s 421548 3526 421604 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
port 215 nsew signal output
rlabel metal2 s 423848 3526 423904 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
port 216 nsew signal output
rlabel metal2 s 426148 3526 426204 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
port 217 nsew signal output
rlabel metal2 s 428448 3526 428504 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
port 218 nsew signal output
rlabel metal2 s 430748 3526 430804 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
port 219 nsew signal output
rlabel metal2 s 383368 575726 383424 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 220 nsew signal output
rlabel metal2 s 433048 3526 433104 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
port 221 nsew signal output
rlabel metal2 s 435348 3526 435404 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
port 222 nsew signal output
rlabel metal2 s 437648 3526 437704 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
port 223 nsew signal output
rlabel metal2 s 439948 3526 440004 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
port 224 nsew signal output
rlabel metal2 s 359172 3526 359228 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
port 225 nsew signal output
rlabel metal2 s 361472 3526 361528 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
port 226 nsew signal output
rlabel metal2 s 363772 3526 363828 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
port 227 nsew signal output
rlabel metal2 s 366072 3526 366128 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
port 228 nsew signal output
rlabel metal2 s 368372 3526 368428 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
port 229 nsew signal output
rlabel metal2 s 370672 3526 370728 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
port 230 nsew signal output
rlabel metal2 s 401860 575726 401916 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 231 nsew signal output
rlabel metal2 s 372972 3526 373028 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
port 232 nsew signal output
rlabel metal2 s 375272 3526 375328 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
port 233 nsew signal output
rlabel metal2 s 377572 3526 377628 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
port 234 nsew signal output
rlabel metal2 s 296796 3526 296852 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
port 235 nsew signal output
rlabel metal2 s 299096 3526 299152 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
port 236 nsew signal output
rlabel metal2 s 301396 3526 301452 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
port 237 nsew signal output
rlabel metal2 s 303696 3526 303752 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
port 238 nsew signal output
rlabel metal2 s 305996 3526 306052 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
port 239 nsew signal output
rlabel metal2 s 308296 3526 308352 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
port 240 nsew signal output
rlabel metal2 s 310596 3526 310652 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
port 241 nsew signal output
rlabel metal2 s 420352 575726 420408 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 242 nsew signal output
rlabel metal2 s 312896 3526 312952 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
port 243 nsew signal output
rlabel metal2 s 315196 3526 315252 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
port 244 nsew signal output
rlabel metal2 s 234420 3526 234476 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
port 245 nsew signal output
rlabel metal2 s 236720 3526 236776 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
port 246 nsew signal output
rlabel metal2 s 239020 3526 239076 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
port 247 nsew signal output
rlabel metal2 s 241320 3526 241376 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
port 248 nsew signal output
rlabel metal2 s 243620 3526 243676 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
port 249 nsew signal output
rlabel metal2 s 245920 3526 245976 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
port 250 nsew signal output
rlabel metal2 s 248220 3526 248276 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
port 251 nsew signal output
rlabel metal2 s 250520 3526 250576 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
port 252 nsew signal output
rlabel metal2 s 438844 575726 438900 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 253 nsew signal output
rlabel metal2 s 252820 3526 252876 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
port 254 nsew signal output
rlabel metal2 s 172044 3526 172100 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
port 255 nsew signal output
rlabel metal2 s 174344 3526 174400 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
port 256 nsew signal output
rlabel metal2 s 176644 3526 176700 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
port 257 nsew signal output
rlabel metal2 s 178944 3526 179000 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
port 258 nsew signal output
rlabel metal2 s 181244 3526 181300 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
port 259 nsew signal output
rlabel metal2 s 183544 3526 183600 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
port 260 nsew signal output
rlabel metal2 s 185844 3526 185900 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
port 261 nsew signal output
rlabel metal2 s 188144 3526 188200 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
port 262 nsew signal output
rlabel metal2 s 190444 3526 190500 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
port 263 nsew signal output
rlabel metal2 s 457336 575726 457392 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 264 nsew signal output
rlabel metal2 s 109668 3526 109724 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
port 265 nsew signal output
rlabel metal2 s 111968 3526 112024 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
port 266 nsew signal output
rlabel metal2 s 114268 3526 114324 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
port 267 nsew signal output
rlabel metal2 s 116568 3526 116624 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
port 268 nsew signal output
rlabel metal2 s 118868 3526 118924 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
port 269 nsew signal output
rlabel metal2 s 121168 3526 121224 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
port 270 nsew signal output
rlabel metal2 s 123468 3526 123524 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
port 271 nsew signal output
rlabel metal2 s 125768 3526 125824 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
port 272 nsew signal output
rlabel metal2 s 128068 3526 128124 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
port 273 nsew signal output
rlabel metal2 s 47292 3526 47348 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
port 274 nsew signal output
rlabel metal2 s 475828 575726 475884 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 275 nsew signal output
rlabel metal2 s 49592 3526 49648 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
port 276 nsew signal output
rlabel metal2 s 51892 3526 51948 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
port 277 nsew signal output
rlabel metal2 s 54192 3526 54248 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
port 278 nsew signal output
rlabel metal2 s 56492 3526 56548 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
port 279 nsew signal output
rlabel metal2 s 58792 3526 58848 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
port 280 nsew signal output
rlabel metal2 s 61092 3526 61148 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
port 281 nsew signal output
rlabel metal2 s 63392 3526 63448 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
port 282 nsew signal output
rlabel metal2 s 65692 3526 65748 4326 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
port 283 nsew signal output
rlabel metal3 s 4586 131782 5386 131902 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
port 284 nsew signal output
rlabel metal3 s 4586 191078 5386 191198 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
port 285 nsew signal output
rlabel metal2 s 494320 575726 494376 576526 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 286 nsew signal output
rlabel metal3 s 4586 250374 5386 250494 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
port 287 nsew signal output
rlabel metal3 s 4586 309670 5386 309790 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
port 288 nsew signal output
rlabel metal3 s 4586 368830 5386 368950 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
port 289 nsew signal output
rlabel metal3 s 4586 428126 5386 428246 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
port 290 nsew signal output
rlabel metal3 s 4586 487422 5386 487542 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
port 291 nsew signal output
rlabel metal3 s 4586 546718 5386 546838 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
port 292 nsew signal output
rlabel metal3 s 502786 86902 503586 87022 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
port 293 nsew signal output
rlabel metal3 s 502786 15366 503586 15486 6 prog_clk
port 294 nsew signal input
rlabel metal3 s 4586 566438 5386 566558 6 sc_head
port 295 nsew signal input
rlabel metal3 s 502786 564398 503586 564518 6 sc_tail
port 296 nsew signal output
rlabel metal4 s 505948 1252 506848 578632 6 VPWR
port 297 nsew power bidirectional
rlabel metal4 s 1240 1252 2140 578632 6 VPWR
port 298 nsew power bidirectional
rlabel metal5 s 1240 577732 506848 578632 6 VPWR
port 299 nsew power bidirectional
rlabel metal5 s 0 572252 508088 573152 6 VPWR
port 300 nsew power bidirectional
rlabel metal5 s 0 563252 508088 564152 6 VPWR
port 301 nsew power bidirectional
rlabel metal5 s 0 554252 508088 555152 6 VPWR
port 302 nsew power bidirectional
rlabel metal5 s 0 545252 508088 546152 6 VPWR
port 303 nsew power bidirectional
rlabel metal5 s 0 536252 508088 537152 6 VPWR
port 304 nsew power bidirectional
rlabel metal5 s 0 527252 508088 528152 6 VPWR
port 305 nsew power bidirectional
rlabel metal5 s 0 518252 508088 519152 6 VPWR
port 306 nsew power bidirectional
rlabel metal5 s 0 509252 508088 510152 6 VPWR
port 307 nsew power bidirectional
rlabel metal5 s 0 500252 508088 501152 6 VPWR
port 308 nsew power bidirectional
rlabel metal5 s 0 491252 508088 492152 6 VPWR
port 309 nsew power bidirectional
rlabel metal5 s 0 482252 508088 483152 6 VPWR
port 310 nsew power bidirectional
rlabel metal5 s 0 473252 508088 474152 6 VPWR
port 311 nsew power bidirectional
rlabel metal5 s 0 464252 508088 465152 6 VPWR
port 312 nsew power bidirectional
rlabel metal5 s 0 455252 508088 456152 6 VPWR
port 313 nsew power bidirectional
rlabel metal5 s 0 446252 508088 447152 6 VPWR
port 314 nsew power bidirectional
rlabel metal5 s 0 437252 508088 438152 6 VPWR
port 315 nsew power bidirectional
rlabel metal5 s 0 428252 508088 429152 6 VPWR
port 316 nsew power bidirectional
rlabel metal5 s 0 419252 508088 420152 6 VPWR
port 317 nsew power bidirectional
rlabel metal5 s 0 410252 508088 411152 6 VPWR
port 318 nsew power bidirectional
rlabel metal5 s 0 401252 508088 402152 6 VPWR
port 319 nsew power bidirectional
rlabel metal5 s 0 392252 508088 393152 6 VPWR
port 320 nsew power bidirectional
rlabel metal5 s 0 383252 508088 384152 6 VPWR
port 321 nsew power bidirectional
rlabel metal5 s 0 374252 508088 375152 6 VPWR
port 322 nsew power bidirectional
rlabel metal5 s 0 365252 508088 366152 6 VPWR
port 323 nsew power bidirectional
rlabel metal5 s 0 356252 508088 357152 6 VPWR
port 324 nsew power bidirectional
rlabel metal5 s 0 347252 508088 348152 6 VPWR
port 325 nsew power bidirectional
rlabel metal5 s 0 338252 508088 339152 6 VPWR
port 326 nsew power bidirectional
rlabel metal5 s 0 329252 508088 330152 6 VPWR
port 327 nsew power bidirectional
rlabel metal5 s 0 320252 508088 321152 6 VPWR
port 328 nsew power bidirectional
rlabel metal5 s 0 311252 508088 312152 6 VPWR
port 329 nsew power bidirectional
rlabel metal5 s 0 302252 508088 303152 6 VPWR
port 330 nsew power bidirectional
rlabel metal5 s 0 293252 508088 294152 6 VPWR
port 331 nsew power bidirectional
rlabel metal5 s 0 284252 508088 285152 6 VPWR
port 332 nsew power bidirectional
rlabel metal5 s 0 275252 508088 276152 6 VPWR
port 333 nsew power bidirectional
rlabel metal5 s 0 266252 508088 267152 6 VPWR
port 334 nsew power bidirectional
rlabel metal5 s 0 257252 508088 258152 6 VPWR
port 335 nsew power bidirectional
rlabel metal5 s 0 248252 508088 249152 6 VPWR
port 336 nsew power bidirectional
rlabel metal5 s 0 239252 508088 240152 6 VPWR
port 337 nsew power bidirectional
rlabel metal5 s 0 230252 508088 231152 6 VPWR
port 338 nsew power bidirectional
rlabel metal5 s 0 221252 508088 222152 6 VPWR
port 339 nsew power bidirectional
rlabel metal5 s 0 212252 508088 213152 6 VPWR
port 340 nsew power bidirectional
rlabel metal5 s 0 203252 508088 204152 6 VPWR
port 341 nsew power bidirectional
rlabel metal5 s 0 194252 508088 195152 6 VPWR
port 342 nsew power bidirectional
rlabel metal5 s 0 185252 508088 186152 6 VPWR
port 343 nsew power bidirectional
rlabel metal5 s 0 176252 508088 177152 6 VPWR
port 344 nsew power bidirectional
rlabel metal5 s 0 167252 508088 168152 6 VPWR
port 345 nsew power bidirectional
rlabel metal5 s 0 158252 508088 159152 6 VPWR
port 346 nsew power bidirectional
rlabel metal5 s 0 149252 508088 150152 6 VPWR
port 347 nsew power bidirectional
rlabel metal5 s 0 140252 508088 141152 6 VPWR
port 348 nsew power bidirectional
rlabel metal5 s 0 131252 508088 132152 6 VPWR
port 349 nsew power bidirectional
rlabel metal5 s 0 122252 508088 123152 6 VPWR
port 350 nsew power bidirectional
rlabel metal5 s 0 113252 508088 114152 6 VPWR
port 351 nsew power bidirectional
rlabel metal5 s 0 104252 508088 105152 6 VPWR
port 352 nsew power bidirectional
rlabel metal5 s 0 95252 508088 96152 6 VPWR
port 353 nsew power bidirectional
rlabel metal5 s 0 86252 508088 87152 6 VPWR
port 354 nsew power bidirectional
rlabel metal5 s 0 77252 508088 78152 6 VPWR
port 355 nsew power bidirectional
rlabel metal5 s 0 68252 508088 69152 6 VPWR
port 356 nsew power bidirectional
rlabel metal5 s 0 59252 508088 60152 6 VPWR
port 357 nsew power bidirectional
rlabel metal5 s 0 50252 508088 51152 6 VPWR
port 358 nsew power bidirectional
rlabel metal5 s 0 41252 508088 42152 6 VPWR
port 359 nsew power bidirectional
rlabel metal5 s 0 32252 508088 33152 6 VPWR
port 360 nsew power bidirectional
rlabel metal5 s 0 23252 508088 24152 6 VPWR
port 361 nsew power bidirectional
rlabel metal5 s 1240 1252 506848 2152 6 VPWR
port 362 nsew power bidirectional
rlabel metal4 s 507188 12 508088 579872 6 VGND
port 363 nsew ground bidirectional
rlabel metal4 s 0 12 900 579872 6 VGND
port 364 nsew ground bidirectional
rlabel metal5 s 0 578972 508088 579872 6 VGND
port 365 nsew ground bidirectional
rlabel metal5 s 0 567752 508088 568652 6 VGND
port 366 nsew ground bidirectional
rlabel metal5 s 0 558752 508088 559652 6 VGND
port 367 nsew ground bidirectional
rlabel metal5 s 0 549752 508088 550652 6 VGND
port 368 nsew ground bidirectional
rlabel metal5 s 0 540752 508088 541652 6 VGND
port 369 nsew ground bidirectional
rlabel metal5 s 0 531752 508088 532652 6 VGND
port 370 nsew ground bidirectional
rlabel metal5 s 0 522752 508088 523652 6 VGND
port 371 nsew ground bidirectional
rlabel metal5 s 0 513752 508088 514652 6 VGND
port 372 nsew ground bidirectional
rlabel metal5 s 0 504752 508088 505652 6 VGND
port 373 nsew ground bidirectional
rlabel metal5 s 0 495752 508088 496652 6 VGND
port 374 nsew ground bidirectional
rlabel metal5 s 0 486752 508088 487652 6 VGND
port 375 nsew ground bidirectional
rlabel metal5 s 0 477752 508088 478652 6 VGND
port 376 nsew ground bidirectional
rlabel metal5 s 0 468752 508088 469652 6 VGND
port 377 nsew ground bidirectional
rlabel metal5 s 0 459752 508088 460652 6 VGND
port 378 nsew ground bidirectional
rlabel metal5 s 0 450752 508088 451652 6 VGND
port 379 nsew ground bidirectional
rlabel metal5 s 0 441752 508088 442652 6 VGND
port 380 nsew ground bidirectional
rlabel metal5 s 0 432752 508088 433652 6 VGND
port 381 nsew ground bidirectional
rlabel metal5 s 0 423752 508088 424652 6 VGND
port 382 nsew ground bidirectional
rlabel metal5 s 0 414752 508088 415652 6 VGND
port 383 nsew ground bidirectional
rlabel metal5 s 0 405752 508088 406652 6 VGND
port 384 nsew ground bidirectional
rlabel metal5 s 0 396752 508088 397652 6 VGND
port 385 nsew ground bidirectional
rlabel metal5 s 0 387752 508088 388652 6 VGND
port 386 nsew ground bidirectional
rlabel metal5 s 0 378752 508088 379652 6 VGND
port 387 nsew ground bidirectional
rlabel metal5 s 0 369752 508088 370652 6 VGND
port 388 nsew ground bidirectional
rlabel metal5 s 0 360752 508088 361652 6 VGND
port 389 nsew ground bidirectional
rlabel metal5 s 0 351752 508088 352652 6 VGND
port 390 nsew ground bidirectional
rlabel metal5 s 0 342752 508088 343652 6 VGND
port 391 nsew ground bidirectional
rlabel metal5 s 0 333752 508088 334652 6 VGND
port 392 nsew ground bidirectional
rlabel metal5 s 0 324752 508088 325652 6 VGND
port 393 nsew ground bidirectional
rlabel metal5 s 0 315752 508088 316652 6 VGND
port 394 nsew ground bidirectional
rlabel metal5 s 0 306752 508088 307652 6 VGND
port 395 nsew ground bidirectional
rlabel metal5 s 0 297752 508088 298652 6 VGND
port 396 nsew ground bidirectional
rlabel metal5 s 0 288752 508088 289652 6 VGND
port 397 nsew ground bidirectional
rlabel metal5 s 0 279752 508088 280652 6 VGND
port 398 nsew ground bidirectional
rlabel metal5 s 0 270752 508088 271652 6 VGND
port 399 nsew ground bidirectional
rlabel metal5 s 0 261752 508088 262652 6 VGND
port 400 nsew ground bidirectional
rlabel metal5 s 0 252752 508088 253652 6 VGND
port 401 nsew ground bidirectional
rlabel metal5 s 0 243752 508088 244652 6 VGND
port 402 nsew ground bidirectional
rlabel metal5 s 0 234752 508088 235652 6 VGND
port 403 nsew ground bidirectional
rlabel metal5 s 0 225752 508088 226652 6 VGND
port 404 nsew ground bidirectional
rlabel metal5 s 0 216752 508088 217652 6 VGND
port 405 nsew ground bidirectional
rlabel metal5 s 0 207752 508088 208652 6 VGND
port 406 nsew ground bidirectional
rlabel metal5 s 0 198752 508088 199652 6 VGND
port 407 nsew ground bidirectional
rlabel metal5 s 0 189752 508088 190652 6 VGND
port 408 nsew ground bidirectional
rlabel metal5 s 0 180752 508088 181652 6 VGND
port 409 nsew ground bidirectional
rlabel metal5 s 0 171752 508088 172652 6 VGND
port 410 nsew ground bidirectional
rlabel metal5 s 0 162752 508088 163652 6 VGND
port 411 nsew ground bidirectional
rlabel metal5 s 0 153752 508088 154652 6 VGND
port 412 nsew ground bidirectional
rlabel metal5 s 0 144752 508088 145652 6 VGND
port 413 nsew ground bidirectional
rlabel metal5 s 0 135752 508088 136652 6 VGND
port 414 nsew ground bidirectional
rlabel metal5 s 0 126752 508088 127652 6 VGND
port 415 nsew ground bidirectional
rlabel metal5 s 0 117752 508088 118652 6 VGND
port 416 nsew ground bidirectional
rlabel metal5 s 0 108752 508088 109652 6 VGND
port 417 nsew ground bidirectional
rlabel metal5 s 0 99752 508088 100652 6 VGND
port 418 nsew ground bidirectional
rlabel metal5 s 0 90752 508088 91652 6 VGND
port 419 nsew ground bidirectional
rlabel metal5 s 0 81752 508088 82652 6 VGND
port 420 nsew ground bidirectional
rlabel metal5 s 0 72752 508088 73652 6 VGND
port 421 nsew ground bidirectional
rlabel metal5 s 0 63752 508088 64652 6 VGND
port 422 nsew ground bidirectional
rlabel metal5 s 0 54752 508088 55652 6 VGND
port 423 nsew ground bidirectional
rlabel metal5 s 0 45752 508088 46652 6 VGND
port 424 nsew ground bidirectional
rlabel metal5 s 0 36752 508088 37652 6 VGND
port 425 nsew ground bidirectional
rlabel metal5 s 0 27752 508088 28652 6 VGND
port 426 nsew ground bidirectional
rlabel metal5 s 0 12 508088 912 6 VGND
port 427 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 508088 579884
string LEFview TRUE
string GDS_FILE /project/openlane/fpga_core/runs/fpga_core/results/magic/fpga_core.gds
string GDS_END 37108538
string GDS_START 19917628
<< end >>

