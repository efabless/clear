magic
tech sky130A
magscale 1 2
timestamp 1680903011
<< viali >>
rect 6561 24361 6595 24395
rect 9137 24361 9171 24395
rect 11713 24361 11747 24395
rect 14289 24361 14323 24395
rect 25789 24361 25823 24395
rect 27169 24361 27203 24395
rect 32321 24361 32355 24395
rect 34161 24361 34195 24395
rect 37933 24361 37967 24395
rect 39313 24361 39347 24395
rect 44741 24361 44775 24395
rect 3985 24293 4019 24327
rect 29009 24293 29043 24327
rect 35909 24293 35943 24327
rect 37473 24293 37507 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 16865 24225 16899 24259
rect 18981 24225 19015 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25145 24225 25179 24259
rect 26341 24225 26375 24259
rect 27721 24225 27755 24259
rect 29745 24225 29779 24259
rect 30021 24225 30055 24259
rect 37013 24225 37047 24259
rect 40049 24225 40083 24259
rect 40325 24225 40359 24259
rect 2237 24157 2271 24191
rect 3893 24157 3927 24191
rect 4169 24157 4203 24191
rect 4629 24157 4663 24191
rect 6469 24157 6503 24191
rect 6745 24157 6779 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 15117 24157 15151 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22017 24157 22051 24191
rect 24041 24157 24075 24191
rect 25053 24157 25087 24191
rect 26249 24157 26283 24191
rect 27537 24157 27571 24191
rect 28549 24157 28583 24191
rect 29193 24157 29227 24191
rect 31493 24157 31527 24191
rect 32505 24157 32539 24191
rect 33333 24157 33367 24191
rect 34069 24157 34103 24191
rect 34989 24157 35023 24191
rect 36553 24157 36587 24191
rect 37657 24157 37691 24191
rect 38485 24157 38519 24191
rect 38669 24157 38703 24191
rect 39221 24157 39255 24191
rect 41429 24157 41463 24191
rect 42809 24157 42843 24191
rect 45201 24157 45235 24191
rect 45937 24157 45971 24191
rect 46673 24157 46707 24191
rect 47225 24157 47259 24191
rect 47777 24157 47811 24191
rect 48605 24157 48639 24191
rect 10977 24089 11011 24123
rect 17141 24089 17175 24123
rect 27629 24089 27663 24123
rect 30941 24089 30975 24123
rect 32781 24089 32815 24123
rect 35725 24089 35759 24123
rect 1593 24021 1627 24055
rect 1685 24021 1719 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 23857 24021 23891 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 26157 24021 26191 24055
rect 28365 24021 28399 24055
rect 31309 24021 31343 24055
rect 31861 24021 31895 24055
rect 33425 24021 33459 24055
rect 35081 24021 35115 24055
rect 36369 24021 36403 24055
rect 36829 24021 36863 24055
rect 42073 24021 42107 24055
rect 42625 24021 42659 24055
rect 45385 24021 45419 24055
rect 46121 24021 46155 24055
rect 46857 24021 46891 24055
rect 47961 24021 47995 24055
rect 49249 24021 49283 24055
rect 1777 23817 1811 23851
rect 12265 23817 12299 23851
rect 12357 23817 12391 23851
rect 24225 23817 24259 23851
rect 29377 23817 29411 23851
rect 30205 23817 30239 23851
rect 36093 23817 36127 23851
rect 38485 23817 38519 23851
rect 39037 23817 39071 23851
rect 39865 23817 39899 23851
rect 40325 23817 40359 23851
rect 42165 23817 42199 23851
rect 43269 23817 43303 23851
rect 45753 23817 45787 23851
rect 47593 23817 47627 23851
rect 47869 23817 47903 23851
rect 1593 23749 1627 23783
rect 3985 23749 4019 23783
rect 9137 23749 9171 23783
rect 10977 23749 11011 23783
rect 14289 23749 14323 23783
rect 16129 23749 16163 23783
rect 18981 23749 19015 23783
rect 21189 23749 21223 23783
rect 22293 23749 22327 23783
rect 30113 23749 30147 23783
rect 32321 23749 32355 23783
rect 32965 23749 32999 23783
rect 34161 23749 34195 23783
rect 34897 23749 34931 23783
rect 35633 23749 35667 23783
rect 38669 23749 38703 23783
rect 2145 23681 2179 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 7113 23681 7147 23715
rect 7205 23681 7239 23715
rect 7941 23681 7975 23715
rect 9873 23681 9907 23715
rect 13277 23681 13311 23715
rect 15117 23681 15151 23715
rect 16957 23681 16991 23715
rect 18705 23681 18739 23715
rect 21005 23681 21039 23715
rect 29561 23681 29595 23715
rect 31493 23681 31527 23715
rect 33425 23681 33459 23715
rect 33977 23681 34011 23715
rect 34713 23681 34747 23715
rect 35449 23681 35483 23715
rect 36277 23681 36311 23715
rect 36921 23681 36955 23715
rect 37289 23681 37323 23715
rect 37933 23681 37967 23715
rect 38209 23681 38243 23715
rect 40877 23681 40911 23715
rect 41521 23681 41555 23715
rect 41797 23681 41831 23715
rect 42625 23681 42659 23715
rect 43729 23681 43763 23715
rect 44465 23681 44499 23715
rect 45017 23681 45051 23715
rect 46765 23681 46799 23715
rect 47317 23681 47351 23715
rect 48053 23681 48087 23715
rect 48329 23681 48363 23715
rect 49065 23681 49099 23715
rect 5457 23613 5491 23647
rect 6469 23613 6503 23647
rect 7389 23613 7423 23647
rect 12541 23613 12575 23647
rect 17877 23613 17911 23647
rect 22017 23613 22051 23647
rect 24869 23613 24903 23647
rect 25145 23613 25179 23647
rect 27169 23613 27203 23647
rect 27445 23613 27479 23647
rect 6745 23545 6779 23579
rect 11897 23545 11931 23579
rect 30849 23545 30883 23579
rect 31033 23545 31067 23579
rect 31769 23545 31803 23579
rect 40693 23545 40727 23579
rect 49249 23545 49283 23579
rect 2237 23477 2271 23511
rect 6561 23477 6595 23511
rect 11529 23477 11563 23511
rect 20453 23477 20487 23511
rect 21649 23477 21683 23511
rect 23765 23477 23799 23511
rect 26617 23477 26651 23511
rect 28917 23477 28951 23511
rect 30573 23477 30607 23511
rect 31309 23477 31343 23511
rect 36737 23477 36771 23511
rect 37749 23477 37783 23511
rect 41337 23477 41371 23511
rect 43913 23477 43947 23511
rect 44649 23477 44683 23511
rect 46949 23477 46983 23511
rect 48513 23477 48547 23511
rect 3801 23273 3835 23307
rect 3985 23273 4019 23307
rect 14473 23273 14507 23307
rect 27524 23273 27558 23307
rect 29009 23273 29043 23307
rect 30002 23273 30036 23307
rect 31861 23273 31895 23307
rect 32505 23273 32539 23307
rect 33241 23273 33275 23307
rect 33977 23273 34011 23307
rect 34437 23273 34471 23307
rect 36829 23273 36863 23307
rect 37289 23273 37323 23307
rect 43637 23273 43671 23307
rect 13645 23205 13679 23239
rect 14933 23205 14967 23239
rect 18889 23205 18923 23239
rect 19441 23205 19475 23239
rect 37013 23205 37047 23239
rect 48421 23205 48455 23239
rect 3617 23137 3651 23171
rect 4721 23137 4755 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11529 23137 11563 23171
rect 13921 23137 13955 23171
rect 20085 23137 20119 23171
rect 22569 23137 22603 23171
rect 25145 23137 25179 23171
rect 26341 23137 26375 23171
rect 27261 23137 27295 23171
rect 29745 23137 29779 23171
rect 1777 23069 1811 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9321 23069 9355 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 19625 23069 19659 23103
rect 22293 23069 22327 23103
rect 25053 23069 25087 23103
rect 33885 23069 33919 23103
rect 35081 23069 35115 23103
rect 35725 23069 35759 23103
rect 41153 23069 41187 23103
rect 43913 23069 43947 23103
rect 48605 23069 48639 23103
rect 49065 23069 49099 23103
rect 2789 23001 2823 23035
rect 3433 23001 3467 23035
rect 4537 23001 4571 23035
rect 9597 23001 9631 23035
rect 11805 23001 11839 23035
rect 14381 23001 14415 23035
rect 16497 23001 16531 23035
rect 17417 23001 17451 23035
rect 20361 23001 20395 23035
rect 26249 23001 26283 23035
rect 32413 23001 32447 23035
rect 33149 23001 33183 23035
rect 36645 23001 36679 23035
rect 48145 23001 48179 23035
rect 4169 22933 4203 22967
rect 4629 22933 4663 22967
rect 9045 22933 9079 22967
rect 11069 22933 11103 22967
rect 13277 22933 13311 22967
rect 21833 22933 21867 22967
rect 24041 22933 24075 22967
rect 24593 22933 24627 22967
rect 24961 22933 24995 22967
rect 25789 22933 25823 22967
rect 26157 22933 26191 22967
rect 26801 22933 26835 22967
rect 29285 22933 29319 22967
rect 31493 22933 31527 22967
rect 31953 22933 31987 22967
rect 34897 22933 34931 22967
rect 35541 22933 35575 22967
rect 36185 22933 36219 22967
rect 42441 22933 42475 22967
rect 44557 22933 44591 22967
rect 49249 22933 49283 22967
rect 14565 22729 14599 22763
rect 21465 22729 21499 22763
rect 25789 22729 25823 22763
rect 27169 22729 27203 22763
rect 30573 22729 30607 22763
rect 33241 22729 33275 22763
rect 35081 22729 35115 22763
rect 48605 22729 48639 22763
rect 10701 22661 10735 22695
rect 12725 22661 12759 22695
rect 16129 22661 16163 22695
rect 17141 22661 17175 22695
rect 22477 22661 22511 22695
rect 27537 22661 27571 22695
rect 31585 22661 31619 22695
rect 31861 22661 31895 22695
rect 38117 22661 38151 22695
rect 39957 22661 39991 22695
rect 1777 22593 1811 22627
rect 3801 22593 3835 22627
rect 4813 22593 4847 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 7941 22593 7975 22627
rect 9965 22593 9999 22627
rect 11805 22593 11839 22627
rect 15117 22593 15151 22627
rect 19257 22593 19291 22627
rect 19717 22593 19751 22627
rect 23121 22593 23155 22627
rect 25697 22593 25731 22627
rect 28365 22593 28399 22627
rect 30941 22593 30975 22627
rect 31033 22593 31067 22627
rect 32413 22593 32447 22627
rect 32965 22593 32999 22627
rect 33609 22593 33643 22627
rect 33885 22593 33919 22627
rect 34989 22593 35023 22627
rect 37565 22593 37599 22627
rect 37841 22593 37875 22627
rect 48789 22593 48823 22627
rect 49065 22593 49099 22627
rect 2789 22525 2823 22559
rect 3893 22525 3927 22559
rect 4077 22525 4111 22559
rect 5089 22525 5123 22559
rect 7389 22525 7423 22559
rect 8677 22525 8711 22559
rect 12449 22525 12483 22559
rect 16865 22525 16899 22559
rect 19993 22525 20027 22559
rect 23397 22525 23431 22559
rect 25881 22525 25915 22559
rect 26433 22525 26467 22559
rect 27629 22525 27663 22559
rect 27721 22525 27755 22559
rect 31125 22525 31159 22559
rect 39589 22525 39623 22559
rect 18613 22457 18647 22491
rect 21925 22457 21959 22491
rect 33057 22457 33091 22491
rect 34713 22457 34747 22491
rect 3433 22389 3467 22423
rect 6469 22389 6503 22423
rect 6745 22389 6779 22423
rect 11897 22389 11931 22423
rect 14197 22389 14231 22423
rect 19073 22389 19107 22423
rect 22201 22389 22235 22423
rect 24869 22389 24903 22423
rect 25329 22389 25363 22423
rect 26525 22389 26559 22423
rect 26709 22389 26743 22423
rect 28628 22389 28662 22423
rect 30113 22389 30147 22423
rect 32505 22389 32539 22423
rect 35357 22389 35391 22423
rect 49249 22389 49283 22423
rect 27537 22185 27571 22219
rect 29561 22185 29595 22219
rect 29745 22185 29779 22219
rect 33885 22185 33919 22219
rect 29193 22117 29227 22151
rect 2053 22049 2087 22083
rect 3525 22049 3559 22083
rect 4445 22049 4479 22083
rect 7297 22049 7331 22083
rect 9965 22049 9999 22083
rect 11253 22049 11287 22083
rect 13369 22049 13403 22083
rect 15669 22049 15703 22083
rect 17141 22049 17175 22083
rect 20085 22049 20119 22083
rect 23949 22049 23983 22083
rect 25145 22049 25179 22083
rect 29285 22049 29319 22083
rect 30665 22049 30699 22083
rect 31861 22049 31895 22083
rect 34253 22049 34287 22083
rect 1777 21981 1811 22015
rect 4169 21981 4203 22015
rect 6285 21981 6319 22015
rect 6929 21981 6963 22015
rect 8769 21981 8803 22015
rect 9781 21981 9815 22015
rect 10517 21981 10551 22015
rect 12541 21981 12575 22015
rect 14565 21981 14599 22015
rect 15209 21981 15243 22015
rect 20361 21981 20395 22015
rect 21281 21981 21315 22015
rect 22293 21981 22327 22015
rect 23673 21981 23707 22015
rect 23765 21981 23799 22015
rect 25053 21981 25087 22015
rect 25789 21981 25823 22015
rect 28825 21981 28859 22015
rect 30481 21981 30515 22015
rect 32597 21981 32631 22015
rect 32873 21981 32907 22015
rect 34069 21981 34103 22015
rect 48789 21981 48823 22015
rect 49065 21981 49099 22015
rect 8585 21913 8619 21947
rect 14381 21913 14415 21947
rect 17417 21913 17451 21947
rect 19533 21913 19567 21947
rect 19717 21913 19751 21947
rect 22661 21913 22695 21947
rect 24961 21913 24995 21947
rect 26065 21913 26099 21947
rect 30573 21913 30607 21947
rect 31401 21913 31435 21947
rect 32229 21913 32263 21947
rect 3433 21845 3467 21879
rect 5825 21845 5859 21879
rect 6101 21845 6135 21879
rect 8953 21845 8987 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 14933 21845 14967 21879
rect 18889 21845 18923 21879
rect 22109 21845 22143 21879
rect 23305 21845 23339 21879
rect 24593 21845 24627 21879
rect 27997 21845 28031 21879
rect 28641 21845 28675 21879
rect 30113 21845 30147 21879
rect 31493 21845 31527 21879
rect 32045 21845 32079 21879
rect 33701 21845 33735 21879
rect 49249 21845 49283 21879
rect 9413 21641 9447 21675
rect 10241 21641 10275 21675
rect 10977 21641 11011 21675
rect 11161 21641 11195 21675
rect 16037 21641 16071 21675
rect 22017 21641 22051 21675
rect 23029 21641 23063 21675
rect 26709 21641 26743 21675
rect 27629 21641 27663 21675
rect 27721 21641 27755 21675
rect 31125 21641 31159 21675
rect 7941 21573 7975 21607
rect 15945 21573 15979 21607
rect 23673 21573 23707 21607
rect 33609 21573 33643 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 5641 21505 5675 21539
rect 7021 21505 7055 21539
rect 7665 21505 7699 21539
rect 12173 21505 12207 21539
rect 16865 21505 16899 21539
rect 21281 21505 21315 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 25973 21505 26007 21539
rect 26065 21505 26099 21539
rect 31033 21505 31067 21539
rect 31953 21505 31987 21539
rect 32413 21505 32447 21539
rect 32873 21505 32907 21539
rect 47961 21505 47995 21539
rect 2789 21437 2823 21471
rect 3893 21437 3927 21471
rect 5733 21437 5767 21471
rect 5825 21437 5859 21471
rect 10333 21437 10367 21471
rect 10517 21437 10551 21471
rect 12265 21437 12299 21471
rect 12357 21437 12391 21471
rect 13093 21437 13127 21471
rect 13369 21437 13403 21471
rect 16221 21437 16255 21471
rect 17325 21437 17359 21471
rect 18705 21437 18739 21471
rect 18981 21437 19015 21471
rect 22477 21437 22511 21471
rect 22661 21437 22695 21471
rect 25145 21437 25179 21471
rect 26249 21437 26283 21471
rect 27813 21437 27847 21471
rect 28457 21437 28491 21471
rect 28733 21437 28767 21471
rect 31217 21437 31251 21471
rect 33425 21437 33459 21471
rect 49157 21437 49191 21471
rect 6469 21369 6503 21403
rect 7205 21369 7239 21403
rect 15577 21369 15611 21403
rect 27261 21369 27295 21403
rect 33241 21369 33275 21403
rect 5273 21301 5307 21335
rect 6653 21301 6687 21335
rect 9689 21301 9723 21335
rect 9873 21301 9907 21335
rect 11345 21301 11379 21335
rect 11805 21301 11839 21335
rect 14841 21301 14875 21335
rect 15301 21301 15335 21335
rect 20453 21301 20487 21335
rect 20821 21301 20855 21335
rect 21005 21301 21039 21335
rect 25605 21301 25639 21335
rect 30205 21301 30239 21335
rect 30665 21301 30699 21335
rect 31769 21301 31803 21335
rect 32505 21301 32539 21335
rect 33057 21301 33091 21335
rect 47685 21301 47719 21335
rect 3433 21097 3467 21131
rect 15761 21097 15795 21131
rect 27813 21097 27847 21131
rect 32505 21097 32539 21131
rect 14289 21029 14323 21063
rect 14565 21029 14599 21063
rect 21833 21029 21867 21063
rect 4261 20961 4295 20995
rect 5733 20961 5767 20995
rect 8309 20961 8343 20995
rect 8493 20961 8527 20995
rect 9597 20961 9631 20995
rect 12633 20961 12667 20995
rect 15117 20961 15151 20995
rect 16405 20961 16439 20995
rect 17417 20961 17451 20995
rect 17601 20961 17635 20995
rect 18613 20961 18647 20995
rect 18705 20961 18739 20995
rect 19717 20961 19751 20995
rect 22661 20961 22695 20995
rect 23857 20961 23891 20995
rect 25329 20961 25363 20995
rect 26341 20961 26375 20995
rect 28549 20961 28583 20995
rect 30021 20961 30055 20995
rect 1777 20893 1811 20927
rect 3985 20893 4019 20927
rect 5457 20893 5491 20927
rect 9321 20893 9355 20927
rect 10977 20893 11011 20927
rect 11989 20893 12023 20927
rect 13737 20893 13771 20927
rect 19441 20893 19475 20927
rect 25697 20893 25731 20927
rect 26065 20893 26099 20927
rect 28273 20893 28307 20927
rect 29745 20893 29779 20927
rect 31125 20893 31159 20927
rect 32689 20893 32723 20927
rect 32965 20893 32999 20927
rect 2789 20825 2823 20859
rect 3617 20825 3651 20859
rect 7757 20825 7791 20859
rect 8217 20825 8251 20859
rect 11345 20825 11379 20859
rect 16221 20825 16255 20859
rect 23765 20825 23799 20859
rect 25053 20825 25087 20859
rect 31861 20825 31895 20859
rect 5181 20757 5215 20791
rect 7205 20757 7239 20791
rect 7573 20757 7607 20791
rect 7849 20757 7883 20791
rect 11437 20757 11471 20791
rect 13921 20757 13955 20791
rect 14933 20757 14967 20791
rect 15025 20757 15059 20791
rect 16129 20757 16163 20791
rect 16957 20757 16991 20791
rect 17325 20757 17359 20791
rect 18153 20757 18187 20791
rect 18521 20757 18555 20791
rect 21189 20757 21223 20791
rect 21649 20757 21683 20791
rect 22109 20757 22143 20791
rect 22477 20757 22511 20791
rect 22569 20757 22603 20791
rect 23305 20757 23339 20791
rect 23673 20757 23707 20791
rect 24685 20757 24719 20791
rect 25145 20757 25179 20791
rect 31217 20757 31251 20791
rect 31953 20757 31987 20791
rect 5641 20553 5675 20587
rect 12909 20553 12943 20587
rect 16129 20553 16163 20587
rect 17509 20553 17543 20587
rect 18153 20553 18187 20587
rect 18521 20553 18555 20587
rect 18889 20553 18923 20587
rect 23397 20553 23431 20587
rect 24041 20553 24075 20587
rect 26525 20553 26559 20587
rect 26801 20553 26835 20587
rect 27629 20553 27663 20587
rect 30941 20553 30975 20587
rect 31769 20553 31803 20587
rect 8769 20485 8803 20519
rect 16773 20485 16807 20519
rect 17417 20485 17451 20519
rect 22753 20485 22787 20519
rect 32137 20485 32171 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 5733 20417 5767 20451
rect 6561 20417 6595 20451
rect 11805 20417 11839 20451
rect 13001 20417 13035 20451
rect 13737 20417 13771 20451
rect 16037 20417 16071 20451
rect 19717 20417 19751 20451
rect 22017 20417 22051 20451
rect 24317 20417 24351 20451
rect 27537 20417 27571 20451
rect 28365 20417 28399 20451
rect 31033 20417 31067 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 5825 20349 5859 20383
rect 7297 20349 7331 20383
rect 9413 20349 9447 20383
rect 9689 20349 9723 20383
rect 13185 20349 13219 20383
rect 14013 20349 14047 20383
rect 16865 20349 16899 20383
rect 17693 20349 17727 20383
rect 18981 20349 19015 20383
rect 19073 20349 19107 20383
rect 19993 20349 20027 20383
rect 24593 20349 24627 20383
rect 26065 20349 26099 20383
rect 27721 20349 27755 20383
rect 28641 20349 28675 20383
rect 31125 20349 31159 20383
rect 8953 20281 8987 20315
rect 17049 20281 17083 20315
rect 27169 20281 27203 20315
rect 31585 20281 31619 20315
rect 5273 20213 5307 20247
rect 8401 20213 8435 20247
rect 11161 20213 11195 20247
rect 11897 20213 11931 20247
rect 12541 20213 12575 20247
rect 15485 20213 15519 20247
rect 21465 20213 21499 20247
rect 26433 20213 26467 20247
rect 30113 20213 30147 20247
rect 30573 20213 30607 20247
rect 11805 20009 11839 20043
rect 14197 20009 14231 20043
rect 17233 20009 17267 20043
rect 18705 20009 18739 20043
rect 19717 20009 19751 20043
rect 6285 19941 6319 19975
rect 16957 19941 16991 19975
rect 27629 19941 27663 19975
rect 29745 19941 29779 19975
rect 4537 19873 4571 19907
rect 6745 19873 6779 19907
rect 7021 19873 7055 19907
rect 9137 19873 9171 19907
rect 10885 19873 10919 19907
rect 12357 19873 12391 19907
rect 13645 19873 13679 19907
rect 14841 19873 14875 19907
rect 16773 19873 16807 19907
rect 17693 19873 17727 19907
rect 17877 19873 17911 19907
rect 20545 19873 20579 19907
rect 22017 19873 22051 19907
rect 23857 19873 23891 19907
rect 25329 19873 25363 19907
rect 28641 19873 28675 19907
rect 31309 19873 31343 19907
rect 1777 19805 1811 19839
rect 12265 19805 12299 19839
rect 14565 19805 14599 19839
rect 18889 19805 18923 19839
rect 20269 19805 20303 19839
rect 22569 19805 22603 19839
rect 23765 19805 23799 19839
rect 25881 19805 25915 19839
rect 28365 19805 28399 19839
rect 29929 19805 29963 19839
rect 30205 19805 30239 19839
rect 31125 19805 31159 19839
rect 2789 19737 2823 19771
rect 3617 19737 3651 19771
rect 4813 19737 4847 19771
rect 9413 19737 9447 19771
rect 11345 19737 11379 19771
rect 11529 19737 11563 19771
rect 13461 19737 13495 19771
rect 19625 19737 19659 19771
rect 22753 19737 22787 19771
rect 25053 19737 25087 19771
rect 26157 19737 26191 19771
rect 3433 19669 3467 19703
rect 3893 19669 3927 19703
rect 4077 19669 4111 19703
rect 4261 19669 4295 19703
rect 8493 19669 8527 19703
rect 12173 19669 12207 19703
rect 13001 19669 13035 19703
rect 13369 19669 13403 19703
rect 16313 19669 16347 19703
rect 17601 19669 17635 19703
rect 18429 19669 18463 19703
rect 23305 19669 23339 19703
rect 23673 19669 23707 19703
rect 24685 19669 24719 19703
rect 25145 19669 25179 19703
rect 27997 19669 28031 19703
rect 30389 19669 30423 19703
rect 30757 19669 30791 19703
rect 31217 19669 31251 19703
rect 5273 19465 5307 19499
rect 5733 19465 5767 19499
rect 10885 19465 10919 19499
rect 14381 19465 14415 19499
rect 14841 19465 14875 19499
rect 17877 19465 17911 19499
rect 18337 19465 18371 19499
rect 19073 19465 19107 19499
rect 21465 19465 21499 19499
rect 22385 19465 22419 19499
rect 26433 19465 26467 19499
rect 27261 19465 27295 19499
rect 27721 19465 27755 19499
rect 30481 19465 30515 19499
rect 4353 19397 4387 19431
rect 5641 19397 5675 19431
rect 9321 19397 9355 19431
rect 13921 19397 13955 19431
rect 16773 19397 16807 19431
rect 22477 19397 22511 19431
rect 28549 19397 28583 19431
rect 1777 19329 1811 19363
rect 2789 19329 2823 19363
rect 3617 19329 3651 19363
rect 6653 19329 6687 19363
rect 7481 19329 7515 19363
rect 8585 19329 8619 19363
rect 10793 19329 10827 19363
rect 11713 19329 11747 19363
rect 14749 19329 14783 19363
rect 15669 19329 15703 19363
rect 17425 19329 17459 19363
rect 17785 19329 17819 19363
rect 18245 19329 18279 19363
rect 19257 19329 19291 19363
rect 24041 19329 24075 19363
rect 24133 19329 24167 19363
rect 24961 19329 24995 19363
rect 30665 19329 30699 19363
rect 31125 19329 31159 19363
rect 5825 19261 5859 19295
rect 10149 19261 10183 19295
rect 10977 19261 11011 19295
rect 11989 19261 12023 19295
rect 14933 19261 14967 19295
rect 16957 19261 16991 19295
rect 18429 19261 18463 19295
rect 19717 19261 19751 19295
rect 19993 19261 20027 19295
rect 22569 19261 22603 19295
rect 23029 19261 23063 19295
rect 24317 19261 24351 19295
rect 25789 19261 25823 19295
rect 26985 19261 27019 19295
rect 27445 19261 27479 19295
rect 28273 19261 28307 19295
rect 31033 19261 31067 19295
rect 10425 19193 10459 19227
rect 17233 19193 17267 19227
rect 22017 19193 22051 19227
rect 23397 19193 23431 19227
rect 10333 19125 10367 19159
rect 13461 19125 13495 19159
rect 14013 19125 14047 19159
rect 15761 19125 15795 19159
rect 16221 19125 16255 19159
rect 16497 19125 16531 19159
rect 23673 19125 23707 19159
rect 27905 19125 27939 19159
rect 30021 19125 30055 19159
rect 3893 18921 3927 18955
rect 22937 18921 22971 18955
rect 8585 18853 8619 18887
rect 11621 18853 11655 18887
rect 14749 18853 14783 18887
rect 18153 18853 18187 18887
rect 20913 18853 20947 18887
rect 30849 18853 30883 18887
rect 2053 18785 2087 18819
rect 3985 18785 4019 18819
rect 6837 18785 6871 18819
rect 9965 18785 9999 18819
rect 12173 18785 12207 18819
rect 13553 18785 13587 18819
rect 15209 18785 15243 18819
rect 17509 18785 17543 18819
rect 18705 18785 18739 18819
rect 20361 18785 20395 18819
rect 21189 18785 21223 18819
rect 21465 18785 21499 18819
rect 24593 18785 24627 18819
rect 25421 18785 25455 18819
rect 27169 18785 27203 18819
rect 30205 18785 30239 18819
rect 30297 18785 30331 18819
rect 1777 18717 1811 18751
rect 4629 18717 4663 18751
rect 9781 18717 9815 18751
rect 9873 18717 9907 18751
rect 10609 18717 10643 18751
rect 18521 18717 18555 18751
rect 19625 18717 19659 18751
rect 23581 18717 23615 18751
rect 27629 18717 27663 18751
rect 27905 18717 27939 18751
rect 4905 18649 4939 18683
rect 7113 18649 7147 18683
rect 10977 18649 11011 18683
rect 12081 18649 12115 18683
rect 12817 18649 12851 18683
rect 14565 18649 14599 18683
rect 15485 18649 15519 18683
rect 24041 18649 24075 18683
rect 25697 18649 25731 18683
rect 3341 18581 3375 18615
rect 3525 18581 3559 18615
rect 6377 18581 6411 18615
rect 9045 18581 9079 18615
rect 9413 18581 9447 18615
rect 11069 18581 11103 18615
rect 11989 18581 12023 18615
rect 14197 18581 14231 18615
rect 16957 18581 16991 18615
rect 18061 18581 18095 18615
rect 18613 18581 18647 18615
rect 19349 18581 19383 18615
rect 23397 18581 23431 18615
rect 24133 18581 24167 18615
rect 25053 18581 25087 18615
rect 29745 18581 29779 18615
rect 30113 18581 30147 18615
rect 10425 18377 10459 18411
rect 15025 18377 15059 18411
rect 16865 18377 16899 18411
rect 22569 18377 22603 18411
rect 22845 18377 22879 18411
rect 24869 18377 24903 18411
rect 26801 18377 26835 18411
rect 27169 18377 27203 18411
rect 30757 18377 30791 18411
rect 31493 18377 31527 18411
rect 9965 18309 9999 18343
rect 14381 18309 14415 18343
rect 15393 18309 15427 18343
rect 15485 18309 15519 18343
rect 18153 18309 18187 18343
rect 22017 18309 22051 18343
rect 26065 18309 26099 18343
rect 28365 18309 28399 18343
rect 30665 18309 30699 18343
rect 31309 18309 31343 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 5641 18241 5675 18275
rect 5733 18241 5767 18275
rect 6745 18241 6779 18275
rect 8493 18241 8527 18275
rect 10793 18241 10827 18275
rect 12357 18241 12391 18275
rect 13645 18241 13679 18275
rect 16221 18241 16255 18275
rect 17233 18241 17267 18275
rect 19901 18241 19935 18275
rect 21097 18241 21131 18275
rect 25329 18241 25363 18275
rect 26525 18241 26559 18275
rect 28089 18241 28123 18275
rect 2053 18173 2087 18207
rect 3893 18173 3927 18207
rect 5917 18173 5951 18207
rect 7205 18173 7239 18207
rect 9229 18173 9263 18207
rect 10885 18173 10919 18207
rect 11069 18173 11103 18207
rect 12449 18173 12483 18207
rect 12633 18173 12667 18207
rect 13185 18173 13219 18207
rect 15669 18173 15703 18207
rect 17325 18173 17359 18207
rect 17417 18173 17451 18207
rect 18889 18173 18923 18207
rect 19993 18173 20027 18207
rect 20177 18173 20211 18207
rect 21189 18173 21223 18207
rect 21281 18173 21315 18207
rect 23121 18173 23155 18207
rect 23397 18173 23431 18207
rect 30849 18173 30883 18207
rect 11989 18105 12023 18139
rect 20729 18105 20763 18139
rect 30297 18105 30331 18139
rect 5273 18037 5307 18071
rect 9689 18037 9723 18071
rect 10057 18037 10091 18071
rect 11713 18037 11747 18071
rect 13277 18037 13311 18071
rect 16037 18037 16071 18071
rect 16497 18037 16531 18071
rect 18245 18037 18279 18071
rect 19533 18037 19567 18071
rect 29837 18037 29871 18071
rect 3433 17833 3467 17867
rect 3617 17833 3651 17867
rect 10609 17833 10643 17867
rect 13737 17833 13771 17867
rect 20729 17833 20763 17867
rect 30941 17833 30975 17867
rect 4445 17765 4479 17799
rect 6653 17765 6687 17799
rect 7849 17765 7883 17799
rect 18337 17765 18371 17799
rect 22017 17765 22051 17799
rect 26617 17765 26651 17799
rect 29745 17765 29779 17799
rect 7389 17697 7423 17731
rect 8493 17697 8527 17731
rect 9873 17697 9907 17731
rect 11161 17697 11195 17731
rect 11621 17697 11655 17731
rect 12265 17697 12299 17731
rect 14565 17697 14599 17731
rect 16313 17697 16347 17731
rect 16589 17697 16623 17731
rect 19441 17697 19475 17731
rect 21189 17697 21223 17731
rect 21281 17697 21315 17731
rect 24869 17697 24903 17731
rect 27077 17697 27111 17731
rect 29193 17697 29227 17731
rect 30297 17697 30331 17731
rect 31493 17697 31527 17731
rect 1777 17629 1811 17663
rect 4905 17629 4939 17663
rect 7205 17629 7239 17663
rect 8217 17629 8251 17663
rect 9137 17629 9171 17663
rect 10977 17629 11011 17663
rect 11989 17629 12023 17663
rect 14381 17629 14415 17663
rect 19717 17629 19751 17663
rect 22293 17629 22327 17663
rect 31309 17629 31343 17663
rect 31401 17629 31435 17663
rect 2513 17561 2547 17595
rect 4261 17561 4295 17595
rect 5181 17561 5215 17595
rect 8309 17561 8343 17595
rect 11069 17561 11103 17595
rect 21097 17561 21131 17595
rect 22569 17561 22603 17595
rect 25145 17561 25179 17595
rect 27353 17561 27387 17595
rect 30113 17561 30147 17595
rect 3801 17493 3835 17527
rect 14841 17493 14875 17527
rect 15117 17493 15151 17527
rect 15393 17493 15427 17527
rect 16037 17493 16071 17527
rect 18061 17493 18095 17527
rect 18705 17493 18739 17527
rect 21833 17493 21867 17527
rect 24041 17493 24075 17527
rect 24409 17493 24443 17527
rect 28825 17493 28859 17527
rect 30205 17493 30239 17527
rect 5273 17289 5307 17323
rect 7297 17289 7331 17323
rect 8033 17289 8067 17323
rect 9965 17289 9999 17323
rect 12541 17289 12575 17323
rect 13737 17289 13771 17323
rect 16865 17289 16899 17323
rect 22017 17289 22051 17323
rect 24317 17289 24351 17323
rect 29837 17289 29871 17323
rect 30573 17289 30607 17323
rect 30941 17289 30975 17323
rect 4629 17221 4663 17255
rect 8401 17221 8435 17255
rect 10977 17221 11011 17255
rect 11805 17221 11839 17255
rect 13001 17221 13035 17255
rect 18429 17221 18463 17255
rect 20177 17221 20211 17255
rect 22477 17221 22511 17255
rect 24961 17221 24995 17255
rect 26801 17221 26835 17255
rect 30849 17221 30883 17255
rect 1777 17153 1811 17187
rect 3617 17153 3651 17187
rect 5641 17153 5675 17187
rect 7205 17153 7239 17187
rect 9873 17153 9907 17187
rect 10793 17153 10827 17187
rect 12909 17153 12943 17187
rect 14105 17153 14139 17187
rect 14749 17153 14783 17187
rect 14933 17153 14967 17187
rect 15209 17153 15243 17187
rect 15669 17153 15703 17187
rect 16313 17153 16347 17187
rect 17233 17153 17267 17187
rect 21097 17153 21131 17187
rect 22385 17153 22419 17187
rect 23673 17153 23707 17187
rect 24685 17153 24719 17187
rect 27813 17153 27847 17187
rect 2053 17085 2087 17119
rect 4997 17085 5031 17119
rect 5181 17085 5215 17119
rect 5733 17085 5767 17119
rect 5825 17085 5859 17119
rect 7481 17085 7515 17119
rect 8493 17085 8527 17119
rect 8677 17085 8711 17119
rect 10149 17085 10183 17119
rect 13185 17085 13219 17119
rect 14197 17085 14231 17119
rect 14381 17085 14415 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 18153 17085 18187 17119
rect 21189 17085 21223 17119
rect 21373 17085 21407 17119
rect 22569 17085 22603 17119
rect 23765 17085 23799 17119
rect 23857 17085 23891 17119
rect 26433 17085 26467 17119
rect 27169 17085 27203 17119
rect 28089 17085 28123 17119
rect 6837 17017 6871 17051
rect 11989 17017 12023 17051
rect 16129 17017 16163 17051
rect 6469 16949 6503 16983
rect 9137 16949 9171 16983
rect 9505 16949 9539 16983
rect 11345 16949 11379 16983
rect 15485 16949 15519 16983
rect 19901 16949 19935 16983
rect 20361 16949 20395 16983
rect 20729 16949 20763 16983
rect 23305 16949 23339 16983
rect 29561 16949 29595 16983
rect 3617 16745 3651 16779
rect 6009 16745 6043 16779
rect 7849 16745 7883 16779
rect 9781 16745 9815 16779
rect 12541 16745 12575 16779
rect 14381 16677 14415 16711
rect 15025 16677 15059 16711
rect 25697 16677 25731 16711
rect 3433 16609 3467 16643
rect 7113 16609 7147 16643
rect 7297 16609 7331 16643
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 10517 16609 10551 16643
rect 10701 16609 10735 16643
rect 11713 16609 11747 16643
rect 11897 16609 11931 16643
rect 12725 16609 12759 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 15485 16609 15519 16643
rect 15669 16609 15703 16643
rect 16405 16609 16439 16643
rect 16773 16609 16807 16643
rect 18705 16609 18739 16643
rect 19717 16609 19751 16643
rect 22477 16609 22511 16643
rect 22661 16609 22695 16643
rect 23765 16609 23799 16643
rect 25145 16609 25179 16643
rect 25329 16609 25363 16643
rect 25881 16609 25915 16643
rect 27077 16609 27111 16643
rect 27261 16609 27295 16643
rect 28273 16609 28307 16643
rect 28457 16609 28491 16643
rect 1777 16541 1811 16575
rect 4077 16541 4111 16575
rect 4905 16541 4939 16575
rect 9413 16541 9447 16575
rect 10425 16541 10459 16575
rect 14565 16541 14599 16575
rect 15393 16541 15427 16575
rect 17601 16541 17635 16575
rect 18245 16541 18279 16575
rect 19441 16541 19475 16575
rect 22385 16541 22419 16575
rect 23581 16541 23615 16575
rect 28181 16541 28215 16575
rect 2513 16473 2547 16507
rect 5917 16473 5951 16507
rect 9229 16473 9263 16507
rect 11621 16473 11655 16507
rect 21465 16473 21499 16507
rect 26985 16473 27019 16507
rect 6653 16405 6687 16439
rect 7021 16405 7055 16439
rect 8217 16405 8251 16439
rect 10057 16405 10091 16439
rect 11253 16405 11287 16439
rect 12265 16405 12299 16439
rect 13001 16405 13035 16439
rect 13369 16405 13403 16439
rect 16129 16405 16163 16439
rect 16313 16405 16347 16439
rect 17417 16405 17451 16439
rect 18061 16405 18095 16439
rect 22017 16405 22051 16439
rect 23213 16405 23247 16439
rect 23673 16405 23707 16439
rect 24685 16405 24719 16439
rect 25053 16405 25087 16439
rect 26617 16405 26651 16439
rect 27813 16405 27847 16439
rect 5733 16201 5767 16235
rect 7297 16201 7331 16235
rect 13737 16201 13771 16235
rect 16773 16201 16807 16235
rect 17141 16201 17175 16235
rect 17417 16201 17451 16235
rect 17877 16201 17911 16235
rect 20453 16201 20487 16235
rect 26617 16201 26651 16235
rect 27721 16201 27755 16235
rect 4353 16133 4387 16167
rect 7757 16133 7791 16167
rect 14657 16133 14691 16167
rect 19717 16133 19751 16167
rect 20545 16133 20579 16167
rect 1777 16065 1811 16099
rect 3525 16065 3559 16099
rect 5641 16065 5675 16099
rect 7665 16065 7699 16099
rect 8493 16065 8527 16099
rect 10609 16065 10643 16099
rect 11161 16065 11195 16099
rect 11989 16065 12023 16099
rect 14749 16065 14783 16099
rect 16313 16065 16347 16099
rect 17785 16065 17819 16099
rect 18613 16065 18647 16099
rect 21465 16065 21499 16099
rect 22293 16065 22327 16099
rect 23673 16065 23707 16099
rect 24317 16065 24351 16099
rect 24593 16065 24627 16099
rect 24869 16065 24903 16099
rect 26985 16065 27019 16099
rect 2053 15997 2087 16031
rect 5917 15997 5951 16031
rect 6653 15997 6687 16031
rect 7941 15997 7975 16031
rect 8769 15997 8803 16031
rect 10241 15997 10275 16031
rect 11713 15997 11747 16031
rect 12265 15997 12299 16031
rect 14841 15997 14875 16031
rect 15485 15997 15519 16031
rect 17969 15997 18003 16031
rect 18889 15997 18923 16031
rect 20637 15997 20671 16031
rect 22017 15997 22051 16031
rect 23765 15997 23799 16031
rect 23949 15997 23983 16031
rect 25145 15997 25179 16031
rect 10977 15929 11011 15963
rect 14289 15929 14323 15963
rect 20085 15929 20119 15963
rect 5273 15861 5307 15895
rect 16129 15861 16163 15895
rect 16957 15861 16991 15895
rect 21281 15861 21315 15895
rect 23305 15861 23339 15895
rect 7849 15657 7883 15691
rect 9321 15657 9355 15691
rect 9781 15657 9815 15691
rect 15853 15657 15887 15691
rect 22477 15657 22511 15691
rect 24501 15657 24535 15691
rect 3433 15589 3467 15623
rect 12081 15589 12115 15623
rect 13553 15589 13587 15623
rect 14473 15589 14507 15623
rect 19901 15589 19935 15623
rect 26341 15589 26375 15623
rect 2053 15521 2087 15555
rect 4445 15521 4479 15555
rect 4629 15521 4663 15555
rect 5641 15521 5675 15555
rect 5733 15521 5767 15555
rect 6929 15521 6963 15555
rect 8309 15521 8343 15555
rect 8401 15521 8435 15555
rect 10241 15521 10275 15555
rect 11437 15521 11471 15555
rect 12725 15521 12759 15555
rect 15025 15521 15059 15555
rect 16497 15521 16531 15555
rect 20269 15521 20303 15555
rect 22753 15521 22787 15555
rect 25789 15521 25823 15555
rect 1777 15453 1811 15487
rect 3617 15453 3651 15487
rect 6837 15453 6871 15487
rect 7481 15453 7515 15487
rect 12449 15453 12483 15487
rect 13277 15453 13311 15487
rect 13737 15453 13771 15487
rect 14841 15453 14875 15487
rect 17049 15453 17083 15487
rect 19625 15453 19659 15487
rect 23121 15453 23155 15487
rect 25605 15453 25639 15487
rect 5549 15385 5583 15419
rect 6745 15385 6779 15419
rect 9229 15385 9263 15419
rect 11345 15385 11379 15419
rect 14933 15385 14967 15419
rect 17325 15385 17359 15419
rect 20545 15385 20579 15419
rect 23949 15385 23983 15419
rect 25697 15385 25731 15419
rect 26433 15385 26467 15419
rect 3985 15317 4019 15351
rect 4353 15317 4387 15351
rect 5181 15317 5215 15351
rect 6377 15317 6411 15351
rect 8217 15317 8251 15351
rect 9873 15317 9907 15351
rect 10885 15317 10919 15351
rect 11253 15317 11287 15351
rect 12541 15317 12575 15351
rect 14105 15317 14139 15351
rect 15485 15317 15519 15351
rect 16221 15317 16255 15351
rect 16313 15317 16347 15351
rect 18797 15317 18831 15351
rect 19441 15317 19475 15351
rect 22017 15317 22051 15351
rect 22385 15317 22419 15351
rect 25237 15317 25271 15351
rect 3525 15113 3559 15147
rect 8677 15113 8711 15147
rect 9229 15113 9263 15147
rect 13001 15113 13035 15147
rect 23765 15113 23799 15147
rect 24041 15113 24075 15147
rect 24225 15113 24259 15147
rect 27077 15113 27111 15147
rect 7665 15045 7699 15079
rect 9689 15045 9723 15079
rect 10793 15045 10827 15079
rect 10885 15045 10919 15079
rect 14197 15045 14231 15079
rect 20177 15045 20211 15079
rect 22293 15045 22327 15079
rect 25145 15045 25179 15079
rect 1777 14977 1811 15011
rect 3709 14977 3743 15011
rect 4169 14977 4203 15011
rect 6653 14977 6687 15011
rect 8585 14977 8619 15011
rect 9597 14977 9631 15011
rect 11989 14977 12023 15011
rect 13369 14977 13403 15011
rect 17141 14977 17175 15011
rect 18889 14977 18923 15011
rect 20085 14977 20119 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 22017 14977 22051 15011
rect 24869 14977 24903 15011
rect 2053 14909 2087 14943
rect 4445 14909 4479 14943
rect 7757 14909 7791 14943
rect 7849 14909 7883 14943
rect 9873 14909 9907 14943
rect 10977 14909 11011 14943
rect 11713 14909 11747 14943
rect 13461 14909 13495 14943
rect 13645 14909 13679 14943
rect 14565 14909 14599 14943
rect 14841 14909 14875 14943
rect 16773 14909 16807 14943
rect 20361 14909 20395 14943
rect 6837 14841 6871 14875
rect 14013 14841 14047 14875
rect 5917 14773 5951 14807
rect 7297 14773 7331 14807
rect 10425 14773 10459 14807
rect 16313 14773 16347 14807
rect 19165 14773 19199 14807
rect 19349 14773 19383 14807
rect 19717 14773 19751 14807
rect 26617 14773 26651 14807
rect 3985 14569 4019 14603
rect 9413 14569 9447 14603
rect 11621 14569 11655 14603
rect 13737 14569 13771 14603
rect 14381 14569 14415 14603
rect 18613 14569 18647 14603
rect 19441 14569 19475 14603
rect 26985 14569 27019 14603
rect 7205 14501 7239 14535
rect 21557 14501 21591 14535
rect 21741 14501 21775 14535
rect 24041 14501 24075 14535
rect 2053 14433 2087 14467
rect 4905 14433 4939 14467
rect 8493 14433 8527 14467
rect 9873 14433 9907 14467
rect 10057 14433 10091 14467
rect 11161 14433 11195 14467
rect 12265 14433 12299 14467
rect 14933 14433 14967 14467
rect 16865 14433 16899 14467
rect 18889 14433 18923 14467
rect 21097 14433 21131 14467
rect 22293 14433 22327 14467
rect 25053 14433 25087 14467
rect 25145 14433 25179 14467
rect 26341 14433 26375 14467
rect 1777 14365 1811 14399
rect 5457 14365 5491 14399
rect 8217 14365 8251 14399
rect 10977 14365 11011 14399
rect 11989 14365 12023 14399
rect 14657 14365 14691 14399
rect 19625 14365 19659 14399
rect 21005 14365 21039 14399
rect 26157 14365 26191 14399
rect 4629 14297 4663 14331
rect 5733 14297 5767 14331
rect 8309 14297 8343 14331
rect 17141 14297 17175 14331
rect 22569 14297 22603 14331
rect 24961 14297 24995 14331
rect 26249 14297 26283 14331
rect 26801 14297 26835 14331
rect 3433 14229 3467 14263
rect 3525 14229 3559 14263
rect 4261 14229 4295 14263
rect 4721 14229 4755 14263
rect 7849 14229 7883 14263
rect 9045 14229 9079 14263
rect 9781 14229 9815 14263
rect 10609 14229 10643 14263
rect 11069 14229 11103 14263
rect 14105 14229 14139 14263
rect 16405 14229 16439 14263
rect 20545 14229 20579 14263
rect 20913 14229 20947 14263
rect 24593 14229 24627 14263
rect 25789 14229 25823 14263
rect 3433 14025 3467 14059
rect 4077 14025 4111 14059
rect 5641 14025 5675 14059
rect 6929 14025 6963 14059
rect 7297 14025 7331 14059
rect 8125 14025 8159 14059
rect 11989 14025 12023 14059
rect 13645 14025 13679 14059
rect 14749 14025 14783 14059
rect 14841 14025 14875 14059
rect 15577 14025 15611 14059
rect 18889 14025 18923 14059
rect 19441 14025 19475 14059
rect 23397 14025 23431 14059
rect 24961 14025 24995 14059
rect 25881 14025 25915 14059
rect 4537 13957 4571 13991
rect 5733 13957 5767 13991
rect 8493 13957 8527 13991
rect 8585 13957 8619 13991
rect 16681 13957 16715 13991
rect 21833 13957 21867 13991
rect 23765 13957 23799 13991
rect 23857 13957 23891 13991
rect 25053 13957 25087 13991
rect 25605 13957 25639 13991
rect 1777 13889 1811 13923
rect 3617 13889 3651 13923
rect 4445 13889 4479 13923
rect 7389 13889 7423 13923
rect 11621 13889 11655 13923
rect 12357 13889 12391 13923
rect 13553 13889 13587 13923
rect 15945 13889 15979 13923
rect 16037 13889 16071 13923
rect 19625 13889 19659 13923
rect 20453 13889 20487 13923
rect 20545 13889 20579 13923
rect 22569 13889 22603 13923
rect 25973 13889 26007 13923
rect 2053 13821 2087 13855
rect 4629 13821 4663 13855
rect 5825 13821 5859 13855
rect 6377 13821 6411 13855
rect 7481 13821 7515 13855
rect 8677 13821 8711 13855
rect 9321 13821 9355 13855
rect 9597 13821 9631 13855
rect 11069 13821 11103 13855
rect 12449 13821 12483 13855
rect 12541 13821 12575 13855
rect 13829 13821 13863 13855
rect 14933 13821 14967 13855
rect 16129 13821 16163 13855
rect 17141 13821 17175 13855
rect 20637 13821 20671 13855
rect 22661 13821 22695 13855
rect 22845 13821 22879 13855
rect 24041 13821 24075 13855
rect 25237 13821 25271 13855
rect 26157 13821 26191 13855
rect 6561 13753 6595 13787
rect 13185 13753 13219 13787
rect 14381 13753 14415 13787
rect 20085 13753 20119 13787
rect 22201 13753 22235 13787
rect 5273 13685 5307 13719
rect 17404 13685 17438 13719
rect 24593 13685 24627 13719
rect 4432 13481 4466 13515
rect 11437 13481 11471 13515
rect 13737 13481 13771 13515
rect 17398 13481 17432 13515
rect 18889 13481 18923 13515
rect 22109 13481 22143 13515
rect 22477 13481 22511 13515
rect 23949 13481 23983 13515
rect 22845 13413 22879 13447
rect 24133 13413 24167 13447
rect 2053 13345 2087 13379
rect 4169 13345 4203 13379
rect 6745 13345 6779 13379
rect 10977 13345 11011 13379
rect 11621 13345 11655 13379
rect 11989 13345 12023 13379
rect 14565 13345 14599 13379
rect 16497 13345 16531 13379
rect 17141 13345 17175 13379
rect 20361 13345 20395 13379
rect 23305 13345 23339 13379
rect 23489 13345 23523 13379
rect 1777 13277 1811 13311
rect 3893 13277 3927 13311
rect 9137 13277 9171 13311
rect 9413 13277 9447 13311
rect 10793 13277 10827 13311
rect 14289 13277 14323 13311
rect 19349 13277 19383 13311
rect 19441 13277 19475 13311
rect 3525 13209 3559 13243
rect 7021 13209 7055 13243
rect 12265 13209 12299 13243
rect 20637 13209 20671 13243
rect 23213 13209 23247 13243
rect 24593 13209 24627 13243
rect 25421 13209 25455 13243
rect 3341 13141 3375 13175
rect 5917 13141 5951 13175
rect 6285 13141 6319 13175
rect 6469 13141 6503 13175
rect 8493 13141 8527 13175
rect 10425 13141 10459 13175
rect 10885 13141 10919 13175
rect 16037 13141 16071 13175
rect 3617 12937 3651 12971
rect 5733 12937 5767 12971
rect 7297 12937 7331 12971
rect 12541 12937 12575 12971
rect 13737 12937 13771 12971
rect 14197 12937 14231 12971
rect 16221 12937 16255 12971
rect 17785 12937 17819 12971
rect 18153 12937 18187 12971
rect 21097 12937 21131 12971
rect 22201 12937 22235 12971
rect 24777 12937 24811 12971
rect 3525 12869 3559 12903
rect 4261 12869 4295 12903
rect 4445 12869 4479 12903
rect 4813 12869 4847 12903
rect 5641 12869 5675 12903
rect 6469 12869 6503 12903
rect 7205 12869 7239 12903
rect 11897 12869 11931 12903
rect 15669 12869 15703 12903
rect 18981 12869 19015 12903
rect 1869 12801 1903 12835
rect 10701 12801 10735 12835
rect 12909 12801 12943 12835
rect 14105 12801 14139 12835
rect 14933 12801 14967 12835
rect 16313 12801 16347 12835
rect 18245 12801 18279 12835
rect 21189 12801 21223 12835
rect 23029 12801 23063 12835
rect 1593 12733 1627 12767
rect 2789 12733 2823 12767
rect 4905 12733 4939 12767
rect 5917 12733 5951 12767
rect 7389 12733 7423 12767
rect 8033 12733 8067 12767
rect 8309 12733 8343 12767
rect 10057 12733 10091 12767
rect 13001 12733 13035 12767
rect 13185 12733 13219 12767
rect 14381 12733 14415 12767
rect 16865 12733 16899 12767
rect 18429 12733 18463 12767
rect 19809 12733 19843 12767
rect 21373 12733 21407 12767
rect 23305 12733 23339 12767
rect 25053 12733 25087 12767
rect 3157 12665 3191 12699
rect 10517 12665 10551 12699
rect 11345 12665 11379 12699
rect 2973 12597 3007 12631
rect 5273 12597 5307 12631
rect 6837 12597 6871 12631
rect 11161 12597 11195 12631
rect 11621 12597 11655 12631
rect 20729 12597 20763 12631
rect 3985 12393 4019 12427
rect 4629 12393 4663 12427
rect 7849 12393 7883 12427
rect 11805 12393 11839 12427
rect 14473 12393 14507 12427
rect 18061 12393 18095 12427
rect 18429 12393 18463 12427
rect 18981 12393 19015 12427
rect 21833 12393 21867 12427
rect 24501 12393 24535 12427
rect 3617 12325 3651 12359
rect 13001 12325 13035 12359
rect 18889 12325 18923 12359
rect 1869 12257 1903 12291
rect 4721 12257 4755 12291
rect 5365 12257 5399 12291
rect 7389 12257 7423 12291
rect 8401 12257 8435 12291
rect 9873 12257 9907 12291
rect 11253 12257 11287 12291
rect 12357 12257 12391 12291
rect 13645 12257 13679 12291
rect 15945 12257 15979 12291
rect 16589 12257 16623 12291
rect 19533 12257 19567 12291
rect 20085 12257 20119 12291
rect 22569 12257 22603 12291
rect 1593 12189 1627 12223
rect 4169 12189 4203 12223
rect 8309 12189 8343 12223
rect 11069 12189 11103 12223
rect 13369 12189 13403 12223
rect 14749 12189 14783 12223
rect 15577 12189 15611 12223
rect 16313 12189 16347 12223
rect 22293 12189 22327 12223
rect 2973 12121 3007 12155
rect 3157 12121 3191 12155
rect 5641 12121 5675 12155
rect 9137 12121 9171 12155
rect 10977 12121 11011 12155
rect 12265 12121 12299 12155
rect 13461 12121 13495 12155
rect 20361 12121 20395 12155
rect 8217 12053 8251 12087
rect 10609 12053 10643 12087
rect 12173 12053 12207 12087
rect 14105 12053 14139 12087
rect 18521 12053 18555 12087
rect 19349 12053 19383 12087
rect 24041 12053 24075 12087
rect 1777 11849 1811 11883
rect 3433 11849 3467 11883
rect 4445 11849 4479 11883
rect 5273 11849 5307 11883
rect 5641 11849 5675 11883
rect 6469 11849 6503 11883
rect 6745 11849 6779 11883
rect 12357 11849 12391 11883
rect 17325 11849 17359 11883
rect 18521 11849 18555 11883
rect 19165 11849 19199 11883
rect 1685 11781 1719 11815
rect 5733 11781 5767 11815
rect 7665 11781 7699 11815
rect 12449 11781 12483 11815
rect 15301 11781 15335 11815
rect 16037 11781 16071 11815
rect 18613 11781 18647 11815
rect 19349 11781 19383 11815
rect 19993 11781 20027 11815
rect 22661 11781 22695 11815
rect 24409 11781 24443 11815
rect 1501 11713 1535 11747
rect 2421 11713 2455 11747
rect 4537 11713 4571 11747
rect 7389 11713 7423 11747
rect 9597 11713 9631 11747
rect 11621 11713 11655 11747
rect 13185 11713 13219 11747
rect 15945 11713 15979 11747
rect 17417 11713 17451 11747
rect 2145 11645 2179 11679
rect 4721 11645 4755 11679
rect 5917 11645 5951 11679
rect 10333 11645 10367 11679
rect 10977 11645 11011 11679
rect 12541 11645 12575 11679
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 17601 11645 17635 11679
rect 18705 11645 18739 11679
rect 19717 11645 19751 11679
rect 21925 11645 21959 11679
rect 22385 11645 22419 11679
rect 9137 11577 9171 11611
rect 16957 11577 16991 11611
rect 18153 11577 18187 11611
rect 4077 11509 4111 11543
rect 11989 11509 12023 11543
rect 14933 11509 14967 11543
rect 15577 11509 15611 11543
rect 21465 11509 21499 11543
rect 24133 11509 24167 11543
rect 3433 11305 3467 11339
rect 3617 11305 3651 11339
rect 4169 11305 4203 11339
rect 6561 11305 6595 11339
rect 7481 11305 7515 11339
rect 7849 11305 7883 11339
rect 13277 11305 13311 11339
rect 13553 11305 13587 11339
rect 13829 11305 13863 11339
rect 16497 11305 16531 11339
rect 18889 11305 18923 11339
rect 22661 11305 22695 11339
rect 23029 11305 23063 11339
rect 32045 11305 32079 11339
rect 1593 11237 1627 11271
rect 10333 11237 10367 11271
rect 2237 11169 2271 11203
rect 5089 11169 5123 11203
rect 8309 11169 8343 11203
rect 8401 11169 8435 11203
rect 9597 11169 9631 11203
rect 9689 11169 9723 11203
rect 10977 11169 11011 11203
rect 11529 11169 11563 11203
rect 14197 11169 14231 11203
rect 29745 11169 29779 11203
rect 1777 11101 1811 11135
rect 2513 11101 2547 11135
rect 4077 11101 4111 11135
rect 4813 11101 4847 11135
rect 8217 11101 8251 11135
rect 9505 11101 9539 11135
rect 14749 11101 14783 11135
rect 17141 11101 17175 11135
rect 19533 11101 19567 11135
rect 20913 11101 20947 11135
rect 7021 11033 7055 11067
rect 10701 11033 10735 11067
rect 11805 11033 11839 11067
rect 15025 11033 15059 11067
rect 17417 11033 17451 11067
rect 20269 11033 20303 11067
rect 21189 11033 21223 11067
rect 30021 11033 30055 11067
rect 31769 11033 31803 11067
rect 9137 10965 9171 10999
rect 10793 10965 10827 10999
rect 16773 10965 16807 10999
rect 4813 10761 4847 10795
rect 5825 10761 5859 10795
rect 9873 10761 9907 10795
rect 14841 10761 14875 10795
rect 15577 10761 15611 10795
rect 19257 10761 19291 10795
rect 21925 10761 21959 10795
rect 22109 10761 22143 10795
rect 1501 10693 1535 10727
rect 10701 10693 10735 10727
rect 10793 10693 10827 10727
rect 12357 10693 12391 10727
rect 17785 10693 17819 10727
rect 3433 10625 3467 10659
rect 5365 10625 5399 10659
rect 7021 10625 7055 10659
rect 9505 10625 9539 10659
rect 14749 10625 14783 10659
rect 15945 10625 15979 10659
rect 17509 10625 17543 10659
rect 1869 10557 1903 10591
rect 2145 10557 2179 10591
rect 2421 10557 2455 10591
rect 3709 10557 3743 10591
rect 7481 10557 7515 10591
rect 7757 10557 7791 10591
rect 10057 10557 10091 10591
rect 10885 10557 10919 10591
rect 12081 10557 12115 10591
rect 15025 10557 15059 10591
rect 16037 10557 16071 10591
rect 16221 10557 16255 10591
rect 16865 10557 16899 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 4629 10489 4663 10523
rect 6561 10489 6595 10523
rect 21465 10489 21499 10523
rect 1593 10421 1627 10455
rect 5181 10421 5215 10455
rect 6837 10421 6871 10455
rect 10333 10421 10367 10455
rect 11621 10421 11655 10455
rect 13829 10421 13863 10455
rect 14381 10421 14415 10455
rect 2697 10217 2731 10251
rect 3249 10217 3283 10251
rect 5457 10217 5491 10251
rect 9137 10217 9171 10251
rect 10057 10217 10091 10251
rect 14105 10217 14139 10251
rect 16313 10217 16347 10251
rect 18889 10217 18923 10251
rect 21557 10217 21591 10251
rect 3893 10149 3927 10183
rect 6377 10149 6411 10183
rect 6469 10149 6503 10183
rect 8585 10149 8619 10183
rect 1593 10081 1627 10115
rect 1869 10081 1903 10115
rect 4261 10081 4295 10115
rect 4537 10081 4571 10115
rect 6837 10081 6871 10115
rect 10701 10081 10735 10115
rect 13553 10081 13587 10115
rect 14565 10081 14599 10115
rect 14841 10081 14875 10115
rect 19441 10081 19475 10115
rect 2881 10013 2915 10047
rect 3157 10013 3191 10047
rect 3433 10013 3467 10047
rect 5825 10013 5859 10047
rect 9413 10013 9447 10047
rect 11253 10013 11287 10047
rect 17141 10013 17175 10047
rect 7113 9945 7147 9979
rect 11529 9945 11563 9979
rect 17417 9945 17451 9979
rect 19717 9945 19751 9979
rect 21649 9945 21683 9979
rect 10425 9877 10459 9911
rect 10517 9877 10551 9911
rect 13001 9877 13035 9911
rect 16681 9877 16715 9911
rect 16865 9877 16899 9911
rect 21189 9877 21223 9911
rect 6469 9673 6503 9707
rect 16221 9673 16255 9707
rect 1501 9605 1535 9639
rect 1685 9605 1719 9639
rect 3249 9605 3283 9639
rect 5733 9605 5767 9639
rect 5825 9605 5859 9639
rect 10793 9605 10827 9639
rect 11989 9605 12023 9639
rect 13829 9605 13863 9639
rect 13921 9605 13955 9639
rect 17141 9605 17175 9639
rect 19533 9605 19567 9639
rect 28641 9605 28675 9639
rect 2237 9537 2271 9571
rect 3801 9537 3835 9571
rect 4261 9537 4295 9571
rect 7113 9537 7147 9571
rect 10701 9537 10735 9571
rect 19441 9537 19475 9571
rect 27537 9537 27571 9571
rect 1961 9469 1995 9503
rect 4537 9469 4571 9503
rect 6837 9469 6871 9503
rect 8125 9469 8159 9503
rect 8401 9469 8435 9503
rect 10885 9469 10919 9503
rect 11713 9469 11747 9503
rect 14473 9469 14507 9503
rect 14749 9469 14783 9503
rect 16865 9469 16899 9503
rect 19717 9469 19751 9503
rect 27997 9469 28031 9503
rect 3617 9401 3651 9435
rect 13461 9401 13495 9435
rect 14105 9401 14139 9435
rect 19073 9401 19107 9435
rect 5549 9333 5583 9367
rect 9873 9333 9907 9367
rect 10333 9333 10367 9367
rect 18613 9333 18647 9367
rect 20085 9333 20119 9367
rect 27813 9333 27847 9367
rect 28457 9333 28491 9367
rect 3433 9129 3467 9163
rect 4629 9129 4663 9163
rect 5457 9129 5491 9163
rect 5549 9129 5583 9163
rect 7205 9129 7239 9163
rect 7849 9129 7883 9163
rect 10149 9129 10183 9163
rect 11575 9129 11609 9163
rect 3617 9061 3651 9095
rect 5181 9061 5215 9095
rect 14289 9061 14323 9095
rect 1593 8993 1627 9027
rect 1869 8993 1903 9027
rect 4721 8993 4755 9027
rect 6193 8993 6227 9027
rect 8401 8993 8435 9027
rect 9413 8993 9447 9027
rect 10793 8993 10827 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 15485 8993 15519 9027
rect 16037 8993 16071 9027
rect 3065 8925 3099 8959
rect 5917 8925 5951 8959
rect 7389 8925 7423 8959
rect 11345 8925 11379 8959
rect 10517 8857 10551 8891
rect 13553 8857 13587 8891
rect 16313 8857 16347 8891
rect 2881 8789 2915 8823
rect 3985 8789 4019 8823
rect 8217 8789 8251 8823
rect 8309 8789 8343 8823
rect 9045 8789 9079 8823
rect 10609 8789 10643 8823
rect 12633 8789 12667 8823
rect 14657 8789 14691 8823
rect 17785 8789 17819 8823
rect 18153 8789 18187 8823
rect 18705 8789 18739 8823
rect 18981 8789 19015 8823
rect 2881 8585 2915 8619
rect 3433 8585 3467 8619
rect 3525 8585 3559 8619
rect 3985 8585 4019 8619
rect 5825 8585 5859 8619
rect 6469 8585 6503 8619
rect 6653 8585 6687 8619
rect 8033 8585 8067 8619
rect 11161 8585 11195 8619
rect 11529 8585 11563 8619
rect 12173 8585 12207 8619
rect 14289 8585 14323 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 7389 8517 7423 8551
rect 16037 8517 16071 8551
rect 1869 8449 1903 8483
rect 3065 8449 3099 8483
rect 4169 8449 4203 8483
rect 4813 8449 4847 8483
rect 6009 8449 6043 8483
rect 6837 8449 6871 8483
rect 7205 8449 7239 8483
rect 8677 8449 8711 8483
rect 9689 8449 9723 8483
rect 10517 8449 10551 8483
rect 12541 8449 12575 8483
rect 13645 8449 13679 8483
rect 14657 8449 14691 8483
rect 1593 8381 1627 8415
rect 5181 8381 5215 8415
rect 7757 8381 7791 8415
rect 8401 8381 8435 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 12633 8381 12667 8415
rect 12817 8381 12851 8415
rect 14749 8381 14783 8415
rect 14933 8381 14967 8415
rect 16221 8381 16255 8415
rect 4629 8313 4663 8347
rect 9873 8313 9907 8347
rect 7849 8245 7883 8279
rect 10149 8245 10183 8279
rect 1593 8041 1627 8075
rect 2237 8041 2271 8075
rect 2881 8041 2915 8075
rect 3893 8041 3927 8075
rect 4261 8041 4295 8075
rect 4629 8041 4663 8075
rect 7573 8041 7607 8075
rect 9597 8041 9631 8075
rect 12449 8041 12483 8075
rect 13001 8041 13035 8075
rect 3985 7973 4019 8007
rect 15209 7973 15243 8007
rect 7757 7905 7791 7939
rect 10241 7905 10275 7939
rect 11253 7905 11287 7939
rect 13645 7905 13679 7939
rect 14289 7905 14323 7939
rect 14841 7905 14875 7939
rect 1777 7837 1811 7871
rect 2421 7837 2455 7871
rect 3065 7837 3099 7871
rect 4445 7837 4479 7871
rect 10057 7837 10091 7871
rect 14197 7837 14231 7871
rect 15025 7837 15059 7871
rect 3433 7769 3467 7803
rect 9229 7769 9263 7803
rect 9965 7769 9999 7803
rect 3525 7701 3559 7735
rect 11483 7701 11517 7735
rect 13369 7701 13403 7735
rect 13461 7701 13495 7735
rect 15853 7701 15887 7735
rect 1593 7497 1627 7531
rect 4353 7497 4387 7531
rect 9137 7497 9171 7531
rect 11897 7497 11931 7531
rect 13461 7497 13495 7531
rect 23949 7497 23983 7531
rect 1777 7361 1811 7395
rect 2421 7361 2455 7395
rect 3065 7361 3099 7395
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 9321 7361 9355 7395
rect 10793 7361 10827 7395
rect 12725 7361 12759 7395
rect 14289 7361 14323 7395
rect 22201 7361 22235 7395
rect 24225 7361 24259 7395
rect 4169 7293 4203 7327
rect 22477 7293 22511 7327
rect 2237 7225 2271 7259
rect 2881 7225 2915 7259
rect 3525 7157 3559 7191
rect 10609 7157 10643 7191
rect 12541 7157 12575 7191
rect 14105 7157 14139 7191
rect 3433 6953 3467 6987
rect 23213 6953 23247 6987
rect 2881 6885 2915 6919
rect 23765 6885 23799 6919
rect 4169 6817 4203 6851
rect 10609 6817 10643 6851
rect 1777 6749 1811 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 3525 6749 3559 6783
rect 22937 6749 22971 6783
rect 3801 6681 3835 6715
rect 1593 6613 1627 6647
rect 2237 6613 2271 6647
rect 3985 6613 4019 6647
rect 23397 6613 23431 6647
rect 2881 6409 2915 6443
rect 22845 6409 22879 6443
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 22452 6273 22486 6307
rect 1593 6205 1627 6239
rect 1869 6205 1903 6239
rect 22523 6069 22557 6103
rect 2697 5865 2731 5899
rect 18889 5865 18923 5899
rect 21005 5865 21039 5899
rect 21741 5797 21775 5831
rect 1869 5729 1903 5763
rect 15577 5729 15611 5763
rect 17141 5729 17175 5763
rect 24869 5729 24903 5763
rect 26985 5729 27019 5763
rect 28825 5729 28859 5763
rect 1593 5661 1627 5695
rect 2881 5661 2915 5695
rect 15761 5661 15795 5695
rect 19349 5661 19383 5695
rect 20913 5661 20947 5695
rect 24685 5661 24719 5695
rect 17417 5593 17451 5627
rect 26525 5593 26559 5627
rect 27169 5593 27203 5627
rect 16221 5525 16255 5559
rect 21373 5525 21407 5559
rect 22891 5321 22925 5355
rect 1593 5185 1627 5219
rect 2697 5185 2731 5219
rect 15669 5185 15703 5219
rect 17509 5185 17543 5219
rect 22176 5185 22210 5219
rect 22788 5185 22822 5219
rect 1869 5117 1903 5151
rect 15853 5117 15887 5151
rect 17693 5117 17727 5151
rect 28641 5117 28675 5151
rect 28825 5117 28859 5151
rect 30021 5117 30055 5151
rect 16313 4981 16347 5015
rect 18153 4981 18187 5015
rect 22247 4981 22281 5015
rect 19533 4777 19567 4811
rect 20269 4777 20303 4811
rect 24731 4777 24765 4811
rect 1593 4641 1627 4675
rect 1869 4641 1903 4675
rect 25789 4641 25823 4675
rect 2881 4573 2915 4607
rect 19441 4573 19475 4607
rect 24628 4573 24662 4607
rect 27629 4573 27663 4607
rect 25973 4505 26007 4539
rect 2789 4437 2823 4471
rect 19901 4437 19935 4471
rect 2237 4233 2271 4267
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 3065 4097 3099 4131
rect 3341 4097 3375 4131
rect 15209 4097 15243 4131
rect 3525 3961 3559 3995
rect 1593 3893 1627 3927
rect 2881 3893 2915 3927
rect 15025 3893 15059 3927
rect 12081 3689 12115 3723
rect 3525 3621 3559 3655
rect 1869 3553 1903 3587
rect 1593 3485 1627 3519
rect 3065 3485 3099 3519
rect 3341 3485 3375 3519
rect 11529 3417 11563 3451
rect 2881 3349 2915 3383
rect 3801 3349 3835 3383
rect 11621 3349 11655 3383
rect 14013 3145 14047 3179
rect 10793 3077 10827 3111
rect 12633 3077 12667 3111
rect 13921 3077 13955 3111
rect 15577 3077 15611 3111
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 4169 3009 4203 3043
rect 6561 3009 6595 3043
rect 8769 3009 8803 3043
rect 17049 3009 17083 3043
rect 18337 3009 18371 3043
rect 20545 3009 20579 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 7205 2941 7239 2975
rect 9045 2941 9079 2975
rect 10517 2941 10551 2975
rect 3985 2873 4019 2907
rect 15761 2873 15795 2907
rect 12725 2805 12759 2839
rect 16865 2805 16899 2839
rect 18153 2805 18187 2839
rect 20361 2805 20395 2839
rect 3341 2601 3375 2635
rect 3801 2601 3835 2635
rect 25513 2601 25547 2635
rect 28181 2601 28215 2635
rect 30849 2601 30883 2635
rect 33517 2601 33551 2635
rect 2881 2533 2915 2567
rect 1593 2465 1627 2499
rect 4629 2465 4663 2499
rect 7297 2465 7331 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 15301 2465 15335 2499
rect 17969 2465 18003 2499
rect 20545 2465 20579 2499
rect 23121 2465 23155 2499
rect 36369 2465 36403 2499
rect 3065 2397 3099 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 9597 2397 9631 2431
rect 12357 2397 12391 2431
rect 15025 2397 15059 2431
rect 17509 2397 17543 2431
rect 20085 2397 20119 2431
rect 22661 2397 22695 2431
rect 25697 2397 25731 2431
rect 25973 2397 26007 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33701 2397 33735 2431
rect 33977 2397 34011 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
rect 3525 2329 3559 2363
rect 1823 2261 1857 2295
<< metal1 >>
rect 8294 26324 8300 26376
rect 8352 26364 8358 26376
rect 23382 26364 23388 26376
rect 8352 26336 23388 26364
rect 8352 26324 8358 26336
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 12066 25712 12072 25764
rect 12124 25752 12130 25764
rect 33962 25752 33968 25764
rect 12124 25724 33968 25752
rect 12124 25712 12130 25724
rect 33962 25712 33968 25724
rect 34020 25712 34026 25764
rect 10594 25644 10600 25696
rect 10652 25684 10658 25696
rect 26878 25684 26884 25696
rect 10652 25656 26884 25684
rect 10652 25644 10658 25656
rect 26878 25644 26884 25656
rect 26936 25644 26942 25696
rect 13722 25576 13728 25628
rect 13780 25616 13786 25628
rect 34882 25616 34888 25628
rect 13780 25588 34888 25616
rect 13780 25576 13786 25588
rect 34882 25576 34888 25588
rect 34940 25576 34946 25628
rect 10042 25508 10048 25560
rect 10100 25548 10106 25560
rect 33594 25548 33600 25560
rect 10100 25520 33600 25548
rect 10100 25508 10106 25520
rect 33594 25508 33600 25520
rect 33652 25508 33658 25560
rect 10778 25440 10784 25492
rect 10836 25480 10842 25492
rect 34974 25480 34980 25492
rect 10836 25452 34980 25480
rect 10836 25440 10842 25452
rect 34974 25440 34980 25452
rect 35032 25440 35038 25492
rect 14642 25372 14648 25424
rect 14700 25412 14706 25424
rect 31110 25412 31116 25424
rect 14700 25384 31116 25412
rect 14700 25372 14706 25384
rect 31110 25372 31116 25384
rect 31168 25372 31174 25424
rect 12250 25304 12256 25356
rect 12308 25344 12314 25356
rect 32306 25344 32312 25356
rect 12308 25316 32312 25344
rect 12308 25304 12314 25316
rect 32306 25304 32312 25316
rect 32364 25304 32370 25356
rect 13906 25236 13912 25288
rect 13964 25276 13970 25288
rect 32490 25276 32496 25288
rect 13964 25248 32496 25276
rect 13964 25236 13970 25248
rect 32490 25236 32496 25248
rect 32548 25236 32554 25288
rect 4062 25168 4068 25220
rect 4120 25208 4126 25220
rect 9122 25208 9128 25220
rect 4120 25180 9128 25208
rect 4120 25168 4126 25180
rect 9122 25168 9128 25180
rect 9180 25168 9186 25220
rect 10410 25168 10416 25220
rect 10468 25208 10474 25220
rect 30190 25208 30196 25220
rect 10468 25180 30196 25208
rect 10468 25168 10474 25180
rect 30190 25168 30196 25180
rect 30248 25168 30254 25220
rect 16666 25100 16672 25152
rect 16724 25140 16730 25152
rect 28534 25140 28540 25152
rect 16724 25112 28540 25140
rect 16724 25100 16730 25112
rect 28534 25100 28540 25112
rect 28592 25100 28598 25152
rect 15654 25032 15660 25084
rect 15712 25072 15718 25084
rect 30374 25072 30380 25084
rect 15712 25044 30380 25072
rect 15712 25032 15718 25044
rect 30374 25032 30380 25044
rect 30432 25032 30438 25084
rect 15930 24964 15936 25016
rect 15988 25004 15994 25016
rect 32858 25004 32864 25016
rect 15988 24976 32864 25004
rect 15988 24964 15994 24976
rect 32858 24964 32864 24976
rect 32916 24964 32922 25016
rect 15194 24896 15200 24948
rect 15252 24936 15258 24948
rect 15252 24908 21680 24936
rect 15252 24896 15258 24908
rect 14734 24828 14740 24880
rect 14792 24868 14798 24880
rect 21542 24868 21548 24880
rect 14792 24840 21548 24868
rect 14792 24828 14798 24840
rect 21542 24828 21548 24840
rect 21600 24828 21606 24880
rect 21652 24868 21680 24908
rect 21910 24896 21916 24948
rect 21968 24936 21974 24948
rect 39298 24936 39304 24948
rect 21968 24908 39304 24936
rect 21968 24896 21974 24908
rect 39298 24896 39304 24908
rect 39356 24896 39362 24948
rect 33502 24868 33508 24880
rect 21652 24840 33508 24868
rect 33502 24828 33508 24840
rect 33560 24828 33566 24880
rect 6546 24760 6552 24812
rect 6604 24800 6610 24812
rect 13538 24800 13544 24812
rect 6604 24772 13544 24800
rect 6604 24760 6610 24772
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 14274 24760 14280 24812
rect 14332 24800 14338 24812
rect 26142 24800 26148 24812
rect 14332 24772 26148 24800
rect 14332 24760 14338 24772
rect 26142 24760 26148 24772
rect 26200 24760 26206 24812
rect 26234 24760 26240 24812
rect 26292 24800 26298 24812
rect 29178 24800 29184 24812
rect 26292 24772 29184 24800
rect 26292 24760 26298 24772
rect 29178 24760 29184 24772
rect 29236 24760 29242 24812
rect 3786 24692 3792 24744
rect 3844 24732 3850 24744
rect 12618 24732 12624 24744
rect 3844 24704 12624 24732
rect 3844 24692 3850 24704
rect 12618 24692 12624 24704
rect 12676 24732 12682 24744
rect 13722 24732 13728 24744
rect 12676 24704 13728 24732
rect 12676 24692 12682 24704
rect 13722 24692 13728 24704
rect 13780 24692 13786 24744
rect 19058 24692 19064 24744
rect 19116 24732 19122 24744
rect 26418 24732 26424 24744
rect 19116 24704 26424 24732
rect 19116 24692 19122 24704
rect 26418 24692 26424 24704
rect 26476 24692 26482 24744
rect 27246 24692 27252 24744
rect 27304 24732 27310 24744
rect 27304 24704 30604 24732
rect 27304 24692 27310 24704
rect 4062 24624 4068 24676
rect 4120 24664 4126 24676
rect 7282 24664 7288 24676
rect 4120 24636 7288 24664
rect 4120 24624 4126 24636
rect 7282 24624 7288 24636
rect 7340 24624 7346 24676
rect 12342 24624 12348 24676
rect 12400 24664 12406 24676
rect 25774 24664 25780 24676
rect 12400 24636 25780 24664
rect 12400 24624 12406 24636
rect 25774 24624 25780 24636
rect 25832 24624 25838 24676
rect 26050 24624 26056 24676
rect 26108 24664 26114 24676
rect 30466 24664 30472 24676
rect 26108 24636 30472 24664
rect 26108 24624 26114 24636
rect 30466 24624 30472 24636
rect 30524 24624 30530 24676
rect 30576 24664 30604 24704
rect 31294 24692 31300 24744
rect 31352 24732 31358 24744
rect 36630 24732 36636 24744
rect 31352 24704 36636 24732
rect 31352 24692 31358 24704
rect 36630 24692 36636 24704
rect 36688 24692 36694 24744
rect 31662 24664 31668 24676
rect 30576 24636 31668 24664
rect 31662 24624 31668 24636
rect 31720 24624 31726 24676
rect 11698 24556 11704 24608
rect 11756 24596 11762 24608
rect 21726 24596 21732 24608
rect 11756 24568 21732 24596
rect 11756 24556 11762 24568
rect 21726 24556 21732 24568
rect 21784 24556 21790 24608
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 30006 24596 30012 24608
rect 21968 24568 30012 24596
rect 21968 24556 21974 24568
rect 30006 24556 30012 24568
rect 30064 24556 30070 24608
rect 30374 24556 30380 24608
rect 30432 24596 30438 24608
rect 34146 24596 34152 24608
rect 30432 24568 34152 24596
rect 30432 24556 30438 24568
rect 34146 24556 34152 24568
rect 34204 24556 34210 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 4890 24392 4896 24404
rect 2832 24364 4896 24392
rect 2832 24352 2838 24364
rect 4890 24352 4896 24364
rect 4948 24352 4954 24404
rect 6546 24352 6552 24404
rect 6604 24352 6610 24404
rect 9125 24395 9183 24401
rect 9125 24361 9137 24395
rect 9171 24392 9183 24395
rect 11054 24392 11060 24404
rect 9171 24364 11060 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 11054 24352 11060 24364
rect 11112 24352 11118 24404
rect 11698 24352 11704 24404
rect 11756 24352 11762 24404
rect 14274 24352 14280 24404
rect 14332 24352 14338 24404
rect 18966 24392 18972 24404
rect 16776 24364 18972 24392
rect 3973 24327 4031 24333
rect 3973 24293 3985 24327
rect 4019 24324 4031 24327
rect 11974 24324 11980 24336
rect 4019 24296 11980 24324
rect 4019 24293 4031 24296
rect 3973 24287 4031 24293
rect 11974 24284 11980 24296
rect 12032 24284 12038 24336
rect 14458 24324 14464 24336
rect 13556 24296 14464 24324
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 5813 24259 5871 24265
rect 3804 24228 5764 24256
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2406 24188 2412 24200
rect 2271 24160 2412 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2406 24148 2412 24160
rect 2464 24148 2470 24200
rect 3418 24148 3424 24200
rect 3476 24188 3482 24200
rect 3804 24188 3832 24228
rect 3476 24160 3832 24188
rect 3881 24191 3939 24197
rect 3476 24148 3482 24160
rect 3881 24157 3893 24191
rect 3927 24188 3939 24191
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 3927 24160 4169 24188
rect 3927 24157 3939 24160
rect 3881 24151 3939 24157
rect 4157 24157 4169 24160
rect 4203 24188 4215 24191
rect 4246 24188 4252 24200
rect 4203 24160 4252 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4246 24148 4252 24160
rect 4304 24148 4310 24200
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 1762 24080 1768 24132
rect 1820 24120 1826 24132
rect 4632 24120 4660 24151
rect 1820 24092 4660 24120
rect 1820 24080 1826 24092
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 1673 24055 1731 24061
rect 1673 24052 1685 24055
rect 1627 24024 1685 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 1673 24021 1685 24024
rect 1719 24052 1731 24055
rect 3694 24052 3700 24064
rect 1719 24024 3700 24052
rect 1719 24021 1731 24024
rect 1673 24015 1731 24021
rect 3694 24012 3700 24024
rect 3752 24012 3758 24064
rect 5736 24052 5764 24228
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6822 24256 6828 24268
rect 5859 24228 6828 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9214 24256 9220 24268
rect 8251 24228 9220 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9214 24216 9220 24228
rect 9272 24216 9278 24268
rect 13556 24265 13584 24296
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 13541 24259 13599 24265
rect 12406 24228 12756 24256
rect 6457 24191 6515 24197
rect 6457 24157 6469 24191
rect 6503 24188 6515 24191
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 6503 24160 6745 24188
rect 6503 24157 6515 24160
rect 6457 24151 6515 24157
rect 6733 24157 6745 24160
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 7377 24191 7435 24197
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 8386 24188 8392 24200
rect 7423 24160 8392 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 6748 24120 6776 24151
rect 8386 24148 8392 24160
rect 8444 24148 8450 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10594 24188 10600 24200
rect 9999 24160 10600 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 8294 24120 8300 24132
rect 6748 24092 8300 24120
rect 8294 24080 8300 24092
rect 8352 24080 8358 24132
rect 9214 24052 9220 24064
rect 5736 24024 9220 24052
rect 9214 24012 9220 24024
rect 9272 24012 9278 24064
rect 9324 24052 9352 24151
rect 10594 24148 10600 24160
rect 10652 24148 10658 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 12406 24188 12434 24228
rect 11931 24160 12434 24188
rect 12529 24191 12587 24197
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12618 24188 12624 24200
rect 12575 24160 12624 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12618 24148 12624 24160
rect 12676 24148 12682 24200
rect 12728 24188 12756 24228
rect 13541 24225 13553 24259
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 16776 24256 16804 24364
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 25130 24392 25136 24404
rect 19306 24364 25136 24392
rect 18414 24284 18420 24336
rect 18472 24324 18478 24336
rect 19306 24324 19334 24364
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 25240 24364 25452 24392
rect 25240 24324 25268 24364
rect 18472 24296 19334 24324
rect 25148 24296 25268 24324
rect 25424 24324 25452 24364
rect 25774 24352 25780 24404
rect 25832 24352 25838 24404
rect 27154 24352 27160 24404
rect 27212 24352 27218 24404
rect 29086 24392 29092 24404
rect 27264 24364 29092 24392
rect 27264 24324 27292 24364
rect 29086 24352 29092 24364
rect 29144 24352 29150 24404
rect 31570 24392 31576 24404
rect 29196 24364 31576 24392
rect 25424 24296 27292 24324
rect 18472 24284 18478 24296
rect 16163 24228 16804 24256
rect 16853 24259 16911 24265
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 18690 24256 18696 24268
rect 16899 24228 18696 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 18966 24216 18972 24268
rect 19024 24256 19030 24268
rect 19242 24256 19248 24268
rect 19024 24228 19248 24256
rect 19024 24216 19030 24228
rect 19242 24216 19248 24228
rect 19300 24216 19306 24268
rect 19886 24216 19892 24268
rect 19944 24256 19950 24268
rect 20806 24256 20812 24268
rect 19944 24228 20812 24256
rect 19944 24216 19950 24228
rect 20806 24216 20812 24228
rect 20864 24216 20870 24268
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 22094 24216 22100 24268
rect 22152 24256 22158 24268
rect 25148 24265 25176 24296
rect 27614 24284 27620 24336
rect 27672 24324 27678 24336
rect 28997 24327 29055 24333
rect 28997 24324 29009 24327
rect 27672 24296 29009 24324
rect 27672 24284 27678 24296
rect 28997 24293 29009 24296
rect 29043 24293 29055 24327
rect 28997 24287 29055 24293
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 22152 24228 22477 24256
rect 22152 24216 22158 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 25222 24216 25228 24268
rect 25280 24256 25286 24268
rect 26329 24259 26387 24265
rect 26329 24256 26341 24259
rect 25280 24228 26341 24256
rect 25280 24216 25286 24228
rect 26329 24225 26341 24228
rect 26375 24225 26387 24259
rect 26329 24219 26387 24225
rect 26418 24216 26424 24268
rect 26476 24256 26482 24268
rect 27709 24259 27767 24265
rect 27709 24256 27721 24259
rect 26476 24228 27721 24256
rect 26476 24216 26482 24228
rect 27709 24225 27721 24228
rect 27755 24225 27767 24259
rect 29196 24256 29224 24364
rect 31570 24352 31576 24364
rect 31628 24352 31634 24404
rect 31662 24352 31668 24404
rect 31720 24392 31726 24404
rect 32309 24395 32367 24401
rect 32309 24392 32321 24395
rect 31720 24364 32321 24392
rect 31720 24352 31726 24364
rect 32309 24361 32321 24364
rect 32355 24361 32367 24395
rect 32309 24355 32367 24361
rect 34146 24352 34152 24404
rect 34204 24352 34210 24404
rect 37921 24395 37979 24401
rect 37921 24392 37933 24395
rect 35268 24364 37933 24392
rect 29748 24296 30328 24324
rect 27709 24219 27767 24225
rect 28552 24228 29224 24256
rect 12728 24160 14044 24188
rect 10965 24123 11023 24129
rect 10965 24089 10977 24123
rect 11011 24120 11023 24123
rect 13814 24120 13820 24132
rect 11011 24092 13820 24120
rect 11011 24089 11023 24092
rect 10965 24083 11023 24089
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 14016 24120 14044 24160
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 15378 24188 15384 24200
rect 15151 24160 15384 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 15378 24148 15384 24160
rect 15436 24148 15442 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 19978 24188 19984 24200
rect 19659 24160 19984 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 19978 24148 19984 24160
rect 20036 24148 20042 24200
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 15838 24120 15844 24132
rect 14016 24092 15844 24120
rect 15838 24080 15844 24092
rect 15896 24080 15902 24132
rect 17126 24080 17132 24132
rect 17184 24080 17190 24132
rect 17586 24080 17592 24132
rect 17644 24080 17650 24132
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 20088 24120 20116 24151
rect 21726 24148 21732 24200
rect 21784 24188 21790 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21784 24160 22017 24188
rect 21784 24148 21790 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 23934 24148 23940 24200
rect 23992 24188 23998 24200
rect 24029 24191 24087 24197
rect 24029 24188 24041 24191
rect 23992 24160 24041 24188
rect 23992 24148 23998 24160
rect 24029 24157 24041 24160
rect 24075 24188 24087 24191
rect 24946 24188 24952 24200
rect 24075 24160 24952 24188
rect 24075 24157 24087 24160
rect 24029 24151 24087 24157
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 25041 24191 25099 24197
rect 25041 24157 25053 24191
rect 25087 24188 25099 24191
rect 26050 24188 26056 24200
rect 25087 24160 26056 24188
rect 25087 24157 25099 24160
rect 25041 24151 25099 24157
rect 26050 24148 26056 24160
rect 26108 24148 26114 24200
rect 26142 24148 26148 24200
rect 26200 24188 26206 24200
rect 28552 24197 28580 24228
rect 29270 24216 29276 24268
rect 29328 24256 29334 24268
rect 29748 24265 29776 24296
rect 29733 24259 29791 24265
rect 29733 24256 29745 24259
rect 29328 24228 29745 24256
rect 29328 24216 29334 24228
rect 29733 24225 29745 24228
rect 29779 24225 29791 24259
rect 29733 24219 29791 24225
rect 30006 24216 30012 24268
rect 30064 24216 30070 24268
rect 30300 24256 30328 24296
rect 30650 24284 30656 24336
rect 30708 24324 30714 24336
rect 33870 24324 33876 24336
rect 30708 24296 33876 24324
rect 30708 24284 30714 24296
rect 33870 24284 33876 24296
rect 33928 24284 33934 24336
rect 34054 24284 34060 24336
rect 34112 24324 34118 24336
rect 35268 24324 35296 24364
rect 37921 24361 37933 24364
rect 37967 24361 37979 24395
rect 37921 24355 37979 24361
rect 39298 24352 39304 24404
rect 39356 24352 39362 24404
rect 44726 24352 44732 24404
rect 44784 24352 44790 24404
rect 34112 24296 35296 24324
rect 34112 24284 34118 24296
rect 35894 24284 35900 24336
rect 35952 24284 35958 24336
rect 36906 24284 36912 24336
rect 36964 24324 36970 24336
rect 37461 24327 37519 24333
rect 37461 24324 37473 24327
rect 36964 24296 37473 24324
rect 36964 24284 36970 24296
rect 37461 24293 37473 24296
rect 37507 24293 37519 24327
rect 37461 24287 37519 24293
rect 37001 24259 37059 24265
rect 37001 24256 37013 24259
rect 30300 24228 37013 24256
rect 37001 24225 37013 24228
rect 37047 24225 37059 24259
rect 37001 24219 37059 24225
rect 39574 24216 39580 24268
rect 39632 24256 39638 24268
rect 40037 24259 40095 24265
rect 40037 24256 40049 24259
rect 39632 24228 40049 24256
rect 39632 24216 39638 24228
rect 40037 24225 40049 24228
rect 40083 24225 40095 24259
rect 40037 24219 40095 24225
rect 40126 24216 40132 24268
rect 40184 24256 40190 24268
rect 40313 24259 40371 24265
rect 40313 24256 40325 24259
rect 40184 24228 40325 24256
rect 40184 24216 40190 24228
rect 40313 24225 40325 24228
rect 40359 24225 40371 24259
rect 40313 24219 40371 24225
rect 26237 24191 26295 24197
rect 26237 24188 26249 24191
rect 26200 24160 26249 24188
rect 26200 24148 26206 24160
rect 26237 24157 26249 24160
rect 26283 24157 26295 24191
rect 26237 24151 26295 24157
rect 27525 24191 27583 24197
rect 27525 24157 27537 24191
rect 27571 24188 27583 24191
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 27571 24160 27752 24188
rect 27571 24157 27583 24160
rect 27525 24151 27583 24157
rect 27724 24132 27752 24160
rect 28276 24160 28549 24188
rect 27617 24123 27675 24129
rect 27617 24120 27629 24123
rect 19392 24092 20116 24120
rect 23860 24092 27629 24120
rect 19392 24080 19398 24092
rect 16758 24052 16764 24064
rect 9324 24024 16764 24052
rect 16758 24012 16764 24024
rect 16816 24012 16822 24064
rect 17402 24012 17408 24064
rect 17460 24052 17466 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 17460 24024 18613 24052
rect 17460 24012 17466 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 18601 24015 18659 24021
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 20438 24052 20444 24064
rect 19475 24024 20444 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 20438 24012 20444 24024
rect 20496 24012 20502 24064
rect 23860 24061 23888 24092
rect 27617 24089 27629 24092
rect 27663 24089 27675 24123
rect 27617 24083 27675 24089
rect 27706 24080 27712 24132
rect 27764 24080 27770 24132
rect 23845 24055 23903 24061
rect 23845 24021 23857 24055
rect 23891 24021 23903 24055
rect 23845 24015 23903 24021
rect 24026 24012 24032 24064
rect 24084 24052 24090 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 24084 24024 24593 24052
rect 24084 24012 24090 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 24946 24012 24952 24064
rect 25004 24012 25010 24064
rect 26050 24012 26056 24064
rect 26108 24052 26114 24064
rect 26145 24055 26203 24061
rect 26145 24052 26157 24055
rect 26108 24024 26157 24052
rect 26108 24012 26114 24024
rect 26145 24021 26157 24024
rect 26191 24021 26203 24055
rect 26145 24015 26203 24021
rect 26970 24012 26976 24064
rect 27028 24052 27034 24064
rect 28276 24052 28304 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 29178 24148 29184 24200
rect 29236 24188 29242 24200
rect 29914 24188 29920 24200
rect 29236 24160 29920 24188
rect 29236 24148 29242 24160
rect 29914 24148 29920 24160
rect 29972 24148 29978 24200
rect 30558 24148 30564 24200
rect 30616 24188 30622 24200
rect 31481 24191 31539 24197
rect 31481 24188 31493 24191
rect 30616 24160 31493 24188
rect 30616 24148 30622 24160
rect 31481 24157 31493 24160
rect 31527 24157 31539 24191
rect 31481 24151 31539 24157
rect 30929 24123 30987 24129
rect 30929 24089 30941 24123
rect 30975 24120 30987 24123
rect 31496 24120 31524 24151
rect 31846 24148 31852 24200
rect 31904 24188 31910 24200
rect 32493 24191 32551 24197
rect 32493 24188 32505 24191
rect 31904 24160 32505 24188
rect 31904 24148 31910 24160
rect 32493 24157 32505 24160
rect 32539 24188 32551 24191
rect 32674 24188 32680 24200
rect 32539 24160 32680 24188
rect 32539 24157 32551 24160
rect 32493 24151 32551 24157
rect 32674 24148 32680 24160
rect 32732 24148 32738 24200
rect 33318 24148 33324 24200
rect 33376 24148 33382 24200
rect 34054 24148 34060 24200
rect 34112 24148 34118 24200
rect 34514 24148 34520 24200
rect 34572 24188 34578 24200
rect 34977 24191 35035 24197
rect 34977 24188 34989 24191
rect 34572 24160 34989 24188
rect 34572 24148 34578 24160
rect 34977 24157 34989 24160
rect 35023 24188 35035 24191
rect 35618 24188 35624 24200
rect 35023 24160 35624 24188
rect 35023 24157 35035 24160
rect 34977 24151 35035 24157
rect 35618 24148 35624 24160
rect 35676 24148 35682 24200
rect 35894 24148 35900 24200
rect 35952 24188 35958 24200
rect 36541 24191 36599 24197
rect 36541 24188 36553 24191
rect 35952 24160 36553 24188
rect 35952 24148 35958 24160
rect 36541 24157 36553 24160
rect 36587 24188 36599 24191
rect 36814 24188 36820 24200
rect 36587 24160 36820 24188
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 36814 24148 36820 24160
rect 36872 24148 36878 24200
rect 37274 24148 37280 24200
rect 37332 24188 37338 24200
rect 37645 24191 37703 24197
rect 37645 24188 37657 24191
rect 37332 24160 37657 24188
rect 37332 24148 37338 24160
rect 37645 24157 37657 24160
rect 37691 24157 37703 24191
rect 37645 24151 37703 24157
rect 38470 24148 38476 24200
rect 38528 24148 38534 24200
rect 38654 24148 38660 24200
rect 38712 24148 38718 24200
rect 39206 24148 39212 24200
rect 39264 24148 39270 24200
rect 41417 24191 41475 24197
rect 41417 24157 41429 24191
rect 41463 24188 41475 24191
rect 41506 24188 41512 24200
rect 41463 24160 41512 24188
rect 41463 24157 41475 24160
rect 41417 24151 41475 24157
rect 41506 24148 41512 24160
rect 41564 24148 41570 24200
rect 42797 24191 42855 24197
rect 42797 24157 42809 24191
rect 42843 24188 42855 24191
rect 43254 24188 43260 24200
rect 42843 24160 43260 24188
rect 42843 24157 42855 24160
rect 42797 24151 42855 24157
rect 43254 24148 43260 24160
rect 43312 24148 43318 24200
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44784 24160 45201 24188
rect 44784 24148 44790 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45925 24191 45983 24197
rect 45925 24188 45937 24191
rect 45612 24160 45937 24188
rect 45612 24148 45618 24160
rect 45925 24157 45937 24160
rect 45971 24157 45983 24191
rect 45925 24151 45983 24157
rect 46014 24148 46020 24200
rect 46072 24188 46078 24200
rect 46661 24191 46719 24197
rect 46661 24188 46673 24191
rect 46072 24160 46673 24188
rect 46072 24148 46078 24160
rect 46661 24157 46673 24160
rect 46707 24188 46719 24191
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 46707 24160 47225 24188
rect 46707 24157 46719 24160
rect 46661 24151 46719 24157
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 47765 24191 47823 24197
rect 47765 24188 47777 24191
rect 47360 24160 47777 24188
rect 47360 24148 47366 24160
rect 47765 24157 47777 24160
rect 47811 24157 47823 24191
rect 47765 24151 47823 24157
rect 48590 24148 48596 24200
rect 48648 24148 48654 24200
rect 31570 24120 31576 24132
rect 30975 24092 31432 24120
rect 31496 24092 31576 24120
rect 30975 24089 30987 24092
rect 30929 24083 30987 24089
rect 27028 24024 28304 24052
rect 27028 24012 27034 24024
rect 28350 24012 28356 24064
rect 28408 24012 28414 24064
rect 29086 24012 29092 24064
rect 29144 24052 29150 24064
rect 31297 24055 31355 24061
rect 31297 24052 31309 24055
rect 29144 24024 31309 24052
rect 29144 24012 29150 24024
rect 31297 24021 31309 24024
rect 31343 24021 31355 24055
rect 31404 24052 31432 24092
rect 31570 24080 31576 24092
rect 31628 24080 31634 24132
rect 31662 24080 31668 24132
rect 31720 24120 31726 24132
rect 32769 24123 32827 24129
rect 32769 24120 32781 24123
rect 31720 24092 32781 24120
rect 31720 24080 31726 24092
rect 32769 24089 32781 24092
rect 32815 24089 32827 24123
rect 32769 24083 32827 24089
rect 35158 24080 35164 24132
rect 35216 24120 35222 24132
rect 35713 24123 35771 24129
rect 35713 24120 35725 24123
rect 35216 24092 35725 24120
rect 35216 24080 35222 24092
rect 35713 24089 35725 24092
rect 35759 24120 35771 24123
rect 36262 24120 36268 24132
rect 35759 24092 36268 24120
rect 35759 24089 35771 24092
rect 35713 24083 35771 24089
rect 36262 24080 36268 24092
rect 36320 24080 36326 24132
rect 36630 24080 36636 24132
rect 36688 24120 36694 24132
rect 36688 24092 45554 24120
rect 36688 24080 36694 24092
rect 31846 24052 31852 24064
rect 31404 24024 31852 24052
rect 31297 24015 31355 24021
rect 31846 24012 31852 24024
rect 31904 24012 31910 24064
rect 33410 24012 33416 24064
rect 33468 24012 33474 24064
rect 35066 24012 35072 24064
rect 35124 24012 35130 24064
rect 35250 24012 35256 24064
rect 35308 24052 35314 24064
rect 36357 24055 36415 24061
rect 36357 24052 36369 24055
rect 35308 24024 36369 24052
rect 35308 24012 35314 24024
rect 36357 24021 36369 24024
rect 36403 24021 36415 24055
rect 36357 24015 36415 24021
rect 36446 24012 36452 24064
rect 36504 24052 36510 24064
rect 36817 24055 36875 24061
rect 36817 24052 36829 24055
rect 36504 24024 36829 24052
rect 36504 24012 36510 24024
rect 36817 24021 36829 24024
rect 36863 24021 36875 24055
rect 36817 24015 36875 24021
rect 42058 24012 42064 24064
rect 42116 24012 42122 24064
rect 42610 24012 42616 24064
rect 42668 24012 42674 24064
rect 45370 24012 45376 24064
rect 45428 24012 45434 24064
rect 45526 24052 45554 24092
rect 46109 24055 46167 24061
rect 46109 24052 46121 24055
rect 45526 24024 46121 24052
rect 46109 24021 46121 24024
rect 46155 24021 46167 24055
rect 46109 24015 46167 24021
rect 46842 24012 46848 24064
rect 46900 24012 46906 24064
rect 47026 24012 47032 24064
rect 47084 24052 47090 24064
rect 47949 24055 48007 24061
rect 47949 24052 47961 24055
rect 47084 24024 47961 24052
rect 47084 24012 47090 24024
rect 47949 24021 47961 24024
rect 47995 24021 48007 24055
rect 47949 24015 48007 24021
rect 48682 24012 48688 24064
rect 48740 24052 48746 24064
rect 49237 24055 49295 24061
rect 49237 24052 49249 24055
rect 48740 24024 49249 24052
rect 48740 24012 48746 24024
rect 49237 24021 49249 24024
rect 49283 24021 49295 24055
rect 49237 24015 49295 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 1765 23851 1823 23857
rect 1765 23817 1777 23851
rect 1811 23848 1823 23851
rect 3418 23848 3424 23860
rect 1811 23820 3424 23848
rect 1811 23817 1823 23820
rect 1765 23811 1823 23817
rect 3418 23808 3424 23820
rect 3476 23808 3482 23860
rect 5994 23848 6000 23860
rect 3896 23820 6000 23848
rect 1581 23783 1639 23789
rect 1581 23749 1593 23783
rect 1627 23780 1639 23783
rect 3896 23780 3924 23820
rect 5994 23808 6000 23820
rect 6052 23808 6058 23860
rect 6638 23808 6644 23860
rect 6696 23848 6702 23860
rect 12250 23848 12256 23860
rect 6696 23820 12256 23848
rect 6696 23808 6702 23820
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12342 23808 12348 23860
rect 12400 23808 12406 23860
rect 12434 23808 12440 23860
rect 12492 23848 12498 23860
rect 21910 23848 21916 23860
rect 12492 23820 21916 23848
rect 12492 23808 12498 23820
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 23842 23848 23848 23860
rect 23400 23820 23848 23848
rect 1627 23752 3924 23780
rect 3973 23783 4031 23789
rect 1627 23749 1639 23752
rect 1581 23743 1639 23749
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4062 23780 4068 23792
rect 4019 23752 4068 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4062 23740 4068 23752
rect 4120 23740 4126 23792
rect 8570 23780 8576 23792
rect 4172 23752 8576 23780
rect 2130 23672 2136 23724
rect 2188 23672 2194 23724
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3510 23712 3516 23724
rect 3007 23684 3516 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 4062 23604 4068 23656
rect 4120 23644 4126 23656
rect 4172 23644 4200 23752
rect 8570 23740 8576 23752
rect 8628 23740 8634 23792
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9950 23780 9956 23792
rect 9171 23752 9956 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 12526 23780 12532 23792
rect 11011 23752 12532 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 15746 23780 15752 23792
rect 14323 23752 15752 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 16117 23783 16175 23789
rect 16117 23749 16129 23783
rect 16163 23780 16175 23783
rect 18322 23780 18328 23792
rect 16163 23752 18328 23780
rect 16163 23749 16175 23752
rect 16117 23743 16175 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 18969 23783 19027 23789
rect 18969 23749 18981 23783
rect 19015 23780 19027 23783
rect 19058 23780 19064 23792
rect 19015 23752 19064 23780
rect 19015 23749 19027 23752
rect 18969 23743 19027 23749
rect 19058 23740 19064 23752
rect 19116 23740 19122 23792
rect 19242 23740 19248 23792
rect 19300 23780 19306 23792
rect 19300 23752 19458 23780
rect 19300 23740 19306 23752
rect 21174 23740 21180 23792
rect 21232 23740 21238 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 21836 23752 22293 23780
rect 21836 23724 21864 23752
rect 22281 23749 22293 23752
rect 22327 23749 22339 23783
rect 22281 23743 22339 23749
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 7101 23715 7159 23721
rect 7101 23712 7113 23715
rect 6604 23684 7113 23712
rect 6604 23672 6610 23684
rect 7101 23681 7113 23684
rect 7147 23681 7159 23715
rect 7101 23675 7159 23681
rect 7193 23715 7251 23721
rect 7193 23681 7205 23715
rect 7239 23712 7251 23715
rect 7742 23712 7748 23724
rect 7239 23684 7748 23712
rect 7239 23681 7251 23684
rect 7193 23675 7251 23681
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23712 9919 23715
rect 11146 23712 11152 23724
rect 9907 23684 11152 23712
rect 9907 23681 9919 23684
rect 9861 23675 9919 23681
rect 11146 23672 11152 23684
rect 11204 23672 11210 23724
rect 13262 23672 13268 23724
rect 13320 23672 13326 23724
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23712 15163 23715
rect 16574 23712 16580 23724
rect 15151 23684 16580 23712
rect 15151 23681 15163 23684
rect 15105 23675 15163 23681
rect 16574 23672 16580 23684
rect 16632 23672 16638 23724
rect 16942 23672 16948 23724
rect 17000 23672 17006 23724
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 18414 23712 18420 23724
rect 17184 23684 18420 23712
rect 17184 23672 17190 23684
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 18690 23672 18696 23724
rect 18748 23672 18754 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 20772 23684 21005 23712
rect 20772 23672 20778 23684
rect 20993 23681 21005 23684
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 21818 23672 21824 23724
rect 21876 23672 21882 23724
rect 23400 23698 23428 23820
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24213 23851 24271 23857
rect 24213 23817 24225 23851
rect 24259 23848 24271 23851
rect 24946 23848 24952 23860
rect 24259 23820 24952 23848
rect 24259 23817 24271 23820
rect 24213 23811 24271 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25774 23808 25780 23860
rect 25832 23848 25838 23860
rect 29365 23851 29423 23857
rect 29365 23848 29377 23851
rect 25832 23820 29377 23848
rect 25832 23808 25838 23820
rect 29365 23817 29377 23820
rect 29411 23817 29423 23851
rect 29365 23811 29423 23817
rect 30190 23808 30196 23860
rect 30248 23808 30254 23860
rect 31018 23808 31024 23860
rect 31076 23848 31082 23860
rect 36081 23851 36139 23857
rect 36081 23848 36093 23851
rect 31076 23820 36093 23848
rect 31076 23808 31082 23820
rect 36081 23817 36093 23820
rect 36127 23817 36139 23851
rect 36081 23811 36139 23817
rect 38470 23808 38476 23860
rect 38528 23808 38534 23860
rect 39025 23851 39083 23857
rect 39025 23817 39037 23851
rect 39071 23848 39083 23851
rect 39206 23848 39212 23860
rect 39071 23820 39212 23848
rect 39071 23817 39083 23820
rect 39025 23811 39083 23817
rect 39206 23808 39212 23820
rect 39264 23808 39270 23860
rect 39574 23808 39580 23860
rect 39632 23848 39638 23860
rect 39853 23851 39911 23857
rect 39853 23848 39865 23851
rect 39632 23820 39865 23848
rect 39632 23808 39638 23820
rect 39853 23817 39865 23820
rect 39899 23817 39911 23851
rect 39853 23811 39911 23817
rect 40310 23808 40316 23860
rect 40368 23808 40374 23860
rect 41506 23808 41512 23860
rect 41564 23848 41570 23860
rect 42153 23851 42211 23857
rect 42153 23848 42165 23851
rect 41564 23820 42165 23848
rect 41564 23808 41570 23820
rect 42153 23817 42165 23820
rect 42199 23817 42211 23851
rect 42153 23811 42211 23817
rect 43254 23808 43260 23860
rect 43312 23808 43318 23860
rect 45554 23808 45560 23860
rect 45612 23848 45618 23860
rect 45741 23851 45799 23857
rect 45741 23848 45753 23851
rect 45612 23820 45753 23848
rect 45612 23808 45618 23820
rect 45741 23817 45753 23820
rect 45787 23817 45799 23851
rect 45741 23811 45799 23817
rect 47302 23808 47308 23860
rect 47360 23848 47366 23860
rect 47581 23851 47639 23857
rect 47581 23848 47593 23851
rect 47360 23820 47593 23848
rect 47360 23808 47366 23820
rect 47581 23817 47593 23820
rect 47627 23817 47639 23851
rect 47581 23811 47639 23817
rect 47854 23808 47860 23860
rect 47912 23808 47918 23860
rect 25406 23780 25412 23792
rect 23584 23752 25412 23780
rect 4120 23616 4200 23644
rect 4120 23604 4126 23616
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6457 23647 6515 23653
rect 6457 23613 6469 23647
rect 6503 23644 6515 23647
rect 6503 23616 7328 23644
rect 6503 23613 6515 23616
rect 6457 23607 6515 23613
rect 1210 23536 1216 23588
rect 1268 23576 1274 23588
rect 6733 23579 6791 23585
rect 6733 23576 6745 23579
rect 1268 23548 2360 23576
rect 1268 23536 1274 23548
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 2225 23511 2283 23517
rect 2225 23508 2237 23511
rect 1820 23480 2237 23508
rect 1820 23468 1826 23480
rect 2225 23477 2237 23480
rect 2271 23477 2283 23511
rect 2332 23508 2360 23548
rect 2746 23548 6745 23576
rect 2746 23508 2774 23548
rect 6733 23545 6745 23548
rect 6779 23545 6791 23579
rect 7300 23576 7328 23616
rect 7374 23604 7380 23656
rect 7432 23604 7438 23656
rect 7466 23604 7472 23656
rect 7524 23644 7530 23656
rect 12529 23647 12587 23653
rect 7524 23616 11928 23644
rect 7524 23604 7530 23616
rect 11330 23576 11336 23588
rect 7300 23548 11336 23576
rect 6733 23539 6791 23545
rect 11330 23536 11336 23548
rect 11388 23536 11394 23588
rect 11900 23585 11928 23616
rect 12529 23613 12541 23647
rect 12575 23644 12587 23647
rect 17402 23644 17408 23656
rect 12575 23616 17408 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 17402 23604 17408 23616
rect 17460 23604 17466 23656
rect 17862 23604 17868 23656
rect 17920 23604 17926 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 20088 23616 22017 23644
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23545 11943 23579
rect 11885 23539 11943 23545
rect 16758 23536 16764 23588
rect 16816 23576 16822 23588
rect 17586 23576 17592 23588
rect 16816 23548 17592 23576
rect 16816 23536 16822 23548
rect 17586 23536 17592 23548
rect 17644 23536 17650 23588
rect 20088 23520 20116 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22370 23604 22376 23656
rect 22428 23644 22434 23656
rect 23584 23644 23612 23752
rect 25406 23740 25412 23752
rect 25464 23740 25470 23792
rect 26418 23780 26424 23792
rect 26358 23752 26424 23780
rect 26418 23740 26424 23752
rect 26476 23740 26482 23792
rect 30098 23740 30104 23792
rect 30156 23740 30162 23792
rect 32306 23740 32312 23792
rect 32364 23740 32370 23792
rect 32858 23740 32864 23792
rect 32916 23780 32922 23792
rect 32953 23783 33011 23789
rect 32953 23780 32965 23783
rect 32916 23752 32965 23780
rect 32916 23740 32922 23752
rect 32953 23749 32965 23752
rect 32999 23749 33011 23783
rect 32953 23743 33011 23749
rect 33594 23740 33600 23792
rect 33652 23780 33658 23792
rect 34149 23783 34207 23789
rect 34149 23780 34161 23783
rect 33652 23752 34161 23780
rect 33652 23740 33658 23752
rect 34149 23749 34161 23752
rect 34195 23749 34207 23783
rect 34149 23743 34207 23749
rect 34882 23740 34888 23792
rect 34940 23740 34946 23792
rect 34974 23740 34980 23792
rect 35032 23780 35038 23792
rect 35621 23783 35679 23789
rect 35621 23780 35633 23783
rect 35032 23752 35633 23780
rect 35032 23740 35038 23752
rect 35621 23749 35633 23752
rect 35667 23749 35679 23783
rect 35621 23743 35679 23749
rect 36538 23740 36544 23792
rect 36596 23780 36602 23792
rect 38657 23783 38715 23789
rect 38657 23780 38669 23783
rect 36596 23752 38669 23780
rect 36596 23740 36602 23752
rect 38657 23749 38669 23752
rect 38703 23749 38715 23783
rect 38657 23743 38715 23749
rect 28534 23672 28540 23724
rect 28592 23672 28598 23724
rect 29549 23715 29607 23721
rect 29549 23681 29561 23715
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 24857 23647 24915 23653
rect 24857 23644 24869 23647
rect 22428 23616 23612 23644
rect 23676 23616 24869 23644
rect 22428 23604 22434 23616
rect 2332 23480 2774 23508
rect 2225 23471 2283 23477
rect 3878 23468 3884 23520
rect 3936 23508 3942 23520
rect 4982 23508 4988 23520
rect 3936 23480 4988 23508
rect 3936 23468 3942 23480
rect 4982 23468 4988 23480
rect 5040 23468 5046 23520
rect 6546 23468 6552 23520
rect 6604 23468 6610 23520
rect 11422 23468 11428 23520
rect 11480 23508 11486 23520
rect 11517 23511 11575 23517
rect 11517 23508 11529 23511
rect 11480 23480 11529 23508
rect 11480 23468 11486 23480
rect 11517 23477 11529 23480
rect 11563 23508 11575 23511
rect 12250 23508 12256 23520
rect 11563 23480 12256 23508
rect 11563 23477 11575 23480
rect 11517 23471 11575 23477
rect 12250 23468 12256 23480
rect 12308 23508 12314 23520
rect 12802 23508 12808 23520
rect 12308 23480 12808 23508
rect 12308 23468 12314 23480
rect 12802 23468 12808 23480
rect 12860 23468 12866 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 20070 23508 20076 23520
rect 18748 23480 20076 23508
rect 18748 23468 18754 23480
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20441 23511 20499 23517
rect 20441 23477 20453 23511
rect 20487 23508 20499 23511
rect 20622 23508 20628 23520
rect 20487 23480 20628 23508
rect 20487 23477 20499 23480
rect 20441 23471 20499 23477
rect 20622 23468 20628 23480
rect 20680 23468 20686 23520
rect 21637 23511 21695 23517
rect 21637 23477 21649 23511
rect 21683 23508 21695 23511
rect 22094 23508 22100 23520
rect 21683 23480 22100 23508
rect 21683 23477 21695 23480
rect 21637 23471 21695 23477
rect 22094 23468 22100 23480
rect 22152 23468 22158 23520
rect 22830 23468 22836 23520
rect 22888 23508 22894 23520
rect 23676 23508 23704 23616
rect 24857 23613 24869 23616
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23644 25191 23647
rect 26142 23644 26148 23656
rect 25179 23616 26148 23644
rect 25179 23613 25191 23616
rect 25133 23607 25191 23613
rect 22888 23480 23704 23508
rect 22888 23468 22894 23480
rect 23750 23468 23756 23520
rect 23808 23468 23814 23520
rect 24872 23508 24900 23607
rect 26142 23604 26148 23616
rect 26200 23604 26206 23656
rect 27154 23644 27160 23656
rect 26252 23616 27160 23644
rect 26252 23508 26280 23616
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 27433 23647 27491 23653
rect 27433 23644 27445 23647
rect 27264 23616 27445 23644
rect 27264 23576 27292 23616
rect 27433 23613 27445 23616
rect 27479 23613 27491 23647
rect 27433 23607 27491 23613
rect 27522 23604 27528 23656
rect 27580 23644 27586 23656
rect 29564 23644 29592 23675
rect 30374 23672 30380 23724
rect 30432 23712 30438 23724
rect 31386 23712 31392 23724
rect 30432 23684 31392 23712
rect 30432 23672 30438 23684
rect 31386 23672 31392 23684
rect 31444 23712 31450 23724
rect 31481 23715 31539 23721
rect 31481 23712 31493 23715
rect 31444 23684 31493 23712
rect 31444 23672 31450 23684
rect 31481 23681 31493 23684
rect 31527 23681 31539 23715
rect 33413 23715 33471 23721
rect 33413 23712 33425 23715
rect 31481 23675 31539 23681
rect 31726 23684 33425 23712
rect 31726 23644 31754 23684
rect 33413 23681 33425 23684
rect 33459 23681 33471 23715
rect 33413 23675 33471 23681
rect 33965 23715 34023 23721
rect 33965 23681 33977 23715
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 27580 23616 31754 23644
rect 27580 23604 27586 23616
rect 32122 23604 32128 23656
rect 32180 23644 32186 23656
rect 33980 23644 34008 23675
rect 34698 23672 34704 23724
rect 34756 23672 34762 23724
rect 35437 23715 35495 23721
rect 35437 23681 35449 23715
rect 35483 23681 35495 23715
rect 35437 23675 35495 23681
rect 35452 23644 35480 23675
rect 36262 23672 36268 23724
rect 36320 23672 36326 23724
rect 36354 23672 36360 23724
rect 36412 23712 36418 23724
rect 36909 23715 36967 23721
rect 36909 23712 36921 23715
rect 36412 23684 36921 23712
rect 36412 23672 36418 23684
rect 36909 23681 36921 23684
rect 36955 23712 36967 23715
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 36955 23684 37289 23712
rect 36955 23681 36967 23684
rect 36909 23675 36967 23681
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 37277 23675 37335 23681
rect 37642 23672 37648 23724
rect 37700 23712 37706 23724
rect 37921 23715 37979 23721
rect 37921 23712 37933 23715
rect 37700 23684 37933 23712
rect 37700 23672 37706 23684
rect 37921 23681 37933 23684
rect 37967 23712 37979 23715
rect 38197 23715 38255 23721
rect 38197 23712 38209 23715
rect 37967 23684 38209 23712
rect 37967 23681 37979 23684
rect 37921 23675 37979 23681
rect 38197 23681 38209 23684
rect 38243 23681 38255 23715
rect 40328 23712 40356 23808
rect 47872 23780 47900 23808
rect 47872 23752 49096 23780
rect 40865 23715 40923 23721
rect 40865 23712 40877 23715
rect 40328 23684 40877 23712
rect 38197 23675 38255 23681
rect 40865 23681 40877 23684
rect 40911 23681 40923 23715
rect 40865 23675 40923 23681
rect 40954 23672 40960 23724
rect 41012 23712 41018 23724
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 41012 23684 41521 23712
rect 41012 23672 41018 23684
rect 41509 23681 41521 23684
rect 41555 23712 41567 23715
rect 41785 23715 41843 23721
rect 41785 23712 41797 23715
rect 41555 23684 41797 23712
rect 41555 23681 41567 23684
rect 41509 23675 41567 23681
rect 41785 23681 41797 23684
rect 41831 23681 41843 23715
rect 41785 23675 41843 23681
rect 42058 23672 42064 23724
rect 42116 23712 42122 23724
rect 42613 23715 42671 23721
rect 42613 23712 42625 23715
rect 42116 23684 42625 23712
rect 42116 23672 42122 23684
rect 42613 23681 42625 23684
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 43714 23672 43720 23724
rect 43772 23672 43778 23724
rect 44174 23672 44180 23724
rect 44232 23712 44238 23724
rect 44453 23715 44511 23721
rect 44453 23712 44465 23715
rect 44232 23684 44465 23712
rect 44232 23672 44238 23684
rect 44453 23681 44465 23684
rect 44499 23712 44511 23715
rect 45005 23715 45063 23721
rect 45005 23712 45017 23715
rect 44499 23684 45017 23712
rect 44499 23681 44511 23684
rect 44453 23675 44511 23681
rect 45005 23681 45017 23684
rect 45051 23681 45063 23715
rect 45005 23675 45063 23681
rect 46658 23672 46664 23724
rect 46716 23712 46722 23724
rect 46753 23715 46811 23721
rect 46753 23712 46765 23715
rect 46716 23684 46765 23712
rect 46716 23672 46722 23684
rect 46753 23681 46765 23684
rect 46799 23712 46811 23715
rect 47305 23715 47363 23721
rect 47305 23712 47317 23715
rect 46799 23684 47317 23712
rect 46799 23681 46811 23684
rect 46753 23675 46811 23681
rect 47305 23681 47317 23684
rect 47351 23681 47363 23715
rect 47305 23675 47363 23681
rect 48041 23715 48099 23721
rect 48041 23681 48053 23715
rect 48087 23712 48099 23715
rect 48314 23712 48320 23724
rect 48087 23684 48320 23712
rect 48087 23681 48099 23684
rect 48041 23675 48099 23681
rect 48314 23672 48320 23684
rect 48372 23672 48378 23724
rect 49068 23721 49096 23752
rect 49053 23715 49111 23721
rect 49053 23681 49065 23715
rect 49099 23681 49111 23715
rect 49053 23675 49111 23681
rect 32180 23616 34008 23644
rect 34072 23616 35480 23644
rect 36096 23616 40724 23644
rect 32180 23604 32186 23616
rect 30650 23576 30656 23588
rect 26620 23548 27292 23576
rect 28460 23548 30656 23576
rect 26620 23520 26648 23548
rect 24872 23480 26280 23508
rect 26602 23468 26608 23520
rect 26660 23468 26666 23520
rect 26786 23468 26792 23520
rect 26844 23508 26850 23520
rect 28460 23508 28488 23548
rect 30650 23536 30656 23548
rect 30708 23536 30714 23588
rect 30742 23536 30748 23588
rect 30800 23576 30806 23588
rect 30837 23579 30895 23585
rect 30837 23576 30849 23579
rect 30800 23548 30849 23576
rect 30800 23536 30806 23548
rect 30837 23545 30849 23548
rect 30883 23576 30895 23579
rect 31021 23579 31079 23585
rect 31021 23576 31033 23579
rect 30883 23548 31033 23576
rect 30883 23545 30895 23548
rect 30837 23539 30895 23545
rect 31021 23545 31033 23548
rect 31067 23576 31079 23579
rect 31662 23576 31668 23588
rect 31067 23548 31668 23576
rect 31067 23545 31079 23548
rect 31021 23539 31079 23545
rect 31662 23536 31668 23548
rect 31720 23536 31726 23588
rect 31754 23536 31760 23588
rect 31812 23536 31818 23588
rect 32582 23536 32588 23588
rect 32640 23576 32646 23588
rect 34072 23576 34100 23616
rect 32640 23548 34100 23576
rect 32640 23536 32646 23548
rect 26844 23480 28488 23508
rect 26844 23468 26850 23480
rect 28718 23468 28724 23520
rect 28776 23508 28782 23520
rect 28905 23511 28963 23517
rect 28905 23508 28917 23511
rect 28776 23480 28917 23508
rect 28776 23468 28782 23480
rect 28905 23477 28917 23480
rect 28951 23477 28963 23511
rect 28905 23471 28963 23477
rect 30558 23468 30564 23520
rect 30616 23468 30622 23520
rect 31110 23468 31116 23520
rect 31168 23508 31174 23520
rect 31297 23511 31355 23517
rect 31297 23508 31309 23511
rect 31168 23480 31309 23508
rect 31168 23468 31174 23480
rect 31297 23477 31309 23480
rect 31343 23477 31355 23511
rect 31297 23471 31355 23477
rect 33870 23468 33876 23520
rect 33928 23508 33934 23520
rect 36096 23508 36124 23616
rect 37182 23536 37188 23588
rect 37240 23576 37246 23588
rect 40696 23585 40724 23616
rect 40681 23579 40739 23585
rect 37240 23548 39160 23576
rect 37240 23536 37246 23548
rect 33928 23480 36124 23508
rect 33928 23468 33934 23480
rect 36722 23468 36728 23520
rect 36780 23468 36786 23520
rect 37734 23468 37740 23520
rect 37792 23468 37798 23520
rect 39132 23508 39160 23548
rect 40681 23545 40693 23579
rect 40727 23545 40739 23579
rect 40681 23539 40739 23545
rect 40770 23536 40776 23588
rect 40828 23576 40834 23588
rect 49237 23579 49295 23585
rect 49237 23576 49249 23579
rect 40828 23548 49249 23576
rect 40828 23536 40834 23548
rect 49237 23545 49249 23548
rect 49283 23545 49295 23579
rect 49237 23539 49295 23545
rect 41325 23511 41383 23517
rect 41325 23508 41337 23511
rect 39132 23480 41337 23508
rect 41325 23477 41337 23480
rect 41371 23477 41383 23511
rect 41325 23471 41383 23477
rect 41414 23468 41420 23520
rect 41472 23508 41478 23520
rect 43901 23511 43959 23517
rect 43901 23508 43913 23511
rect 41472 23480 43913 23508
rect 41472 23468 41478 23480
rect 43901 23477 43913 23480
rect 43947 23477 43959 23511
rect 43901 23471 43959 23477
rect 44634 23468 44640 23520
rect 44692 23468 44698 23520
rect 46934 23468 46940 23520
rect 46992 23468 46998 23520
rect 48498 23468 48504 23520
rect 48556 23468 48562 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 3694 23264 3700 23316
rect 3752 23304 3758 23316
rect 3789 23307 3847 23313
rect 3789 23304 3801 23307
rect 3752 23276 3801 23304
rect 3752 23264 3758 23276
rect 3789 23273 3801 23276
rect 3835 23304 3847 23307
rect 3878 23304 3884 23316
rect 3835 23276 3884 23304
rect 3835 23273 3847 23276
rect 3789 23267 3847 23273
rect 3878 23264 3884 23276
rect 3936 23264 3942 23316
rect 3970 23264 3976 23316
rect 4028 23264 4034 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 4080 23276 14473 23304
rect 3418 23196 3424 23248
rect 3476 23236 3482 23248
rect 4080 23236 4108 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 24118 23304 24124 23316
rect 18012 23276 24124 23304
rect 18012 23264 18018 23276
rect 24118 23264 24124 23276
rect 24176 23264 24182 23316
rect 24394 23264 24400 23316
rect 24452 23304 24458 23316
rect 26602 23304 26608 23316
rect 24452 23276 26608 23304
rect 24452 23264 24458 23276
rect 26602 23264 26608 23276
rect 26660 23264 26666 23316
rect 27062 23304 27068 23316
rect 26896 23276 27068 23304
rect 6638 23236 6644 23248
rect 3476 23208 4108 23236
rect 4632 23208 6644 23236
rect 3476 23196 3482 23208
rect 3605 23171 3663 23177
rect 3605 23137 3617 23171
rect 3651 23168 3663 23171
rect 3786 23168 3792 23180
rect 3651 23140 3792 23168
rect 3651 23137 3663 23140
rect 3605 23131 3663 23137
rect 3786 23128 3792 23140
rect 3844 23128 3850 23180
rect 4632 23168 4660 23208
rect 6638 23196 6644 23208
rect 6696 23196 6702 23248
rect 12802 23196 12808 23248
rect 12860 23236 12866 23248
rect 13633 23239 13691 23245
rect 13633 23236 13645 23239
rect 12860 23208 13645 23236
rect 12860 23196 12866 23208
rect 13633 23205 13645 23208
rect 13679 23236 13691 23239
rect 14921 23239 14979 23245
rect 14921 23236 14933 23239
rect 13679 23208 14933 23236
rect 13679 23205 13691 23208
rect 13633 23199 13691 23205
rect 14921 23205 14933 23208
rect 14967 23205 14979 23239
rect 14921 23199 14979 23205
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 19058 23236 19064 23248
rect 18923 23208 19064 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 19058 23196 19064 23208
rect 19116 23196 19122 23248
rect 19426 23196 19432 23248
rect 19484 23196 19490 23248
rect 19610 23196 19616 23248
rect 19668 23196 19674 23248
rect 23750 23196 23756 23248
rect 23808 23236 23814 23248
rect 23808 23208 25268 23236
rect 23808 23196 23814 23208
rect 3988 23140 4660 23168
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 1811 23072 3372 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 3344 22964 3372 23072
rect 3421 23035 3479 23041
rect 3421 23001 3433 23035
rect 3467 23032 3479 23035
rect 3988 23032 4016 23140
rect 4706 23128 4712 23180
rect 4764 23128 4770 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 9030 23128 9036 23180
rect 9088 23168 9094 23180
rect 11422 23168 11428 23180
rect 9088 23140 11428 23168
rect 9088 23128 9094 23140
rect 3467 23004 4016 23032
rect 4080 23072 5304 23100
rect 3467 23001 3479 23004
rect 3421 22995 3479 23001
rect 4080 22964 4108 23072
rect 4246 22992 4252 23044
rect 4304 23032 4310 23044
rect 4525 23035 4583 23041
rect 4525 23032 4537 23035
rect 4304 23004 4537 23032
rect 4304 22992 4310 23004
rect 4525 23001 4537 23004
rect 4571 23032 4583 23035
rect 5166 23032 5172 23044
rect 4571 23004 5172 23032
rect 4571 23001 4583 23004
rect 4525 22995 4583 23001
rect 5166 22992 5172 23004
rect 5224 22992 5230 23044
rect 5276 23032 5304 23072
rect 5350 23060 5356 23112
rect 5408 23060 5414 23112
rect 7190 23060 7196 23112
rect 7248 23060 7254 23112
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 8904 23072 9321 23100
rect 8904 23060 8910 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 10704 23086 10732 23140
rect 11422 23128 11428 23140
rect 11480 23128 11486 23180
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 12434 23168 12440 23180
rect 11563 23140 12440 23168
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 12526 23128 12532 23180
rect 12584 23168 12590 23180
rect 13909 23171 13967 23177
rect 12584 23140 13032 23168
rect 12584 23128 12590 23140
rect 13004 23100 13032 23140
rect 13909 23137 13921 23171
rect 13955 23168 13967 23171
rect 17770 23168 17776 23180
rect 13955 23140 17776 23168
rect 13955 23137 13967 23140
rect 13909 23131 13967 23137
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 17862 23128 17868 23180
rect 17920 23168 17926 23180
rect 19628 23168 19656 23196
rect 17920 23140 19656 23168
rect 17920 23128 17926 23140
rect 20070 23128 20076 23180
rect 20128 23128 20134 23180
rect 22557 23171 22615 23177
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 23768 23168 23796 23196
rect 22603 23140 23796 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 25240 23168 25268 23208
rect 26142 23196 26148 23248
rect 26200 23236 26206 23248
rect 26896 23236 26924 23276
rect 27062 23264 27068 23276
rect 27120 23264 27126 23316
rect 27338 23264 27344 23316
rect 27396 23264 27402 23316
rect 27512 23307 27570 23313
rect 27512 23273 27524 23307
rect 27558 23304 27570 23307
rect 28718 23304 28724 23316
rect 27558 23276 28724 23304
rect 27558 23273 27570 23276
rect 27512 23267 27570 23273
rect 28718 23264 28724 23276
rect 28776 23264 28782 23316
rect 28994 23264 29000 23316
rect 29052 23304 29058 23316
rect 29990 23307 30048 23313
rect 29990 23304 30002 23307
rect 29052 23276 30002 23304
rect 29052 23264 29058 23276
rect 29990 23273 30002 23276
rect 30036 23273 30048 23307
rect 29990 23267 30048 23273
rect 30558 23264 30564 23316
rect 30616 23304 30622 23316
rect 30616 23276 31754 23304
rect 30616 23264 30622 23276
rect 27356 23236 27384 23264
rect 26200 23208 26924 23236
rect 26988 23208 27384 23236
rect 31726 23236 31754 23276
rect 31846 23264 31852 23316
rect 31904 23304 31910 23316
rect 32306 23304 32312 23316
rect 31904 23276 32312 23304
rect 31904 23264 31910 23276
rect 32306 23264 32312 23276
rect 32364 23264 32370 23316
rect 32490 23264 32496 23316
rect 32548 23264 32554 23316
rect 33229 23307 33287 23313
rect 33229 23273 33241 23307
rect 33275 23304 33287 23307
rect 33502 23304 33508 23316
rect 33275 23276 33508 23304
rect 33275 23273 33287 23276
rect 33229 23267 33287 23273
rect 33502 23264 33508 23276
rect 33560 23264 33566 23316
rect 33962 23264 33968 23316
rect 34020 23264 34026 23316
rect 34422 23264 34428 23316
rect 34480 23304 34486 23316
rect 34480 23276 35388 23304
rect 34480 23264 34486 23276
rect 35066 23236 35072 23248
rect 31726 23208 35072 23236
rect 26200 23196 26206 23208
rect 26329 23171 26387 23177
rect 26329 23168 26341 23171
rect 25240 23140 26341 23168
rect 26329 23137 26341 23140
rect 26375 23137 26387 23171
rect 26329 23131 26387 23137
rect 15473 23103 15531 23109
rect 13004 23072 14412 23100
rect 9309 23063 9367 23069
rect 14384 23044 14412 23072
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 16666 23100 16672 23112
rect 15519 23072 16672 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 16908 23072 17141 23100
rect 16908 23060 16914 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 7558 23032 7564 23044
rect 5276 23004 7564 23032
rect 7558 22992 7564 23004
rect 7616 22992 7622 23044
rect 8478 22992 8484 23044
rect 8536 23032 8542 23044
rect 8536 23004 9536 23032
rect 8536 22992 8542 23004
rect 3344 22936 4108 22964
rect 4154 22924 4160 22976
rect 4212 22924 4218 22976
rect 4617 22967 4675 22973
rect 4617 22933 4629 22967
rect 4663 22964 4675 22967
rect 7466 22964 7472 22976
rect 4663 22936 7472 22964
rect 4663 22933 4675 22936
rect 4617 22927 4675 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 9030 22924 9036 22976
rect 9088 22924 9094 22976
rect 9508 22964 9536 23004
rect 9582 22992 9588 23044
rect 9640 22992 9646 23044
rect 11793 23035 11851 23041
rect 11793 23032 11805 23035
rect 11256 23004 11805 23032
rect 11057 22967 11115 22973
rect 11057 22964 11069 22967
rect 9508 22936 11069 22964
rect 11057 22933 11069 22936
rect 11103 22964 11115 22967
rect 11256 22964 11284 23004
rect 11793 23001 11805 23004
rect 11839 23001 11851 23035
rect 11793 22995 11851 23001
rect 12250 22992 12256 23044
rect 12308 22992 12314 23044
rect 14366 22992 14372 23044
rect 14424 22992 14430 23044
rect 16485 23035 16543 23041
rect 16485 23001 16497 23035
rect 16531 23001 16543 23035
rect 16485 22995 16543 23001
rect 11103 22936 11284 22964
rect 11103 22933 11115 22936
rect 11057 22927 11115 22933
rect 11330 22924 11336 22976
rect 11388 22964 11394 22976
rect 12526 22964 12532 22976
rect 11388 22936 12532 22964
rect 11388 22924 11394 22936
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 12710 22924 12716 22976
rect 12768 22964 12774 22976
rect 13265 22967 13323 22973
rect 13265 22964 13277 22967
rect 12768 22936 13277 22964
rect 12768 22924 12774 22936
rect 13265 22933 13277 22936
rect 13311 22964 13323 22967
rect 13538 22964 13544 22976
rect 13311 22936 13544 22964
rect 13311 22933 13323 22936
rect 13265 22927 13323 22933
rect 13538 22924 13544 22936
rect 13596 22924 13602 22976
rect 16500 22964 16528 22995
rect 17402 22992 17408 23044
rect 17460 22992 17466 23044
rect 17494 22992 17500 23044
rect 17552 23032 17558 23044
rect 17552 23004 17894 23032
rect 17552 22992 17558 23004
rect 17678 22964 17684 22976
rect 16500 22936 17684 22964
rect 17678 22924 17684 22936
rect 17736 22924 17742 22976
rect 19628 22964 19656 23063
rect 22278 23060 22284 23112
rect 22336 23060 22342 23112
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23100 25099 23103
rect 26988 23100 27016 23208
rect 35066 23196 35072 23208
rect 35124 23196 35130 23248
rect 27154 23128 27160 23180
rect 27212 23168 27218 23180
rect 27249 23171 27307 23177
rect 27249 23168 27261 23171
rect 27212 23140 27261 23168
rect 27212 23128 27218 23140
rect 27249 23137 27261 23140
rect 27295 23168 27307 23171
rect 27614 23168 27620 23180
rect 27295 23140 27620 23168
rect 27295 23137 27307 23140
rect 27249 23131 27307 23137
rect 27614 23128 27620 23140
rect 27672 23168 27678 23180
rect 29733 23171 29791 23177
rect 29733 23168 29745 23171
rect 27672 23140 29745 23168
rect 27672 23128 27678 23140
rect 29733 23137 29745 23140
rect 29779 23168 29791 23171
rect 30742 23168 30748 23180
rect 29779 23140 30748 23168
rect 29779 23137 29791 23140
rect 29733 23131 29791 23137
rect 30742 23128 30748 23140
rect 30800 23128 30806 23180
rect 35360 23168 35388 23276
rect 36814 23264 36820 23316
rect 36872 23264 36878 23316
rect 37274 23264 37280 23316
rect 37332 23264 37338 23316
rect 43625 23307 43683 23313
rect 43625 23273 43637 23307
rect 43671 23304 43683 23307
rect 43714 23304 43720 23316
rect 43671 23276 43720 23304
rect 43671 23273 43683 23276
rect 43625 23267 43683 23273
rect 43714 23264 43720 23276
rect 43772 23264 43778 23316
rect 35618 23196 35624 23248
rect 35676 23236 35682 23248
rect 37001 23239 37059 23245
rect 37001 23236 37013 23239
rect 35676 23208 37013 23236
rect 35676 23196 35682 23208
rect 37001 23205 37013 23208
rect 37047 23205 37059 23239
rect 48409 23239 48467 23245
rect 48409 23236 48421 23239
rect 37001 23199 37059 23205
rect 45526 23208 48421 23236
rect 31956 23140 35112 23168
rect 35360 23140 39988 23168
rect 25087 23072 27016 23100
rect 25087 23069 25099 23072
rect 25041 23063 25099 23069
rect 28534 23060 28540 23112
rect 28592 23100 28598 23112
rect 31846 23100 31852 23112
rect 28592 23086 28658 23100
rect 28592 23072 28672 23086
rect 31142 23072 31852 23100
rect 28592 23060 28598 23072
rect 20346 22992 20352 23044
rect 20404 22992 20410 23044
rect 22094 23032 22100 23044
rect 21574 23004 22100 23032
rect 22094 22992 22100 23004
rect 22152 22992 22158 23044
rect 23842 23032 23848 23044
rect 23782 23004 23848 23032
rect 23842 22992 23848 23004
rect 23900 23032 23906 23044
rect 24486 23032 24492 23044
rect 23900 23004 24492 23032
rect 23900 22992 23906 23004
rect 24486 22992 24492 23004
rect 24544 22992 24550 23044
rect 26237 23035 26295 23041
rect 26237 23001 26249 23035
rect 26283 23032 26295 23035
rect 26283 23004 27292 23032
rect 26283 23001 26295 23004
rect 26237 22995 26295 23001
rect 20530 22964 20536 22976
rect 19628 22936 20536 22964
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 21818 22924 21824 22976
rect 21876 22924 21882 22976
rect 23198 22924 23204 22976
rect 23256 22964 23262 22976
rect 24029 22967 24087 22973
rect 24029 22964 24041 22967
rect 23256 22936 24041 22964
rect 23256 22924 23262 22936
rect 24029 22933 24041 22936
rect 24075 22933 24087 22967
rect 24029 22927 24087 22933
rect 24118 22924 24124 22976
rect 24176 22964 24182 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 24176 22936 24593 22964
rect 24176 22924 24182 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 24946 22924 24952 22976
rect 25004 22924 25010 22976
rect 25406 22924 25412 22976
rect 25464 22964 25470 22976
rect 25777 22967 25835 22973
rect 25777 22964 25789 22967
rect 25464 22936 25789 22964
rect 25464 22924 25470 22936
rect 25777 22933 25789 22936
rect 25823 22933 25835 22967
rect 25777 22927 25835 22933
rect 26050 22924 26056 22976
rect 26108 22964 26114 22976
rect 26145 22967 26203 22973
rect 26145 22964 26157 22967
rect 26108 22936 26157 22964
rect 26108 22924 26114 22936
rect 26145 22933 26157 22936
rect 26191 22964 26203 22967
rect 26510 22964 26516 22976
rect 26191 22936 26516 22964
rect 26191 22933 26203 22936
rect 26145 22927 26203 22933
rect 26510 22924 26516 22936
rect 26568 22924 26574 22976
rect 26786 22924 26792 22976
rect 26844 22924 26850 22976
rect 27264 22964 27292 23004
rect 28350 22964 28356 22976
rect 27264 22936 28356 22964
rect 28350 22924 28356 22936
rect 28408 22924 28414 22976
rect 28644 22964 28672 23072
rect 31846 23060 31852 23072
rect 31904 23060 31910 23112
rect 28810 22992 28816 23044
rect 28868 23032 28874 23044
rect 31956 23032 31984 23140
rect 32030 23060 32036 23112
rect 32088 23100 32094 23112
rect 33873 23103 33931 23109
rect 33873 23100 33885 23103
rect 32088 23072 33885 23100
rect 32088 23060 32094 23072
rect 33873 23069 33885 23072
rect 33919 23069 33931 23103
rect 33873 23063 33931 23069
rect 34974 23060 34980 23112
rect 35032 23100 35038 23112
rect 35084 23109 35112 23140
rect 35069 23103 35127 23109
rect 35069 23100 35081 23103
rect 35032 23072 35081 23100
rect 35032 23060 35038 23072
rect 35069 23069 35081 23072
rect 35115 23069 35127 23103
rect 35069 23063 35127 23069
rect 35710 23060 35716 23112
rect 35768 23060 35774 23112
rect 28868 23004 30420 23032
rect 28868 22992 28874 23004
rect 28902 22964 28908 22976
rect 28644 22936 28908 22964
rect 28902 22924 28908 22936
rect 28960 22964 28966 22976
rect 29178 22964 29184 22976
rect 28960 22936 29184 22964
rect 28960 22924 28966 22936
rect 29178 22924 29184 22936
rect 29236 22964 29242 22976
rect 29273 22967 29331 22973
rect 29273 22964 29285 22967
rect 29236 22936 29285 22964
rect 29236 22924 29242 22936
rect 29273 22933 29285 22936
rect 29319 22933 29331 22967
rect 30392 22964 30420 23004
rect 31312 23004 31984 23032
rect 32401 23035 32459 23041
rect 31312 22964 31340 23004
rect 32401 23001 32413 23035
rect 32447 23032 32459 23035
rect 32858 23032 32864 23044
rect 32447 23004 32864 23032
rect 32447 23001 32459 23004
rect 32401 22995 32459 23001
rect 32858 22992 32864 23004
rect 32916 22992 32922 23044
rect 33137 23035 33195 23041
rect 33137 23001 33149 23035
rect 33183 23032 33195 23035
rect 33318 23032 33324 23044
rect 33183 23004 33324 23032
rect 33183 23001 33195 23004
rect 33137 22995 33195 23001
rect 33318 22992 33324 23004
rect 33376 22992 33382 23044
rect 36262 23032 36268 23044
rect 33888 23004 36268 23032
rect 30392 22936 31340 22964
rect 29273 22927 29331 22933
rect 31478 22924 31484 22976
rect 31536 22924 31542 22976
rect 31938 22924 31944 22976
rect 31996 22924 32002 22976
rect 32490 22924 32496 22976
rect 32548 22964 32554 22976
rect 33888 22964 33916 23004
rect 36262 22992 36268 23004
rect 36320 23032 36326 23044
rect 36633 23035 36691 23041
rect 36633 23032 36645 23035
rect 36320 23004 36645 23032
rect 36320 22992 36326 23004
rect 36633 23001 36645 23004
rect 36679 23001 36691 23035
rect 36633 22995 36691 23001
rect 39960 22976 39988 23140
rect 41141 23103 41199 23109
rect 41141 23069 41153 23103
rect 41187 23100 41199 23103
rect 42610 23100 42616 23112
rect 41187 23072 42616 23100
rect 41187 23069 41199 23072
rect 41141 23063 41199 23069
rect 42610 23060 42616 23072
rect 42668 23060 42674 23112
rect 43901 23103 43959 23109
rect 43901 23069 43913 23103
rect 43947 23100 43959 23103
rect 45526 23100 45554 23208
rect 48409 23205 48421 23208
rect 48455 23205 48467 23239
rect 48409 23199 48467 23205
rect 43947 23072 45554 23100
rect 48593 23103 48651 23109
rect 43947 23069 43959 23072
rect 43901 23063 43959 23069
rect 48593 23069 48605 23103
rect 48639 23100 48651 23103
rect 48682 23100 48688 23112
rect 48639 23072 48688 23100
rect 48639 23069 48651 23072
rect 48593 23063 48651 23069
rect 48682 23060 48688 23072
rect 48740 23060 48746 23112
rect 49050 23060 49056 23112
rect 49108 23060 49114 23112
rect 48133 23035 48191 23041
rect 48133 23001 48145 23035
rect 48179 23032 48191 23035
rect 49068 23032 49096 23060
rect 48179 23004 49096 23032
rect 48179 23001 48191 23004
rect 48133 22995 48191 23001
rect 32548 22936 33916 22964
rect 32548 22924 32554 22936
rect 34882 22924 34888 22976
rect 34940 22924 34946 22976
rect 35066 22924 35072 22976
rect 35124 22964 35130 22976
rect 35529 22967 35587 22973
rect 35529 22964 35541 22967
rect 35124 22936 35541 22964
rect 35124 22924 35130 22936
rect 35529 22933 35541 22936
rect 35575 22933 35587 22967
rect 35529 22927 35587 22933
rect 36170 22924 36176 22976
rect 36228 22924 36234 22976
rect 39942 22924 39948 22976
rect 40000 22964 40006 22976
rect 42429 22967 42487 22973
rect 42429 22964 42441 22967
rect 40000 22936 42441 22964
rect 40000 22924 40006 22936
rect 42429 22933 42441 22936
rect 42475 22933 42487 22967
rect 42429 22927 42487 22933
rect 44542 22924 44548 22976
rect 44600 22924 44606 22976
rect 47210 22924 47216 22976
rect 47268 22964 47274 22976
rect 49237 22967 49295 22973
rect 49237 22964 49249 22967
rect 47268 22936 49249 22964
rect 47268 22924 47274 22936
rect 49237 22933 49249 22936
rect 49283 22933 49295 22967
rect 49237 22927 49295 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 1026 22720 1032 22772
rect 1084 22760 1090 22772
rect 5350 22760 5356 22772
rect 1084 22732 5356 22760
rect 1084 22720 1090 22732
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 7558 22720 7564 22772
rect 7616 22760 7622 22772
rect 7616 22732 10824 22760
rect 7616 22720 7622 22732
rect 10686 22652 10692 22704
rect 10744 22652 10750 22704
rect 10796 22692 10824 22732
rect 11882 22720 11888 22772
rect 11940 22760 11946 22772
rect 12526 22760 12532 22772
rect 11940 22732 12532 22760
rect 11940 22720 11946 22732
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 14553 22763 14611 22769
rect 14553 22760 14565 22763
rect 13096 22732 14565 22760
rect 12618 22692 12624 22704
rect 10796 22664 12624 22692
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 12710 22652 12716 22704
rect 12768 22652 12774 22704
rect 12802 22652 12808 22704
rect 12860 22692 12866 22704
rect 13096 22692 13124 22732
rect 14553 22729 14565 22732
rect 14599 22729 14611 22763
rect 14553 22723 14611 22729
rect 18506 22720 18512 22772
rect 18564 22760 18570 22772
rect 18564 22732 20208 22760
rect 18564 22720 18570 22732
rect 12860 22664 13202 22692
rect 12860 22652 12866 22664
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 16666 22652 16672 22704
rect 16724 22692 16730 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16724 22664 17141 22692
rect 16724 22652 16730 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 17129 22655 17187 22661
rect 17678 22652 17684 22704
rect 17736 22652 17742 22704
rect 20070 22692 20076 22704
rect 19720 22664 20076 22692
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 3418 22624 3424 22636
rect 1811 22596 3424 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 3418 22584 3424 22596
rect 3476 22584 3482 22636
rect 3786 22584 3792 22636
rect 3844 22584 3850 22636
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 6638 22584 6644 22636
rect 6696 22624 6702 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 6696 22596 7113 22624
rect 6696 22584 6702 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22624 7251 22627
rect 7834 22624 7840 22636
rect 7239 22596 7840 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 7929 22627 7987 22633
rect 7929 22593 7941 22627
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3881 22559 3939 22565
rect 3881 22525 3893 22559
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22525 4123 22559
rect 4065 22519 4123 22525
rect 2590 22380 2596 22432
rect 2648 22420 2654 22432
rect 3421 22423 3479 22429
rect 3421 22420 3433 22423
rect 2648 22392 3433 22420
rect 2648 22380 2654 22392
rect 3421 22389 3433 22392
rect 3467 22389 3479 22423
rect 3896 22420 3924 22519
rect 4080 22488 4108 22519
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 7377 22559 7435 22565
rect 7377 22525 7389 22559
rect 7423 22556 7435 22559
rect 7650 22556 7656 22568
rect 7423 22528 7656 22556
rect 7423 22525 7435 22528
rect 7377 22519 7435 22525
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 4614 22488 4620 22500
rect 4080 22460 4620 22488
rect 4614 22448 4620 22460
rect 4672 22448 4678 22500
rect 7098 22448 7104 22500
rect 7156 22488 7162 22500
rect 7944 22488 7972 22587
rect 8202 22584 8208 22636
rect 8260 22624 8266 22636
rect 9953 22627 10011 22633
rect 9953 22624 9965 22627
rect 8260 22596 9965 22624
rect 8260 22584 8266 22596
rect 9953 22593 9965 22596
rect 9999 22624 10011 22627
rect 10042 22624 10048 22636
rect 9999 22596 10048 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 12342 22624 12348 22636
rect 11839 22596 12348 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 8662 22516 8668 22568
rect 8720 22516 8726 22568
rect 9858 22516 9864 22568
rect 9916 22556 9922 22568
rect 11698 22556 11704 22568
rect 9916 22528 11704 22556
rect 9916 22516 9922 22528
rect 11698 22516 11704 22528
rect 11756 22556 11762 22568
rect 11808 22556 11836 22587
rect 12342 22584 12348 22596
rect 12400 22584 12406 22636
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22624 15163 22627
rect 16758 22624 16764 22636
rect 15151 22596 16764 22624
rect 15151 22593 15163 22596
rect 15105 22587 15163 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19720 22633 19748 22664
rect 20070 22652 20076 22664
rect 20128 22652 20134 22704
rect 20180 22692 20208 22732
rect 20346 22720 20352 22772
rect 20404 22760 20410 22772
rect 21453 22763 21511 22769
rect 21453 22760 21465 22763
rect 20404 22732 21465 22760
rect 20404 22720 20410 22732
rect 21453 22729 21465 22732
rect 21499 22760 21511 22763
rect 25130 22760 25136 22772
rect 21499 22732 25136 22760
rect 21499 22729 21511 22732
rect 21453 22723 21511 22729
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 25774 22720 25780 22772
rect 25832 22720 25838 22772
rect 27157 22763 27215 22769
rect 27157 22729 27169 22763
rect 27203 22729 27215 22763
rect 27157 22723 27215 22729
rect 22465 22695 22523 22701
rect 20180 22664 20470 22692
rect 22465 22661 22477 22695
rect 22511 22692 22523 22695
rect 23658 22692 23664 22704
rect 22511 22664 23664 22692
rect 22511 22661 22523 22664
rect 22465 22655 22523 22661
rect 23658 22652 23664 22664
rect 23716 22652 23722 22704
rect 24670 22652 24676 22704
rect 24728 22692 24734 22704
rect 27172 22692 27200 22723
rect 28442 22720 28448 22772
rect 28500 22760 28506 22772
rect 30374 22760 30380 22772
rect 28500 22732 30380 22760
rect 28500 22720 28506 22732
rect 30374 22720 30380 22732
rect 30432 22720 30438 22772
rect 30466 22720 30472 22772
rect 30524 22760 30530 22772
rect 30561 22763 30619 22769
rect 30561 22760 30573 22763
rect 30524 22732 30573 22760
rect 30524 22720 30530 22732
rect 30561 22729 30573 22732
rect 30607 22729 30619 22763
rect 30561 22723 30619 22729
rect 31662 22720 31668 22772
rect 31720 22760 31726 22772
rect 33229 22763 33287 22769
rect 33229 22760 33241 22763
rect 31720 22732 33241 22760
rect 31720 22720 31726 22732
rect 33229 22729 33241 22732
rect 33275 22729 33287 22763
rect 33229 22723 33287 22729
rect 34698 22720 34704 22772
rect 34756 22760 34762 22772
rect 35066 22760 35072 22772
rect 34756 22732 35072 22760
rect 34756 22720 34762 22732
rect 35066 22720 35072 22732
rect 35124 22720 35130 22772
rect 44542 22760 44548 22772
rect 38120 22732 44548 22760
rect 24728 22664 27200 22692
rect 24728 22652 24734 22664
rect 27522 22652 27528 22704
rect 27580 22652 27586 22704
rect 27614 22652 27620 22704
rect 27672 22692 27678 22704
rect 27672 22664 28396 22692
rect 27672 22652 27678 22664
rect 19705 22627 19763 22633
rect 19705 22624 19717 22627
rect 19484 22596 19717 22624
rect 19484 22584 19490 22596
rect 19705 22593 19717 22596
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 22278 22584 22284 22636
rect 22336 22624 22342 22636
rect 22830 22624 22836 22636
rect 22336 22596 22836 22624
rect 22336 22584 22342 22596
rect 22830 22584 22836 22596
rect 22888 22624 22894 22636
rect 23109 22627 23167 22633
rect 23109 22624 23121 22627
rect 22888 22596 23121 22624
rect 22888 22584 22894 22596
rect 23109 22593 23121 22596
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 24486 22584 24492 22636
rect 24544 22584 24550 22636
rect 25685 22627 25743 22633
rect 25685 22593 25697 22627
rect 25731 22624 25743 22627
rect 26786 22624 26792 22636
rect 25731 22596 26792 22624
rect 25731 22593 25743 22596
rect 25685 22587 25743 22593
rect 26786 22584 26792 22596
rect 26844 22624 26850 22636
rect 27430 22624 27436 22636
rect 26844 22596 27436 22624
rect 26844 22584 26850 22596
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 28368 22633 28396 22664
rect 28902 22652 28908 22704
rect 28960 22692 28966 22704
rect 28960 22664 29118 22692
rect 28960 22652 28966 22664
rect 29914 22652 29920 22704
rect 29972 22692 29978 22704
rect 31573 22695 31631 22701
rect 29972 22664 31524 22692
rect 29972 22652 29978 22664
rect 28353 22627 28411 22633
rect 28353 22593 28365 22627
rect 28399 22593 28411 22627
rect 28353 22587 28411 22593
rect 30926 22584 30932 22636
rect 30984 22584 30990 22636
rect 31018 22584 31024 22636
rect 31076 22584 31082 22636
rect 31496 22624 31524 22664
rect 31573 22661 31585 22695
rect 31619 22692 31631 22695
rect 31754 22692 31760 22704
rect 31619 22664 31760 22692
rect 31619 22661 31631 22664
rect 31573 22655 31631 22661
rect 31754 22652 31760 22664
rect 31812 22692 31818 22704
rect 38120 22701 38148 22732
rect 44542 22720 44548 22732
rect 44600 22720 44606 22772
rect 48590 22720 48596 22772
rect 48648 22720 48654 22772
rect 31849 22695 31907 22701
rect 31849 22692 31861 22695
rect 31812 22664 31861 22692
rect 31812 22652 31818 22664
rect 31849 22661 31861 22664
rect 31895 22692 31907 22695
rect 38105 22695 38163 22701
rect 31895 22664 37596 22692
rect 31895 22661 31907 22664
rect 31849 22655 31907 22661
rect 31662 22624 31668 22636
rect 31496 22596 31668 22624
rect 31662 22584 31668 22596
rect 31720 22584 31726 22636
rect 32398 22584 32404 22636
rect 32456 22584 32462 22636
rect 32490 22584 32496 22636
rect 32548 22624 32554 22636
rect 32953 22627 33011 22633
rect 32953 22624 32965 22627
rect 32548 22596 32965 22624
rect 32548 22584 32554 22596
rect 32953 22593 32965 22596
rect 32999 22624 33011 22627
rect 32999 22596 33548 22624
rect 32999 22593 33011 22596
rect 32953 22587 33011 22593
rect 11756 22528 11836 22556
rect 11756 22516 11762 22528
rect 12434 22516 12440 22568
rect 12492 22516 12498 22568
rect 16850 22516 16856 22568
rect 16908 22516 16914 22568
rect 19981 22559 20039 22565
rect 19981 22556 19993 22559
rect 16960 22528 19993 22556
rect 7156 22460 7972 22488
rect 7156 22448 7162 22460
rect 16206 22448 16212 22500
rect 16264 22488 16270 22500
rect 16960 22488 16988 22528
rect 19981 22525 19993 22528
rect 20027 22556 20039 22559
rect 20622 22556 20628 22568
rect 20027 22528 20628 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 20622 22516 20628 22528
rect 20680 22516 20686 22568
rect 23385 22559 23443 22565
rect 23385 22556 23397 22559
rect 23216 22528 23397 22556
rect 16264 22460 16988 22488
rect 16264 22448 16270 22460
rect 18414 22448 18420 22500
rect 18472 22488 18478 22500
rect 18601 22491 18659 22497
rect 18601 22488 18613 22491
rect 18472 22460 18613 22488
rect 18472 22448 18478 22460
rect 18601 22457 18613 22460
rect 18647 22457 18659 22491
rect 18601 22451 18659 22457
rect 21542 22448 21548 22500
rect 21600 22488 21606 22500
rect 21913 22491 21971 22497
rect 21913 22488 21925 22491
rect 21600 22460 21925 22488
rect 21600 22448 21606 22460
rect 21913 22457 21925 22460
rect 21959 22488 21971 22491
rect 22278 22488 22284 22500
rect 21959 22460 22284 22488
rect 21959 22457 21971 22460
rect 21913 22451 21971 22457
rect 22278 22448 22284 22460
rect 22336 22448 22342 22500
rect 23106 22448 23112 22500
rect 23164 22488 23170 22500
rect 23216 22488 23244 22528
rect 23385 22525 23397 22528
rect 23431 22525 23443 22559
rect 23385 22519 23443 22525
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 23532 22528 25820 22556
rect 23532 22516 23538 22528
rect 25682 22488 25688 22500
rect 23164 22460 23244 22488
rect 24872 22460 25688 22488
rect 23164 22448 23170 22460
rect 5258 22420 5264 22432
rect 3896 22392 5264 22420
rect 3421 22383 3479 22389
rect 5258 22380 5264 22392
rect 5316 22380 5322 22432
rect 6454 22380 6460 22432
rect 6512 22380 6518 22432
rect 6730 22380 6736 22432
rect 6788 22380 6794 22432
rect 6822 22380 6828 22432
rect 6880 22420 6886 22432
rect 11885 22423 11943 22429
rect 11885 22420 11897 22423
rect 6880 22392 11897 22420
rect 6880 22380 6886 22392
rect 11885 22389 11897 22392
rect 11931 22389 11943 22423
rect 11885 22383 11943 22389
rect 13446 22380 13452 22432
rect 13504 22420 13510 22432
rect 14185 22423 14243 22429
rect 14185 22420 14197 22423
rect 13504 22392 14197 22420
rect 13504 22380 13510 22392
rect 14185 22389 14197 22392
rect 14231 22389 14243 22423
rect 14185 22383 14243 22389
rect 17494 22380 17500 22432
rect 17552 22420 17558 22432
rect 17678 22420 17684 22432
rect 17552 22392 17684 22420
rect 17552 22380 17558 22392
rect 17678 22380 17684 22392
rect 17736 22420 17742 22432
rect 18506 22420 18512 22432
rect 17736 22392 18512 22420
rect 17736 22380 17742 22392
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 19061 22423 19119 22429
rect 19061 22389 19073 22423
rect 19107 22420 19119 22423
rect 19150 22420 19156 22432
rect 19107 22392 19156 22420
rect 19107 22389 19119 22392
rect 19061 22383 19119 22389
rect 19150 22380 19156 22392
rect 19208 22380 19214 22432
rect 19794 22380 19800 22432
rect 19852 22420 19858 22432
rect 20162 22420 20168 22432
rect 19852 22392 20168 22420
rect 19852 22380 19858 22392
rect 20162 22380 20168 22392
rect 20220 22380 20226 22432
rect 22094 22380 22100 22432
rect 22152 22420 22158 22432
rect 22189 22423 22247 22429
rect 22189 22420 22201 22423
rect 22152 22392 22201 22420
rect 22152 22380 22158 22392
rect 22189 22389 22201 22392
rect 22235 22420 22247 22423
rect 23842 22420 23848 22432
rect 22235 22392 23848 22420
rect 22235 22389 22247 22392
rect 22189 22383 22247 22389
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 23934 22380 23940 22432
rect 23992 22420 23998 22432
rect 24872 22429 24900 22460
rect 25682 22448 25688 22460
rect 25740 22448 25746 22500
rect 25792 22488 25820 22528
rect 25866 22516 25872 22568
rect 25924 22516 25930 22568
rect 26418 22516 26424 22568
rect 26476 22556 26482 22568
rect 26970 22556 26976 22568
rect 26476 22528 26976 22556
rect 26476 22516 26482 22528
rect 26970 22516 26976 22528
rect 27028 22516 27034 22568
rect 27246 22516 27252 22568
rect 27304 22556 27310 22568
rect 27617 22559 27675 22565
rect 27617 22556 27629 22559
rect 27304 22528 27629 22556
rect 27304 22516 27310 22528
rect 27617 22525 27629 22528
rect 27663 22525 27675 22559
rect 27617 22519 27675 22525
rect 27709 22559 27767 22565
rect 27709 22525 27721 22559
rect 27755 22525 27767 22559
rect 27709 22519 27767 22525
rect 25792 22460 27016 22488
rect 24857 22423 24915 22429
rect 24857 22420 24869 22423
rect 23992 22392 24869 22420
rect 23992 22380 23998 22392
rect 24857 22389 24869 22392
rect 24903 22389 24915 22423
rect 24857 22383 24915 22389
rect 25314 22380 25320 22432
rect 25372 22380 25378 22432
rect 26510 22380 26516 22432
rect 26568 22420 26574 22432
rect 26697 22423 26755 22429
rect 26697 22420 26709 22423
rect 26568 22392 26709 22420
rect 26568 22380 26574 22392
rect 26697 22389 26709 22392
rect 26743 22389 26755 22423
rect 26988 22420 27016 22460
rect 27338 22448 27344 22500
rect 27396 22488 27402 22500
rect 27724 22488 27752 22519
rect 28718 22516 28724 22568
rect 28776 22556 28782 22568
rect 31113 22559 31171 22565
rect 31113 22556 31125 22559
rect 28776 22528 31125 22556
rect 28776 22516 28782 22528
rect 31113 22525 31125 22528
rect 31159 22525 31171 22559
rect 31113 22519 31171 22525
rect 31202 22516 31208 22568
rect 31260 22556 31266 22568
rect 33520 22556 33548 22596
rect 33594 22584 33600 22636
rect 33652 22584 33658 22636
rect 33870 22584 33876 22636
rect 33928 22584 33934 22636
rect 34974 22584 34980 22636
rect 35032 22584 35038 22636
rect 37568 22633 37596 22664
rect 38105 22661 38117 22695
rect 38151 22661 38163 22695
rect 39942 22692 39948 22704
rect 39330 22664 39948 22692
rect 38105 22655 38163 22661
rect 39942 22652 39948 22664
rect 40000 22652 40006 22704
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22624 37611 22627
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37599 22596 37841 22624
rect 37599 22593 37611 22596
rect 37553 22587 37611 22593
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 48777 22627 48835 22633
rect 48777 22593 48789 22627
rect 48823 22624 48835 22627
rect 49053 22627 49111 22633
rect 49053 22624 49065 22627
rect 48823 22596 49065 22624
rect 48823 22593 48835 22596
rect 48777 22587 48835 22593
rect 49053 22593 49065 22596
rect 49099 22624 49111 22627
rect 49234 22624 49240 22636
rect 49099 22596 49240 22624
rect 49099 22593 49111 22596
rect 49053 22587 49111 22593
rect 49234 22584 49240 22596
rect 49292 22584 49298 22636
rect 34422 22556 34428 22568
rect 31260 22528 33364 22556
rect 33520 22528 34428 22556
rect 31260 22516 31266 22528
rect 31478 22488 31484 22500
rect 27396 22460 27752 22488
rect 30024 22460 31484 22488
rect 27396 22448 27402 22460
rect 28258 22420 28264 22432
rect 26988 22392 28264 22420
rect 26697 22383 26755 22389
rect 28258 22380 28264 22392
rect 28316 22380 28322 22432
rect 28616 22423 28674 22429
rect 28616 22389 28628 22423
rect 28662 22420 28674 22423
rect 30024 22420 30052 22460
rect 31478 22448 31484 22460
rect 31536 22448 31542 22500
rect 33045 22491 33103 22497
rect 33045 22488 33057 22491
rect 31726 22460 33057 22488
rect 28662 22392 30052 22420
rect 28662 22389 28674 22392
rect 28616 22383 28674 22389
rect 30098 22380 30104 22432
rect 30156 22380 30162 22432
rect 30926 22380 30932 22432
rect 30984 22420 30990 22432
rect 31726 22420 31754 22460
rect 33045 22457 33057 22460
rect 33091 22457 33103 22491
rect 33045 22451 33103 22457
rect 30984 22392 31754 22420
rect 30984 22380 30990 22392
rect 32490 22380 32496 22432
rect 32548 22380 32554 22432
rect 33336 22420 33364 22528
rect 34422 22516 34428 22528
rect 34480 22516 34486 22568
rect 34606 22516 34612 22568
rect 34664 22556 34670 22568
rect 39577 22559 39635 22565
rect 39577 22556 39589 22559
rect 34664 22528 39589 22556
rect 34664 22516 34670 22528
rect 39577 22525 39589 22528
rect 39623 22525 39635 22559
rect 39577 22519 39635 22525
rect 33410 22448 33416 22500
rect 33468 22488 33474 22500
rect 34701 22491 34759 22497
rect 34701 22488 34713 22491
rect 33468 22460 34713 22488
rect 33468 22448 33474 22460
rect 34701 22457 34713 22460
rect 34747 22457 34759 22491
rect 34701 22451 34759 22457
rect 35345 22423 35403 22429
rect 35345 22420 35357 22423
rect 33336 22392 35357 22420
rect 35345 22389 35357 22392
rect 35391 22420 35403 22423
rect 35710 22420 35716 22432
rect 35391 22392 35716 22420
rect 35391 22389 35403 22392
rect 35345 22383 35403 22389
rect 35710 22380 35716 22392
rect 35768 22380 35774 22432
rect 48314 22380 48320 22432
rect 48372 22420 48378 22432
rect 49237 22423 49295 22429
rect 49237 22420 49249 22423
rect 48372 22392 49249 22420
rect 48372 22380 48378 22392
rect 49237 22389 49249 22392
rect 49283 22389 49295 22423
rect 49237 22383 49295 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 2280 22188 2774 22216
rect 2280 22176 2286 22188
rect 2746 22148 2774 22188
rect 6454 22176 6460 22228
rect 6512 22216 6518 22228
rect 14182 22216 14188 22228
rect 6512 22188 14188 22216
rect 6512 22176 6518 22188
rect 14182 22176 14188 22188
rect 14240 22176 14246 22228
rect 16114 22216 16120 22228
rect 14292 22188 16120 22216
rect 3694 22148 3700 22160
rect 2746 22120 3700 22148
rect 3694 22108 3700 22120
rect 3752 22108 3758 22160
rect 3988 22120 4568 22148
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3234 22040 3240 22092
rect 3292 22080 3298 22092
rect 3513 22083 3571 22089
rect 3513 22080 3525 22083
rect 3292 22052 3525 22080
rect 3292 22040 3298 22052
rect 3513 22049 3525 22052
rect 3559 22049 3571 22083
rect 3513 22043 3571 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 3988 22012 4016 22120
rect 4246 22040 4252 22092
rect 4304 22080 4310 22092
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 4304 22052 4445 22080
rect 4304 22040 4310 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4540 22080 4568 22120
rect 4798 22108 4804 22160
rect 4856 22148 4862 22160
rect 14292 22148 14320 22188
rect 16114 22176 16120 22188
rect 16172 22176 16178 22228
rect 16390 22176 16396 22228
rect 16448 22216 16454 22228
rect 16448 22188 19656 22216
rect 16448 22176 16454 22188
rect 4856 22120 14320 22148
rect 4856 22108 4862 22120
rect 15102 22108 15108 22160
rect 15160 22148 15166 22160
rect 15160 22120 15700 22148
rect 15160 22108 15166 22120
rect 6822 22080 6828 22092
rect 4540 22052 6828 22080
rect 4433 22043 4491 22049
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 7006 22040 7012 22092
rect 7064 22080 7070 22092
rect 7285 22083 7343 22089
rect 7285 22080 7297 22083
rect 7064 22052 7297 22080
rect 7064 22040 7070 22052
rect 7285 22049 7297 22052
rect 7331 22049 7343 22083
rect 9858 22080 9864 22092
rect 7285 22043 7343 22049
rect 8496 22052 9864 22080
rect 1811 21984 4016 22012
rect 4157 22015 4215 22021
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 4157 21981 4169 22015
rect 4203 21981 4215 22015
rect 4157 21975 4215 21981
rect 6273 22015 6331 22021
rect 6273 21981 6285 22015
rect 6319 22012 6331 22015
rect 6546 22012 6552 22024
rect 6319 21984 6552 22012
rect 6319 21981 6331 21984
rect 6273 21975 6331 21981
rect 2498 21904 2504 21956
rect 2556 21944 2562 21956
rect 4172 21944 4200 21975
rect 6546 21972 6552 21984
rect 6604 21972 6610 22024
rect 6917 22015 6975 22021
rect 6917 21981 6929 22015
rect 6963 22012 6975 22015
rect 7558 22012 7564 22024
rect 6963 21984 7564 22012
rect 6963 21981 6975 21984
rect 6917 21975 6975 21981
rect 7558 21972 7564 21984
rect 7616 21972 7622 22024
rect 8496 21944 8524 22052
rect 9858 22040 9864 22052
rect 9916 22040 9922 22092
rect 9953 22083 10011 22089
rect 9953 22049 9965 22083
rect 9999 22049 10011 22083
rect 9953 22043 10011 22049
rect 8754 21972 8760 22024
rect 8812 21972 8818 22024
rect 9766 21972 9772 22024
rect 9824 21972 9830 22024
rect 9968 22012 9996 22043
rect 11238 22040 11244 22092
rect 11296 22040 11302 22092
rect 12618 22040 12624 22092
rect 12676 22080 12682 22092
rect 12676 22052 12756 22080
rect 12676 22040 12682 22052
rect 10042 22012 10048 22024
rect 9968 21984 10048 22012
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10502 21972 10508 22024
rect 10560 22012 10566 22024
rect 10778 22012 10784 22024
rect 10560 21984 10784 22012
rect 10560 21972 10566 21984
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 21981 12587 22015
rect 12728 22012 12756 22052
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 13538 22040 13544 22092
rect 13596 22080 13602 22092
rect 15672 22089 15700 22120
rect 18506 22108 18512 22160
rect 18564 22148 18570 22160
rect 19628 22148 19656 22188
rect 20254 22176 20260 22228
rect 20312 22216 20318 22228
rect 21266 22216 21272 22228
rect 20312 22188 21272 22216
rect 20312 22176 20318 22188
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 23290 22216 23296 22228
rect 21376 22188 23296 22216
rect 21376 22148 21404 22188
rect 23290 22176 23296 22188
rect 23348 22176 23354 22228
rect 26234 22216 26240 22228
rect 25148 22188 26240 22216
rect 18564 22120 19564 22148
rect 19628 22120 21404 22148
rect 18564 22108 18570 22120
rect 15657 22083 15715 22089
rect 13596 22052 14780 22080
rect 13596 22040 13602 22052
rect 14553 22015 14611 22021
rect 14553 22012 14565 22015
rect 12728 21984 14565 22012
rect 12529 21975 12587 21981
rect 14553 21981 14565 21984
rect 14599 21981 14611 22015
rect 14553 21975 14611 21981
rect 2556 21916 4200 21944
rect 5736 21916 8524 21944
rect 8573 21947 8631 21953
rect 2556 21904 2562 21916
rect 3421 21879 3479 21885
rect 3421 21845 3433 21879
rect 3467 21876 3479 21879
rect 5736 21876 5764 21916
rect 8573 21913 8585 21947
rect 8619 21944 8631 21947
rect 12544 21944 12572 21975
rect 13906 21944 13912 21956
rect 8619 21916 9812 21944
rect 8619 21913 8631 21916
rect 8573 21907 8631 21913
rect 3467 21848 5764 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 5810 21836 5816 21888
rect 5868 21836 5874 21888
rect 6086 21836 6092 21888
rect 6144 21836 6150 21888
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 8202 21876 8208 21888
rect 6972 21848 8208 21876
rect 6972 21836 6978 21848
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 8662 21836 8668 21888
rect 8720 21876 8726 21888
rect 8941 21879 8999 21885
rect 8941 21876 8953 21879
rect 8720 21848 8953 21876
rect 8720 21836 8726 21848
rect 8941 21845 8953 21848
rect 8987 21876 8999 21879
rect 9030 21876 9036 21888
rect 8987 21848 9036 21876
rect 8987 21845 8999 21848
rect 8941 21839 8999 21845
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9674 21836 9680 21888
rect 9732 21836 9738 21888
rect 9784 21876 9812 21916
rect 9968 21916 13912 21944
rect 9968 21876 9996 21916
rect 13906 21904 13912 21916
rect 13964 21904 13970 21956
rect 14369 21947 14427 21953
rect 14369 21913 14381 21947
rect 14415 21944 14427 21947
rect 14642 21944 14648 21956
rect 14415 21916 14648 21944
rect 14415 21913 14427 21916
rect 14369 21907 14427 21913
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 14752 21944 14780 22052
rect 15657 22049 15669 22083
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 17129 22083 17187 22089
rect 17129 22049 17141 22083
rect 17175 22080 17187 22083
rect 19426 22080 19432 22092
rect 17175 22052 19432 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 19536 22080 19564 22120
rect 22002 22108 22008 22160
rect 22060 22148 22066 22160
rect 23750 22148 23756 22160
rect 22060 22120 23756 22148
rect 22060 22108 22066 22120
rect 23750 22108 23756 22120
rect 23808 22108 23814 22160
rect 24394 22148 24400 22160
rect 23952 22120 24400 22148
rect 20073 22083 20131 22089
rect 19536 22052 19748 22080
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 19610 22012 19616 22024
rect 18932 21984 19616 22012
rect 18932 21972 18938 21984
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 19720 22012 19748 22052
rect 20073 22049 20085 22083
rect 20119 22080 20131 22083
rect 21542 22080 21548 22092
rect 20119 22052 21548 22080
rect 20119 22049 20131 22052
rect 20073 22043 20131 22049
rect 21542 22040 21548 22052
rect 21600 22040 21606 22092
rect 23952 22089 23980 22120
rect 24394 22108 24400 22120
rect 24452 22108 24458 22160
rect 25148 22089 25176 22188
rect 26234 22176 26240 22188
rect 26292 22176 26298 22228
rect 27338 22176 27344 22228
rect 27396 22216 27402 22228
rect 27525 22219 27583 22225
rect 27525 22216 27537 22219
rect 27396 22188 27537 22216
rect 27396 22176 27402 22188
rect 27525 22185 27537 22188
rect 27571 22185 27583 22219
rect 27525 22179 27583 22185
rect 28350 22176 28356 22228
rect 28408 22216 28414 22228
rect 29549 22219 29607 22225
rect 29549 22216 29561 22219
rect 28408 22188 29561 22216
rect 28408 22176 28414 22188
rect 29549 22185 29561 22188
rect 29595 22216 29607 22219
rect 29733 22219 29791 22225
rect 29733 22216 29745 22219
rect 29595 22188 29745 22216
rect 29595 22185 29607 22188
rect 29549 22179 29607 22185
rect 29733 22185 29745 22188
rect 29779 22185 29791 22219
rect 31846 22216 31852 22228
rect 29733 22179 29791 22185
rect 30300 22188 31852 22216
rect 30300 22160 30328 22188
rect 31846 22176 31852 22188
rect 31904 22176 31910 22228
rect 32214 22176 32220 22228
rect 32272 22216 32278 22228
rect 32858 22216 32864 22228
rect 32272 22188 32864 22216
rect 32272 22176 32278 22188
rect 32858 22176 32864 22188
rect 32916 22216 32922 22228
rect 33873 22219 33931 22225
rect 33873 22216 33885 22219
rect 32916 22188 33885 22216
rect 32916 22176 32922 22188
rect 33873 22185 33885 22188
rect 33919 22185 33931 22219
rect 33873 22179 33931 22185
rect 28994 22108 29000 22160
rect 29052 22108 29058 22160
rect 29178 22108 29184 22160
rect 29236 22148 29242 22160
rect 30282 22148 30288 22160
rect 29236 22120 30288 22148
rect 29236 22108 29242 22120
rect 30282 22108 30288 22120
rect 30340 22108 30346 22160
rect 31478 22148 31484 22160
rect 30668 22120 31484 22148
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22049 23995 22083
rect 23937 22043 23995 22049
rect 25133 22083 25191 22089
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 26694 22080 26700 22092
rect 25133 22043 25191 22049
rect 25700 22052 26700 22080
rect 20254 22012 20260 22024
rect 19720 21984 20260 22012
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 21266 21972 21272 22024
rect 21324 21972 21330 22024
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 22244 21984 22293 22012
rect 22244 21972 22250 21984
rect 22281 21981 22293 21984
rect 22327 22012 22339 22015
rect 23566 22012 23572 22024
rect 22327 21984 23572 22012
rect 22327 21981 22339 21984
rect 22281 21975 22339 21981
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 23658 21972 23664 22024
rect 23716 21972 23722 22024
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 24670 22012 24676 22024
rect 23799 21984 24676 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 24670 21972 24676 21984
rect 24728 21972 24734 22024
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 22012 25099 22015
rect 25700 22012 25728 22052
rect 26694 22040 26700 22052
rect 26752 22040 26758 22092
rect 26786 22040 26792 22092
rect 26844 22080 26850 22092
rect 29012 22080 29040 22108
rect 29273 22083 29331 22089
rect 29273 22080 29285 22083
rect 26844 22052 28948 22080
rect 29012 22052 29285 22080
rect 26844 22040 26850 22052
rect 25087 21984 25728 22012
rect 25087 21981 25099 21984
rect 25041 21975 25099 21981
rect 25774 21972 25780 22024
rect 25832 21972 25838 22024
rect 27062 21972 27068 22024
rect 27120 22012 27126 22024
rect 27338 22012 27344 22024
rect 27120 21984 27344 22012
rect 27120 21972 27126 21984
rect 27338 21972 27344 21984
rect 27396 21972 27402 22024
rect 28258 21972 28264 22024
rect 28316 22012 28322 22024
rect 28813 22015 28871 22021
rect 28813 22012 28825 22015
rect 28316 21984 28825 22012
rect 28316 21972 28322 21984
rect 28813 21981 28825 21984
rect 28859 21981 28871 22015
rect 28920 22012 28948 22052
rect 29273 22049 29285 22052
rect 29319 22049 29331 22083
rect 29273 22043 29331 22049
rect 29822 22040 29828 22092
rect 29880 22080 29886 22092
rect 30374 22080 30380 22092
rect 29880 22052 30380 22080
rect 29880 22040 29886 22052
rect 30374 22040 30380 22052
rect 30432 22040 30438 22092
rect 30668 22089 30696 22120
rect 31478 22108 31484 22120
rect 31536 22108 31542 22160
rect 30653 22083 30711 22089
rect 30653 22049 30665 22083
rect 30699 22049 30711 22083
rect 30653 22043 30711 22049
rect 31110 22040 31116 22092
rect 31168 22080 31174 22092
rect 31849 22083 31907 22089
rect 31849 22080 31861 22083
rect 31168 22052 31861 22080
rect 31168 22040 31174 22052
rect 31849 22049 31861 22052
rect 31895 22049 31907 22083
rect 31849 22043 31907 22049
rect 32674 22040 32680 22092
rect 32732 22080 32738 22092
rect 34241 22083 34299 22089
rect 34241 22080 34253 22083
rect 32732 22052 34253 22080
rect 32732 22040 32738 22052
rect 34241 22049 34253 22052
rect 34287 22049 34299 22083
rect 34241 22043 34299 22049
rect 28920 21984 30328 22012
rect 28813 21975 28871 21981
rect 17126 21944 17132 21956
rect 14752 21916 17132 21944
rect 17126 21904 17132 21916
rect 17184 21904 17190 21956
rect 17402 21904 17408 21956
rect 17460 21904 17466 21956
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 17862 21944 17868 21956
rect 17736 21916 17868 21944
rect 17736 21904 17742 21916
rect 17862 21904 17868 21916
rect 17920 21904 17926 21956
rect 19521 21947 19579 21953
rect 19521 21944 19533 21947
rect 18800 21916 19533 21944
rect 9784 21848 9996 21876
rect 11514 21836 11520 21888
rect 11572 21876 11578 21888
rect 14090 21876 14096 21888
rect 11572 21848 14096 21876
rect 11572 21836 11578 21848
rect 14090 21836 14096 21848
rect 14148 21836 14154 21888
rect 14918 21836 14924 21888
rect 14976 21876 14982 21888
rect 18800 21876 18828 21916
rect 19521 21913 19533 21916
rect 19567 21913 19579 21947
rect 19521 21907 19579 21913
rect 19705 21947 19763 21953
rect 19705 21913 19717 21947
rect 19751 21944 19763 21947
rect 19794 21944 19800 21956
rect 19751 21916 19800 21944
rect 19751 21913 19763 21916
rect 19705 21907 19763 21913
rect 19794 21904 19800 21916
rect 19852 21904 19858 21956
rect 22649 21947 22707 21953
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 22695 21916 24961 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 26053 21947 26111 21953
rect 26053 21913 26065 21947
rect 26099 21944 26111 21947
rect 26326 21944 26332 21956
rect 26099 21916 26332 21944
rect 26099 21913 26111 21916
rect 26053 21907 26111 21913
rect 26326 21904 26332 21916
rect 26384 21904 26390 21956
rect 28828 21944 28856 21975
rect 29914 21944 29920 21956
rect 28828 21916 29920 21944
rect 29914 21904 29920 21916
rect 29972 21904 29978 21956
rect 14976 21848 18828 21876
rect 18877 21879 18935 21885
rect 14976 21836 14982 21848
rect 18877 21845 18889 21879
rect 18923 21876 18935 21879
rect 18966 21876 18972 21888
rect 18923 21848 18972 21876
rect 18923 21845 18935 21848
rect 18877 21839 18935 21845
rect 18966 21836 18972 21848
rect 19024 21836 19030 21888
rect 19058 21836 19064 21888
rect 19116 21876 19122 21888
rect 22002 21876 22008 21888
rect 19116 21848 22008 21876
rect 19116 21836 19122 21848
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 22094 21836 22100 21888
rect 22152 21836 22158 21888
rect 23290 21836 23296 21888
rect 23348 21836 23354 21888
rect 24302 21836 24308 21888
rect 24360 21876 24366 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 24360 21848 24593 21876
rect 24360 21836 24366 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25958 21836 25964 21888
rect 26016 21876 26022 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 26016 21848 27997 21876
rect 26016 21836 26022 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 27985 21839 28043 21845
rect 28442 21836 28448 21888
rect 28500 21876 28506 21888
rect 28629 21879 28687 21885
rect 28629 21876 28641 21879
rect 28500 21848 28641 21876
rect 28500 21836 28506 21848
rect 28629 21845 28641 21848
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 28994 21836 29000 21888
rect 29052 21876 29058 21888
rect 30101 21879 30159 21885
rect 30101 21876 30113 21879
rect 29052 21848 30113 21876
rect 29052 21836 29058 21848
rect 30101 21845 30113 21848
rect 30147 21845 30159 21879
rect 30300 21876 30328 21984
rect 30466 21972 30472 22024
rect 30524 21972 30530 22024
rect 32585 22015 32643 22021
rect 31128 21984 32536 22012
rect 30561 21947 30619 21953
rect 30561 21913 30573 21947
rect 30607 21944 30619 21947
rect 31128 21944 31156 21984
rect 30607 21916 31156 21944
rect 30607 21913 30619 21916
rect 30561 21907 30619 21913
rect 31202 21904 31208 21956
rect 31260 21944 31266 21956
rect 31389 21947 31447 21953
rect 31389 21944 31401 21947
rect 31260 21916 31401 21944
rect 31260 21904 31266 21916
rect 31389 21913 31401 21916
rect 31435 21944 31447 21947
rect 32217 21947 32275 21953
rect 32217 21944 32229 21947
rect 31435 21916 32229 21944
rect 31435 21913 31447 21916
rect 31389 21907 31447 21913
rect 32217 21913 32229 21916
rect 32263 21913 32275 21947
rect 32508 21944 32536 21984
rect 32585 21981 32597 22015
rect 32631 22012 32643 22015
rect 32766 22012 32772 22024
rect 32631 21984 32772 22012
rect 32631 21981 32643 21984
rect 32585 21975 32643 21981
rect 32766 21972 32772 21984
rect 32824 21972 32830 22024
rect 32858 21972 32864 22024
rect 32916 21972 32922 22024
rect 33318 21972 33324 22024
rect 33376 22012 33382 22024
rect 34057 22015 34115 22021
rect 34057 22012 34069 22015
rect 33376 21984 34069 22012
rect 33376 21972 33382 21984
rect 34057 21981 34069 21984
rect 34103 21981 34115 22015
rect 34057 21975 34115 21981
rect 48777 22015 48835 22021
rect 48777 21981 48789 22015
rect 48823 22012 48835 22015
rect 49050 22012 49056 22024
rect 48823 21984 49056 22012
rect 48823 21981 48835 21984
rect 48777 21975 48835 21981
rect 49050 21972 49056 21984
rect 49108 21972 49114 22024
rect 35250 21944 35256 21956
rect 32508 21916 35256 21944
rect 32217 21907 32275 21913
rect 35250 21904 35256 21916
rect 35308 21904 35314 21956
rect 31481 21879 31539 21885
rect 31481 21876 31493 21879
rect 30300 21848 31493 21876
rect 30101 21839 30159 21845
rect 31481 21845 31493 21848
rect 31527 21845 31539 21879
rect 31481 21839 31539 21845
rect 31662 21836 31668 21888
rect 31720 21876 31726 21888
rect 32033 21879 32091 21885
rect 32033 21876 32045 21879
rect 31720 21848 32045 21876
rect 31720 21836 31726 21848
rect 32033 21845 32045 21848
rect 32079 21845 32091 21879
rect 32033 21839 32091 21845
rect 32398 21836 32404 21888
rect 32456 21876 32462 21888
rect 33689 21879 33747 21885
rect 33689 21876 33701 21879
rect 32456 21848 33701 21876
rect 32456 21836 32462 21848
rect 33689 21845 33701 21848
rect 33735 21845 33747 21879
rect 33689 21839 33747 21845
rect 49234 21836 49240 21888
rect 49292 21836 49298 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 5718 21672 5724 21684
rect 1780 21644 5724 21672
rect 1780 21545 1808 21644
rect 5718 21632 5724 21644
rect 5776 21632 5782 21684
rect 5810 21632 5816 21684
rect 5868 21672 5874 21684
rect 9401 21675 9459 21681
rect 5868 21644 9352 21672
rect 5868 21632 5874 21644
rect 3970 21564 3976 21616
rect 4028 21604 4034 21616
rect 6178 21604 6184 21616
rect 4028 21576 6184 21604
rect 4028 21564 4034 21576
rect 6178 21564 6184 21576
rect 6236 21564 6242 21616
rect 6270 21564 6276 21616
rect 6328 21604 6334 21616
rect 7374 21604 7380 21616
rect 6328 21576 7380 21604
rect 6328 21564 6334 21576
rect 7374 21564 7380 21576
rect 7432 21604 7438 21616
rect 7929 21607 7987 21613
rect 7929 21604 7941 21607
rect 7432 21576 7941 21604
rect 7432 21564 7438 21576
rect 7929 21573 7941 21576
rect 7975 21573 7987 21607
rect 7929 21567 7987 21573
rect 8662 21564 8668 21616
rect 8720 21564 8726 21616
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 2222 21496 2228 21548
rect 2280 21536 2286 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 2280 21508 3433 21536
rect 2280 21496 2286 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 7006 21496 7012 21548
rect 7064 21496 7070 21548
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7576 21508 7665 21536
rect 2774 21428 2780 21480
rect 2832 21428 2838 21480
rect 3326 21428 3332 21480
rect 3384 21468 3390 21480
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 3384 21440 3893 21468
rect 3384 21428 3390 21440
rect 3881 21437 3893 21440
rect 3927 21437 3939 21471
rect 5258 21468 5264 21480
rect 3881 21431 3939 21437
rect 4448 21440 5264 21468
rect 3418 21360 3424 21412
rect 3476 21400 3482 21412
rect 4448 21400 4476 21440
rect 5258 21428 5264 21440
rect 5316 21428 5322 21480
rect 5350 21428 5356 21480
rect 5408 21468 5414 21480
rect 5721 21471 5779 21477
rect 5721 21468 5733 21471
rect 5408 21440 5733 21468
rect 5408 21428 5414 21440
rect 5721 21437 5733 21440
rect 5767 21437 5779 21471
rect 5721 21431 5779 21437
rect 5810 21428 5816 21480
rect 5868 21428 5874 21480
rect 5920 21440 6960 21468
rect 5920 21400 5948 21440
rect 3476 21372 4476 21400
rect 4540 21372 5948 21400
rect 6457 21403 6515 21409
rect 3476 21360 3482 21372
rect 2130 21292 2136 21344
rect 2188 21332 2194 21344
rect 4540 21332 4568 21372
rect 6457 21369 6469 21403
rect 6503 21400 6515 21403
rect 6822 21400 6828 21412
rect 6503 21372 6828 21400
rect 6503 21369 6515 21372
rect 6457 21363 6515 21369
rect 6822 21360 6828 21372
rect 6880 21360 6886 21412
rect 6932 21400 6960 21440
rect 7193 21403 7251 21409
rect 7193 21400 7205 21403
rect 6932 21372 7205 21400
rect 7193 21369 7205 21372
rect 7239 21369 7251 21403
rect 7576 21400 7604 21508
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 8938 21496 8944 21548
rect 8996 21496 9002 21548
rect 9324 21536 9352 21644
rect 9401 21641 9413 21675
rect 9447 21641 9459 21675
rect 9401 21635 9459 21641
rect 9416 21604 9444 21635
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 9732 21644 10241 21672
rect 9732 21632 9738 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 10229 21635 10287 21641
rect 10962 21632 10968 21684
rect 11020 21632 11026 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 16025 21675 16083 21681
rect 11195 21644 15976 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 15948 21616 15976 21644
rect 16025 21641 16037 21675
rect 16071 21672 16083 21675
rect 16298 21672 16304 21684
rect 16071 21644 16304 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 16666 21632 16672 21684
rect 16724 21672 16730 21684
rect 18966 21672 18972 21684
rect 16724 21644 18972 21672
rect 16724 21632 16730 21644
rect 18966 21632 18972 21644
rect 19024 21632 19030 21684
rect 19610 21632 19616 21684
rect 19668 21672 19674 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 19668 21644 22017 21672
rect 19668 21632 19674 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22005 21635 22063 21641
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23017 21675 23075 21681
rect 23017 21672 23029 21675
rect 22888 21644 23029 21672
rect 22888 21632 22894 21644
rect 23017 21641 23029 21644
rect 23063 21641 23075 21675
rect 23017 21635 23075 21641
rect 9582 21604 9588 21616
rect 9416 21576 9588 21604
rect 9582 21564 9588 21576
rect 9640 21604 9646 21616
rect 15286 21604 15292 21616
rect 9640 21576 12388 21604
rect 14582 21576 15292 21604
rect 9640 21564 9646 21576
rect 9324 21508 10640 21536
rect 8956 21468 8984 21496
rect 7760 21440 8984 21468
rect 7760 21400 7788 21440
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 10321 21471 10379 21477
rect 10321 21468 10333 21471
rect 9456 21440 10333 21468
rect 9456 21428 9462 21440
rect 10321 21437 10333 21440
rect 10367 21437 10379 21471
rect 10321 21431 10379 21437
rect 10505 21471 10563 21477
rect 10505 21437 10517 21471
rect 10551 21437 10563 21471
rect 10612 21468 10640 21508
rect 12158 21496 12164 21548
rect 12216 21496 12222 21548
rect 12250 21468 12256 21480
rect 10612 21440 12256 21468
rect 10505 21431 10563 21437
rect 7576 21372 7788 21400
rect 10520 21400 10548 21431
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 12360 21477 12388 21576
rect 15286 21564 15292 21576
rect 15344 21564 15350 21616
rect 15930 21564 15936 21616
rect 15988 21564 15994 21616
rect 16574 21564 16580 21616
rect 16632 21604 16638 21616
rect 16758 21604 16764 21616
rect 16632 21576 16764 21604
rect 16632 21564 16638 21576
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 17494 21564 17500 21616
rect 17552 21604 17558 21616
rect 19058 21604 19064 21616
rect 17552 21576 19064 21604
rect 17552 21564 17558 21576
rect 19058 21564 19064 21576
rect 19116 21564 19122 21616
rect 20254 21604 20260 21616
rect 20194 21576 20260 21604
rect 20254 21564 20260 21576
rect 20312 21604 20318 21616
rect 20990 21604 20996 21616
rect 20312 21576 20996 21604
rect 20312 21564 20318 21576
rect 20990 21564 20996 21576
rect 21048 21564 21054 21616
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 14568 21508 16865 21536
rect 12345 21471 12403 21477
rect 12345 21437 12357 21471
rect 12391 21437 12403 21471
rect 12345 21431 12403 21437
rect 12434 21428 12440 21480
rect 12492 21468 12498 21480
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12492 21440 13093 21468
rect 12492 21428 12498 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 12710 21400 12716 21412
rect 10520 21372 12716 21400
rect 7193 21363 7251 21369
rect 12710 21360 12716 21372
rect 12768 21360 12774 21412
rect 2188 21304 4568 21332
rect 5261 21335 5319 21341
rect 2188 21292 2194 21304
rect 5261 21301 5273 21335
rect 5307 21332 5319 21335
rect 5534 21332 5540 21344
rect 5307 21304 5540 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 6178 21292 6184 21344
rect 6236 21332 6242 21344
rect 6641 21335 6699 21341
rect 6641 21332 6653 21335
rect 6236 21304 6653 21332
rect 6236 21292 6242 21304
rect 6641 21301 6653 21304
rect 6687 21301 6699 21335
rect 6641 21295 6699 21301
rect 9674 21292 9680 21344
rect 9732 21292 9738 21344
rect 9861 21335 9919 21341
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 11054 21332 11060 21344
rect 9907 21304 11060 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11514 21332 11520 21344
rect 11379 21304 11520 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 11790 21292 11796 21344
rect 11848 21292 11854 21344
rect 13096 21332 13124 21431
rect 13354 21428 13360 21480
rect 13412 21428 13418 21480
rect 14090 21428 14096 21480
rect 14148 21468 14154 21480
rect 14568 21468 14596 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21536 21327 21539
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 21315 21508 22385 21536
rect 21315 21505 21327 21508
rect 21269 21499 21327 21505
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 23032 21536 23060 21635
rect 24486 21632 24492 21684
rect 24544 21672 24550 21684
rect 24544 21644 24992 21672
rect 24544 21632 24550 21644
rect 23661 21607 23719 21613
rect 23661 21573 23673 21607
rect 23707 21604 23719 21607
rect 23934 21604 23940 21616
rect 23707 21576 23940 21604
rect 23707 21573 23719 21576
rect 23661 21567 23719 21573
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 24964 21604 24992 21644
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 26697 21675 26755 21681
rect 26697 21672 26709 21675
rect 25096 21644 26709 21672
rect 25096 21632 25102 21644
rect 26697 21641 26709 21644
rect 26743 21672 26755 21675
rect 27522 21672 27528 21684
rect 26743 21644 27528 21672
rect 26743 21641 26755 21644
rect 26697 21635 26755 21641
rect 27522 21632 27528 21644
rect 27580 21672 27586 21684
rect 27617 21675 27675 21681
rect 27617 21672 27629 21675
rect 27580 21644 27629 21672
rect 27580 21632 27586 21644
rect 27617 21641 27629 21644
rect 27663 21641 27675 21675
rect 27617 21635 27675 21641
rect 27709 21675 27767 21681
rect 27709 21641 27721 21675
rect 27755 21672 27767 21675
rect 30558 21672 30564 21684
rect 27755 21644 30564 21672
rect 27755 21641 27767 21644
rect 27709 21635 27767 21641
rect 30558 21632 30564 21644
rect 30616 21632 30622 21684
rect 31113 21675 31171 21681
rect 31113 21641 31125 21675
rect 31159 21672 31171 21675
rect 36722 21672 36728 21684
rect 31159 21644 36728 21672
rect 31159 21641 31171 21644
rect 31113 21635 31171 21641
rect 36722 21632 36728 21644
rect 36780 21632 36786 21684
rect 25682 21604 25688 21616
rect 24886 21576 25688 21604
rect 25682 21564 25688 21576
rect 25740 21564 25746 21616
rect 28994 21604 29000 21616
rect 27540 21576 29000 21604
rect 23382 21536 23388 21548
rect 23032 21508 23388 21536
rect 22373 21499 22431 21505
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 25958 21496 25964 21548
rect 26016 21496 26022 21548
rect 26053 21539 26111 21545
rect 26053 21505 26065 21539
rect 26099 21536 26111 21539
rect 27540 21536 27568 21576
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 31570 21564 31576 21616
rect 31628 21604 31634 21616
rect 33597 21607 33655 21613
rect 33597 21604 33609 21607
rect 31628 21576 33609 21604
rect 31628 21564 31634 21576
rect 33597 21573 33609 21576
rect 33643 21573 33655 21607
rect 33597 21567 33655 21573
rect 26099 21508 27568 21536
rect 26099 21505 26111 21508
rect 26053 21499 26111 21505
rect 29822 21496 29828 21548
rect 29880 21496 29886 21548
rect 31021 21539 31079 21545
rect 31021 21505 31033 21539
rect 31067 21536 31079 21539
rect 31938 21536 31944 21548
rect 31067 21508 31944 21536
rect 31067 21505 31079 21508
rect 31021 21499 31079 21505
rect 31938 21496 31944 21508
rect 31996 21496 32002 21548
rect 32306 21496 32312 21548
rect 32364 21536 32370 21548
rect 32401 21539 32459 21545
rect 32401 21536 32413 21539
rect 32364 21508 32413 21536
rect 32364 21496 32370 21508
rect 32401 21505 32413 21508
rect 32447 21536 32459 21539
rect 32861 21539 32919 21545
rect 32861 21536 32873 21539
rect 32447 21508 32873 21536
rect 32447 21505 32459 21508
rect 32401 21499 32459 21505
rect 32861 21505 32873 21508
rect 32907 21505 32919 21539
rect 32861 21499 32919 21505
rect 47854 21496 47860 21548
rect 47912 21536 47918 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47912 21508 47961 21536
rect 47912 21496 47918 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 14148 21440 14596 21468
rect 14148 21428 14154 21440
rect 16206 21428 16212 21480
rect 16264 21428 16270 21480
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21468 18751 21471
rect 18739 21440 18828 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 14366 21360 14372 21412
rect 14424 21400 14430 21412
rect 14424 21372 15332 21400
rect 14424 21360 14430 21372
rect 13722 21332 13728 21344
rect 13096 21304 13728 21332
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 14550 21292 14556 21344
rect 14608 21332 14614 21344
rect 15304 21341 15332 21372
rect 15562 21360 15568 21412
rect 15620 21360 15626 21412
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 14608 21304 14841 21332
rect 14608 21292 14614 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 14829 21295 14887 21301
rect 15289 21335 15347 21341
rect 15289 21301 15301 21335
rect 15335 21332 15347 21335
rect 18690 21332 18696 21344
rect 15335 21304 18696 21332
rect 15335 21301 15347 21304
rect 15289 21295 15347 21301
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 18800 21332 18828 21440
rect 18966 21428 18972 21480
rect 19024 21428 19030 21480
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 21910 21468 21916 21480
rect 19116 21440 21916 21468
rect 19116 21428 19122 21440
rect 21910 21428 21916 21440
rect 21968 21428 21974 21480
rect 22462 21428 22468 21480
rect 22520 21428 22526 21480
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 24670 21468 24676 21480
rect 22695 21440 24676 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 24670 21428 24676 21440
rect 24728 21468 24734 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24728 21440 25145 21468
rect 24728 21428 24734 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 26234 21428 26240 21480
rect 26292 21428 26298 21480
rect 26694 21428 26700 21480
rect 26752 21468 26758 21480
rect 26752 21440 27292 21468
rect 26752 21428 26758 21440
rect 20162 21360 20168 21412
rect 20220 21400 20226 21412
rect 22370 21400 22376 21412
rect 20220 21372 22376 21400
rect 20220 21360 20226 21372
rect 22370 21360 22376 21372
rect 22428 21360 22434 21412
rect 24762 21360 24768 21412
rect 24820 21400 24826 21412
rect 27264 21409 27292 21440
rect 27798 21428 27804 21480
rect 27856 21428 27862 21480
rect 28350 21428 28356 21480
rect 28408 21468 28414 21480
rect 28445 21471 28503 21477
rect 28445 21468 28457 21471
rect 28408 21440 28457 21468
rect 28408 21428 28414 21440
rect 28445 21437 28457 21440
rect 28491 21437 28503 21471
rect 28445 21431 28503 21437
rect 28718 21428 28724 21480
rect 28776 21468 28782 21480
rect 30098 21468 30104 21480
rect 28776 21440 30104 21468
rect 28776 21428 28782 21440
rect 30098 21428 30104 21440
rect 30156 21428 30162 21480
rect 31205 21471 31263 21477
rect 31205 21468 31217 21471
rect 30208 21440 31217 21468
rect 27249 21403 27307 21409
rect 24820 21372 25728 21400
rect 24820 21360 24826 21372
rect 19426 21332 19432 21344
rect 18800 21304 19432 21332
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 19702 21292 19708 21344
rect 19760 21332 19766 21344
rect 20441 21335 20499 21341
rect 20441 21332 20453 21335
rect 19760 21304 20453 21332
rect 19760 21292 19766 21304
rect 20441 21301 20453 21304
rect 20487 21301 20499 21335
rect 20441 21295 20499 21301
rect 20809 21335 20867 21341
rect 20809 21301 20821 21335
rect 20855 21332 20867 21335
rect 20990 21332 20996 21344
rect 20855 21304 20996 21332
rect 20855 21301 20867 21304
rect 20809 21295 20867 21301
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 21910 21292 21916 21344
rect 21968 21332 21974 21344
rect 24118 21332 24124 21344
rect 21968 21304 24124 21332
rect 21968 21292 21974 21304
rect 24118 21292 24124 21304
rect 24176 21292 24182 21344
rect 25222 21292 25228 21344
rect 25280 21332 25286 21344
rect 25593 21335 25651 21341
rect 25593 21332 25605 21335
rect 25280 21304 25605 21332
rect 25280 21292 25286 21304
rect 25593 21301 25605 21304
rect 25639 21301 25651 21335
rect 25700 21332 25728 21372
rect 27249 21369 27261 21403
rect 27295 21369 27307 21403
rect 27249 21363 27307 21369
rect 30208 21344 30236 21440
rect 31205 21437 31217 21440
rect 31251 21437 31263 21471
rect 33413 21471 33471 21477
rect 33413 21468 33425 21471
rect 31205 21431 31263 21437
rect 31312 21440 33425 21468
rect 30282 21360 30288 21412
rect 30340 21400 30346 21412
rect 31312 21400 31340 21440
rect 33413 21437 33425 21440
rect 33459 21437 33471 21471
rect 33413 21431 33471 21437
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 30340 21372 31340 21400
rect 30340 21360 30346 21372
rect 31386 21360 31392 21412
rect 31444 21400 31450 21412
rect 33229 21403 33287 21409
rect 33229 21400 33241 21403
rect 31444 21372 33241 21400
rect 31444 21360 31450 21372
rect 33229 21369 33241 21372
rect 33275 21369 33287 21403
rect 33229 21363 33287 21369
rect 34514 21360 34520 21412
rect 34572 21400 34578 21412
rect 37734 21400 37740 21412
rect 34572 21372 37740 21400
rect 34572 21360 34578 21372
rect 37734 21360 37740 21372
rect 37792 21360 37798 21412
rect 28442 21332 28448 21344
rect 25700 21304 28448 21332
rect 25593 21295 25651 21301
rect 28442 21292 28448 21304
rect 28500 21292 28506 21344
rect 30190 21292 30196 21344
rect 30248 21292 30254 21344
rect 30650 21292 30656 21344
rect 30708 21292 30714 21344
rect 31757 21335 31815 21341
rect 31757 21301 31769 21335
rect 31803 21332 31815 21335
rect 31846 21332 31852 21344
rect 31803 21304 31852 21332
rect 31803 21301 31815 21304
rect 31757 21295 31815 21301
rect 31846 21292 31852 21304
rect 31904 21292 31910 21344
rect 32490 21292 32496 21344
rect 32548 21292 32554 21344
rect 32766 21292 32772 21344
rect 32824 21332 32830 21344
rect 33045 21335 33103 21341
rect 33045 21332 33057 21335
rect 32824 21304 33057 21332
rect 32824 21292 32830 21304
rect 33045 21301 33057 21304
rect 33091 21301 33103 21335
rect 33045 21295 33103 21301
rect 47673 21335 47731 21341
rect 47673 21301 47685 21335
rect 47719 21332 47731 21335
rect 47854 21332 47860 21344
rect 47719 21304 47860 21332
rect 47719 21301 47731 21304
rect 47673 21295 47731 21301
rect 47854 21292 47860 21304
rect 47912 21292 47918 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 3421 21131 3479 21137
rect 3421 21097 3433 21131
rect 3467 21128 3479 21131
rect 6914 21128 6920 21140
rect 3467 21100 6920 21128
rect 3467 21097 3479 21100
rect 3421 21091 3479 21097
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 12158 21128 12164 21140
rect 7024 21100 12164 21128
rect 7024 21072 7052 21100
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 12342 21088 12348 21140
rect 12400 21128 12406 21140
rect 14918 21128 14924 21140
rect 12400 21100 14924 21128
rect 12400 21088 12406 21100
rect 14918 21088 14924 21100
rect 14976 21088 14982 21140
rect 15102 21088 15108 21140
rect 15160 21128 15166 21140
rect 15749 21131 15807 21137
rect 15749 21128 15761 21131
rect 15160 21100 15761 21128
rect 15160 21088 15166 21100
rect 15749 21097 15761 21100
rect 15795 21097 15807 21131
rect 15749 21091 15807 21097
rect 17512 21100 22416 21128
rect 7006 21020 7012 21072
rect 7064 21020 7070 21072
rect 11790 21060 11796 21072
rect 8312 21032 11796 21060
rect 4246 20952 4252 21004
rect 4304 20952 4310 21004
rect 8312 21001 8340 21032
rect 11790 21020 11796 21032
rect 11848 21020 11854 21072
rect 12250 21020 12256 21072
rect 12308 21060 12314 21072
rect 14182 21060 14188 21072
rect 12308 21032 14188 21060
rect 12308 21020 12314 21032
rect 14182 21020 14188 21032
rect 14240 21020 14246 21072
rect 14277 21063 14335 21069
rect 14277 21029 14289 21063
rect 14323 21060 14335 21063
rect 14366 21060 14372 21072
rect 14323 21032 14372 21060
rect 14323 21029 14335 21032
rect 14277 21023 14335 21029
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 14553 21063 14611 21069
rect 14553 21029 14565 21063
rect 14599 21060 14611 21063
rect 17310 21060 17316 21072
rect 14599 21032 17316 21060
rect 14599 21029 14611 21032
rect 14553 21023 14611 21029
rect 17310 21020 17316 21032
rect 17368 21020 17374 21072
rect 5721 20995 5779 21001
rect 5721 20961 5733 20995
rect 5767 20992 5779 20995
rect 8297 20995 8355 21001
rect 5767 20964 7696 20992
rect 5767 20961 5779 20964
rect 5721 20955 5779 20961
rect 7668 20936 7696 20964
rect 8297 20961 8309 20995
rect 8343 20961 8355 20995
rect 8297 20955 8355 20961
rect 8478 20952 8484 21004
rect 8536 20952 8542 21004
rect 8570 20952 8576 21004
rect 8628 20992 8634 21004
rect 9585 20995 9643 21001
rect 9585 20992 9597 20995
rect 8628 20964 9597 20992
rect 8628 20952 8634 20964
rect 9585 20961 9597 20964
rect 9631 20961 9643 20995
rect 9585 20955 9643 20961
rect 11238 20952 11244 21004
rect 11296 20992 11302 21004
rect 12066 20992 12072 21004
rect 11296 20964 12072 20992
rect 11296 20952 11302 20964
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 11992 20933 12020 20964
rect 12066 20952 12072 20964
rect 12124 20952 12130 21004
rect 12618 20952 12624 21004
rect 12676 20952 12682 21004
rect 15010 20952 15016 21004
rect 15068 20992 15074 21004
rect 15105 20995 15163 21001
rect 15105 20992 15117 20995
rect 15068 20964 15117 20992
rect 15068 20952 15074 20964
rect 15105 20961 15117 20964
rect 15151 20961 15163 20995
rect 15286 20992 15292 21004
rect 15105 20955 15163 20961
rect 15212 20964 15292 20992
rect 9309 20927 9367 20933
rect 7708 20896 8616 20924
rect 7708 20884 7714 20896
rect 8588 20868 8616 20896
rect 9309 20893 9321 20927
rect 9355 20924 9367 20927
rect 10965 20927 11023 20933
rect 9355 20896 9628 20924
rect 9355 20893 9367 20896
rect 9309 20887 9367 20893
rect 9600 20868 9628 20896
rect 10965 20893 10977 20927
rect 11011 20924 11023 20927
rect 11977 20927 12035 20933
rect 11011 20896 11652 20924
rect 11011 20893 11023 20896
rect 10965 20887 11023 20893
rect 2777 20859 2835 20865
rect 2777 20825 2789 20859
rect 2823 20856 2835 20859
rect 2866 20856 2872 20868
rect 2823 20828 2872 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 3605 20859 3663 20865
rect 3605 20825 3617 20859
rect 3651 20856 3663 20859
rect 3786 20856 3792 20868
rect 3651 20828 3792 20856
rect 3651 20825 3663 20828
rect 3605 20819 3663 20825
rect 3786 20816 3792 20828
rect 3844 20856 3850 20868
rect 5626 20856 5632 20868
rect 3844 20828 5632 20856
rect 3844 20816 3850 20828
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 6178 20856 6184 20868
rect 5736 20828 6184 20856
rect 5169 20791 5227 20797
rect 5169 20757 5181 20791
rect 5215 20788 5227 20791
rect 5736 20788 5764 20828
rect 6178 20816 6184 20828
rect 6236 20816 6242 20868
rect 7745 20859 7803 20865
rect 7745 20825 7757 20859
rect 7791 20856 7803 20859
rect 8202 20856 8208 20868
rect 7791 20828 8208 20856
rect 7791 20825 7803 20828
rect 7745 20819 7803 20825
rect 8202 20816 8208 20828
rect 8260 20816 8266 20868
rect 8570 20816 8576 20868
rect 8628 20816 8634 20868
rect 9582 20816 9588 20868
rect 9640 20816 9646 20868
rect 11330 20816 11336 20868
rect 11388 20816 11394 20868
rect 11624 20856 11652 20896
rect 11977 20893 11989 20927
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20924 13783 20927
rect 15212 20924 15240 20964
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 16390 20952 16396 21004
rect 16448 20952 16454 21004
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 17512 20992 17540 21100
rect 21821 21063 21879 21069
rect 17604 21032 18920 21060
rect 17604 21001 17632 21032
rect 17451 20964 17540 20992
rect 17589 20995 17647 21001
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 17589 20961 17601 20995
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 18690 20952 18696 21004
rect 18748 20952 18754 21004
rect 18892 20992 18920 21032
rect 21821 21029 21833 21063
rect 21867 21060 21879 21063
rect 22278 21060 22284 21072
rect 21867 21032 22284 21060
rect 21867 21029 21879 21032
rect 21821 21023 21879 21029
rect 22278 21020 22284 21032
rect 22336 21020 22342 21072
rect 22388 21060 22416 21100
rect 22462 21088 22468 21140
rect 22520 21128 22526 21140
rect 25314 21128 25320 21140
rect 22520 21100 25320 21128
rect 22520 21088 22526 21100
rect 25314 21088 25320 21100
rect 25372 21088 25378 21140
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 27801 21131 27859 21137
rect 27801 21128 27813 21131
rect 26384 21100 27813 21128
rect 26384 21088 26390 21100
rect 27801 21097 27813 21100
rect 27847 21097 27859 21131
rect 31938 21128 31944 21140
rect 27801 21091 27859 21097
rect 28966 21100 31944 21128
rect 24762 21060 24768 21072
rect 22388 21032 24768 21060
rect 24762 21020 24768 21032
rect 24820 21020 24826 21072
rect 27522 21020 27528 21072
rect 27580 21060 27586 21072
rect 28810 21060 28816 21072
rect 27580 21032 28816 21060
rect 27580 21020 27586 21032
rect 28810 21020 28816 21032
rect 28868 21060 28874 21072
rect 28966 21060 28994 21100
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 32493 21131 32551 21137
rect 32493 21097 32505 21131
rect 32539 21128 32551 21131
rect 32582 21128 32588 21140
rect 32539 21100 32588 21128
rect 32539 21097 32551 21100
rect 32493 21091 32551 21097
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 28868 21032 28994 21060
rect 28868 21020 28874 21032
rect 29178 21020 29184 21072
rect 29236 21060 29242 21072
rect 32766 21060 32772 21072
rect 29236 21032 32772 21060
rect 29236 21020 29242 21032
rect 32766 21020 32772 21032
rect 32824 21020 32830 21072
rect 19702 20992 19708 21004
rect 18892 20964 19708 20992
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 22646 20952 22652 21004
rect 22704 20952 22710 21004
rect 23842 20952 23848 21004
rect 23900 20952 23906 21004
rect 25314 20952 25320 21004
rect 25372 20952 25378 21004
rect 26329 20995 26387 21001
rect 26329 20961 26341 20995
rect 26375 20992 26387 20995
rect 27798 20992 27804 21004
rect 26375 20964 27804 20992
rect 26375 20961 26387 20964
rect 26329 20955 26387 20961
rect 27798 20952 27804 20964
rect 27856 20952 27862 21004
rect 28534 20952 28540 21004
rect 28592 20952 28598 21004
rect 30006 20952 30012 21004
rect 30064 20952 30070 21004
rect 30558 20952 30564 21004
rect 30616 20992 30622 21004
rect 31202 20992 31208 21004
rect 30616 20964 31208 20992
rect 30616 20952 30622 20964
rect 31202 20952 31208 20964
rect 31260 20952 31266 21004
rect 31662 20952 31668 21004
rect 31720 20992 31726 21004
rect 36446 20992 36452 21004
rect 31720 20964 36452 20992
rect 31720 20952 31726 20964
rect 36446 20952 36452 20964
rect 36504 20952 36510 21004
rect 19058 20924 19064 20936
rect 13771 20896 15240 20924
rect 15304 20896 19064 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 15194 20856 15200 20868
rect 11624 20828 15200 20856
rect 15194 20816 15200 20828
rect 15252 20816 15258 20868
rect 5215 20760 5764 20788
rect 5215 20757 5227 20760
rect 5169 20751 5227 20757
rect 5810 20748 5816 20800
rect 5868 20788 5874 20800
rect 6362 20788 6368 20800
rect 5868 20760 6368 20788
rect 5868 20748 5874 20760
rect 6362 20748 6368 20760
rect 6420 20748 6426 20800
rect 7006 20748 7012 20800
rect 7064 20788 7070 20800
rect 7193 20791 7251 20797
rect 7193 20788 7205 20791
rect 7064 20760 7205 20788
rect 7064 20748 7070 20760
rect 7193 20757 7205 20760
rect 7239 20757 7251 20791
rect 7193 20751 7251 20757
rect 7558 20748 7564 20800
rect 7616 20748 7622 20800
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 9398 20788 9404 20800
rect 7883 20760 9404 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 11422 20748 11428 20800
rect 11480 20748 11486 20800
rect 11606 20748 11612 20800
rect 11664 20788 11670 20800
rect 11882 20788 11888 20800
rect 11664 20760 11888 20788
rect 11664 20748 11670 20760
rect 11882 20748 11888 20760
rect 11940 20788 11946 20800
rect 13538 20788 13544 20800
rect 11940 20760 13544 20788
rect 11940 20748 11946 20760
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 13906 20748 13912 20800
rect 13964 20748 13970 20800
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 14921 20791 14979 20797
rect 14921 20788 14933 20791
rect 14424 20760 14933 20788
rect 14424 20748 14430 20760
rect 14921 20757 14933 20760
rect 14967 20757 14979 20791
rect 14921 20751 14979 20757
rect 15013 20791 15071 20797
rect 15013 20757 15025 20791
rect 15059 20788 15071 20791
rect 15304 20788 15332 20896
rect 19058 20884 19064 20896
rect 19116 20884 19122 20936
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 24210 20884 24216 20936
rect 24268 20924 24274 20936
rect 25685 20927 25743 20933
rect 25685 20924 25697 20927
rect 24268 20896 25697 20924
rect 24268 20884 24274 20896
rect 25685 20893 25697 20896
rect 25731 20924 25743 20927
rect 25774 20924 25780 20936
rect 25731 20896 25780 20924
rect 25731 20893 25743 20896
rect 25685 20887 25743 20893
rect 25774 20884 25780 20896
rect 25832 20924 25838 20936
rect 26050 20924 26056 20936
rect 25832 20896 26056 20924
rect 25832 20884 25838 20896
rect 26050 20884 26056 20896
rect 26108 20884 26114 20936
rect 28261 20927 28319 20933
rect 28261 20893 28273 20927
rect 28307 20924 28319 20927
rect 28442 20924 28448 20936
rect 28307 20896 28448 20924
rect 28307 20893 28319 20896
rect 28261 20887 28319 20893
rect 28442 20884 28448 20896
rect 28500 20924 28506 20936
rect 28902 20924 28908 20936
rect 28500 20896 28908 20924
rect 28500 20884 28506 20896
rect 28902 20884 28908 20896
rect 28960 20884 28966 20936
rect 29546 20884 29552 20936
rect 29604 20924 29610 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29604 20896 29745 20924
rect 29604 20884 29610 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 31110 20884 31116 20936
rect 31168 20884 31174 20936
rect 32674 20884 32680 20936
rect 32732 20924 32738 20936
rect 32953 20927 33011 20933
rect 32953 20924 32965 20927
rect 32732 20896 32965 20924
rect 32732 20884 32738 20896
rect 32953 20893 32965 20896
rect 32999 20893 33011 20927
rect 32953 20887 33011 20893
rect 16209 20859 16267 20865
rect 16209 20825 16221 20859
rect 16255 20856 16267 20859
rect 19702 20856 19708 20868
rect 16255 20828 19708 20856
rect 16255 20825 16267 20828
rect 16209 20819 16267 20825
rect 19702 20816 19708 20828
rect 19760 20816 19766 20868
rect 20990 20856 20996 20868
rect 20930 20828 20996 20856
rect 20990 20816 20996 20828
rect 21048 20856 21054 20868
rect 21048 20828 21680 20856
rect 21048 20816 21054 20828
rect 15059 20760 15332 20788
rect 16117 20791 16175 20797
rect 15059 20757 15071 20760
rect 15013 20751 15071 20757
rect 16117 20757 16129 20791
rect 16163 20788 16175 20791
rect 16758 20788 16764 20800
rect 16163 20760 16764 20788
rect 16163 20757 16175 20760
rect 16117 20751 16175 20757
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17313 20791 17371 20797
rect 17313 20757 17325 20791
rect 17359 20788 17371 20791
rect 17494 20788 17500 20800
rect 17359 20760 17500 20788
rect 17359 20757 17371 20760
rect 17313 20751 17371 20757
rect 17494 20748 17500 20760
rect 17552 20748 17558 20800
rect 17678 20748 17684 20800
rect 17736 20788 17742 20800
rect 18141 20791 18199 20797
rect 18141 20788 18153 20791
rect 17736 20760 18153 20788
rect 17736 20748 17742 20760
rect 18141 20757 18153 20760
rect 18187 20757 18199 20791
rect 18141 20751 18199 20757
rect 18509 20791 18567 20797
rect 18509 20757 18521 20791
rect 18555 20788 18567 20791
rect 18874 20788 18880 20800
rect 18555 20760 18880 20788
rect 18555 20757 18567 20760
rect 18509 20751 18567 20757
rect 18874 20748 18880 20760
rect 18932 20748 18938 20800
rect 21174 20748 21180 20800
rect 21232 20748 21238 20800
rect 21652 20797 21680 20828
rect 21818 20816 21824 20868
rect 21876 20856 21882 20868
rect 21876 20828 22140 20856
rect 21876 20816 21882 20828
rect 21637 20791 21695 20797
rect 21637 20757 21649 20791
rect 21683 20788 21695 20791
rect 21910 20788 21916 20800
rect 21683 20760 21916 20788
rect 21683 20757 21695 20760
rect 21637 20751 21695 20757
rect 21910 20748 21916 20760
rect 21968 20748 21974 20800
rect 22112 20797 22140 20828
rect 23566 20816 23572 20868
rect 23624 20856 23630 20868
rect 23753 20859 23811 20865
rect 23753 20856 23765 20859
rect 23624 20828 23765 20856
rect 23624 20816 23630 20828
rect 23753 20825 23765 20828
rect 23799 20825 23811 20859
rect 23753 20819 23811 20825
rect 25041 20859 25099 20865
rect 25041 20825 25053 20859
rect 25087 20856 25099 20859
rect 26234 20856 26240 20868
rect 25087 20828 26240 20856
rect 25087 20825 25099 20828
rect 25041 20819 25099 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 27338 20816 27344 20868
rect 27396 20816 27402 20868
rect 30650 20856 30656 20868
rect 27724 20828 30656 20856
rect 22097 20791 22155 20797
rect 22097 20757 22109 20791
rect 22143 20757 22155 20791
rect 22097 20751 22155 20757
rect 22462 20748 22468 20800
rect 22520 20748 22526 20800
rect 22554 20748 22560 20800
rect 22612 20748 22618 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 22704 20760 23305 20788
rect 22704 20748 22710 20760
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 23293 20751 23351 20757
rect 23658 20748 23664 20800
rect 23716 20748 23722 20800
rect 23934 20748 23940 20800
rect 23992 20788 23998 20800
rect 24673 20791 24731 20797
rect 24673 20788 24685 20791
rect 23992 20760 24685 20788
rect 23992 20748 23998 20760
rect 24673 20757 24685 20760
rect 24719 20757 24731 20791
rect 24673 20751 24731 20757
rect 25133 20791 25191 20797
rect 25133 20757 25145 20791
rect 25179 20788 25191 20791
rect 27724 20788 27752 20828
rect 30650 20816 30656 20828
rect 30708 20816 30714 20868
rect 31846 20816 31852 20868
rect 31904 20816 31910 20868
rect 25179 20760 27752 20788
rect 25179 20757 25191 20760
rect 25133 20751 25191 20757
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 31938 20748 31944 20800
rect 31996 20748 32002 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5629 20587 5687 20593
rect 5629 20553 5641 20587
rect 5675 20584 5687 20587
rect 5675 20556 6776 20584
rect 5675 20553 5687 20556
rect 5629 20547 5687 20553
rect 3878 20476 3884 20528
rect 3936 20516 3942 20528
rect 4338 20516 4344 20528
rect 3936 20488 4344 20516
rect 3936 20476 3942 20488
rect 4338 20476 4344 20488
rect 4396 20476 4402 20528
rect 6748 20516 6776 20556
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 6880 20556 11836 20584
rect 6880 20544 6886 20556
rect 6914 20516 6920 20528
rect 6748 20488 6920 20516
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 8757 20519 8815 20525
rect 8757 20485 8769 20519
rect 8803 20516 8815 20519
rect 9214 20516 9220 20528
rect 8803 20488 9220 20516
rect 8803 20485 8815 20488
rect 8757 20479 8815 20485
rect 9214 20476 9220 20488
rect 9272 20476 9278 20528
rect 9398 20476 9404 20528
rect 9456 20516 9462 20528
rect 9456 20488 10166 20516
rect 9456 20476 9462 20488
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20448 3663 20451
rect 3970 20448 3976 20460
rect 3651 20420 3976 20448
rect 3651 20417 3663 20420
rect 3605 20411 3663 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 5721 20451 5779 20457
rect 5721 20417 5733 20451
rect 5767 20448 5779 20451
rect 5767 20420 5948 20448
rect 5767 20417 5779 20420
rect 5721 20411 5779 20417
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20380 2835 20383
rect 3326 20380 3332 20392
rect 2823 20352 3332 20380
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 3326 20340 3332 20352
rect 3384 20340 3390 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5810 20340 5816 20392
rect 5868 20340 5874 20392
rect 5920 20380 5948 20420
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6144 20420 6561 20448
rect 6144 20408 6150 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 9416 20448 9444 20476
rect 11808 20457 11836 20556
rect 12406 20556 12909 20584
rect 8720 20420 9444 20448
rect 11793 20451 11851 20457
rect 8720 20408 8726 20420
rect 11793 20417 11805 20451
rect 11839 20448 11851 20451
rect 11974 20448 11980 20460
rect 11839 20420 11980 20448
rect 11839 20417 11851 20420
rect 11793 20411 11851 20417
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 6822 20380 6828 20392
rect 5920 20352 6828 20380
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7282 20340 7288 20392
rect 7340 20340 7346 20392
rect 8846 20340 8852 20392
rect 8904 20380 8910 20392
rect 9398 20380 9404 20392
rect 8904 20352 9404 20380
rect 8904 20340 8910 20352
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 10962 20380 10968 20392
rect 9723 20352 10968 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 5902 20272 5908 20324
rect 5960 20312 5966 20324
rect 8941 20315 8999 20321
rect 8941 20312 8953 20315
rect 5960 20284 8953 20312
rect 5960 20272 5966 20284
rect 8941 20281 8953 20284
rect 8987 20281 8999 20315
rect 8941 20275 8999 20281
rect 10686 20272 10692 20324
rect 10744 20312 10750 20324
rect 12406 20312 12434 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17000 20556 17509 20584
rect 17000 20544 17006 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 17497 20547 17555 20553
rect 17770 20544 17776 20596
rect 17828 20584 17834 20596
rect 18141 20587 18199 20593
rect 18141 20584 18153 20587
rect 17828 20556 18153 20584
rect 17828 20544 17834 20556
rect 18141 20553 18153 20556
rect 18187 20553 18199 20587
rect 18141 20547 18199 20553
rect 18506 20544 18512 20596
rect 18564 20544 18570 20596
rect 18874 20544 18880 20596
rect 18932 20544 18938 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19484 20556 22094 20584
rect 19484 20544 19490 20556
rect 15286 20516 15292 20528
rect 15226 20488 15292 20516
rect 15286 20476 15292 20488
rect 15344 20516 15350 20528
rect 16761 20519 16819 20525
rect 16761 20516 16773 20519
rect 15344 20488 16773 20516
rect 15344 20476 15350 20488
rect 16761 20485 16773 20488
rect 16807 20516 16819 20519
rect 17218 20516 17224 20528
rect 16807 20488 17224 20516
rect 16807 20485 16819 20488
rect 16761 20479 16819 20485
rect 17218 20476 17224 20488
rect 17276 20476 17282 20528
rect 17405 20519 17463 20525
rect 17405 20516 17417 20519
rect 17328 20488 17417 20516
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20448 13047 20451
rect 13538 20448 13544 20460
rect 13035 20420 13544 20448
rect 13035 20417 13047 20420
rect 12989 20411 13047 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 13722 20408 13728 20460
rect 13780 20408 13786 20460
rect 15378 20408 15384 20460
rect 15436 20448 15442 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15436 20420 16037 20448
rect 15436 20408 15442 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 14001 20383 14059 20389
rect 13219 20352 13860 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 10744 20284 12434 20312
rect 10744 20272 10750 20284
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 7650 20244 7656 20256
rect 5307 20216 7656 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 8389 20247 8447 20253
rect 8389 20213 8401 20247
rect 8435 20244 8447 20247
rect 8478 20244 8484 20256
rect 8435 20216 8484 20244
rect 8435 20213 8447 20216
rect 8389 20207 8447 20213
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 9030 20204 9036 20256
rect 9088 20244 9094 20256
rect 10042 20244 10048 20256
rect 9088 20216 10048 20244
rect 9088 20204 9094 20216
rect 10042 20204 10048 20216
rect 10100 20244 10106 20256
rect 10870 20244 10876 20256
rect 10100 20216 10876 20244
rect 10100 20204 10106 20216
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 11146 20204 11152 20256
rect 11204 20204 11210 20256
rect 11606 20204 11612 20256
rect 11664 20244 11670 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 11664 20216 11897 20244
rect 11664 20204 11670 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11885 20207 11943 20213
rect 12529 20247 12587 20253
rect 12529 20213 12541 20247
rect 12575 20244 12587 20247
rect 13630 20244 13636 20256
rect 12575 20216 13636 20244
rect 12575 20213 12587 20216
rect 12529 20207 12587 20213
rect 13630 20204 13636 20216
rect 13688 20204 13694 20256
rect 13832 20244 13860 20352
rect 14001 20349 14013 20383
rect 14047 20380 14059 20383
rect 14550 20380 14556 20392
rect 14047 20352 14556 20380
rect 14047 20349 14059 20352
rect 14001 20343 14059 20349
rect 14550 20340 14556 20352
rect 14608 20380 14614 20392
rect 15010 20380 15016 20392
rect 14608 20352 15016 20380
rect 14608 20340 14614 20352
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 16853 20383 16911 20389
rect 16853 20380 16865 20383
rect 15252 20352 16865 20380
rect 15252 20340 15258 20352
rect 16853 20349 16865 20352
rect 16899 20380 16911 20383
rect 17328 20380 17356 20488
rect 17405 20485 17417 20488
rect 17451 20485 17463 20519
rect 17405 20479 17463 20485
rect 19720 20457 19748 20556
rect 21910 20516 21916 20528
rect 21206 20488 21916 20516
rect 21910 20476 21916 20488
rect 21968 20476 21974 20528
rect 22066 20516 22094 20556
rect 22462 20544 22468 20596
rect 22520 20584 22526 20596
rect 23385 20587 23443 20593
rect 23385 20584 23397 20587
rect 22520 20556 23397 20584
rect 22520 20544 22526 20556
rect 23385 20553 23397 20556
rect 23431 20553 23443 20587
rect 23385 20547 23443 20553
rect 23750 20544 23756 20596
rect 23808 20584 23814 20596
rect 24029 20587 24087 20593
rect 24029 20584 24041 20587
rect 23808 20556 24041 20584
rect 23808 20544 23814 20556
rect 24029 20553 24041 20556
rect 24075 20584 24087 20587
rect 24075 20556 25912 20584
rect 24075 20553 24087 20556
rect 24029 20547 24087 20553
rect 22741 20519 22799 20525
rect 22741 20516 22753 20519
rect 22066 20488 22753 20516
rect 22741 20485 22753 20488
rect 22787 20485 22799 20519
rect 22741 20479 22799 20485
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20448 22063 20451
rect 22094 20448 22100 20460
rect 22051 20420 22100 20448
rect 22051 20417 22063 20420
rect 22005 20411 22063 20417
rect 22094 20408 22100 20420
rect 22152 20408 22158 20460
rect 23382 20408 23388 20460
rect 23440 20448 23446 20460
rect 24210 20448 24216 20460
rect 23440 20420 24216 20448
rect 23440 20408 23446 20420
rect 24210 20408 24216 20420
rect 24268 20448 24274 20460
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 24268 20420 24317 20448
rect 24268 20408 24274 20420
rect 24305 20417 24317 20420
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 25682 20408 25688 20460
rect 25740 20408 25746 20460
rect 25884 20448 25912 20556
rect 26050 20544 26056 20596
rect 26108 20584 26114 20596
rect 26513 20587 26571 20593
rect 26513 20584 26525 20587
rect 26108 20556 26525 20584
rect 26108 20544 26114 20556
rect 26513 20553 26525 20556
rect 26559 20553 26571 20587
rect 26513 20547 26571 20553
rect 26528 20516 26556 20547
rect 26602 20544 26608 20596
rect 26660 20584 26666 20596
rect 26789 20587 26847 20593
rect 26789 20584 26801 20587
rect 26660 20556 26801 20584
rect 26660 20544 26666 20556
rect 26789 20553 26801 20556
rect 26835 20584 26847 20587
rect 27522 20584 27528 20596
rect 26835 20556 27528 20584
rect 26835 20553 26847 20556
rect 26789 20547 26847 20553
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 27617 20587 27675 20593
rect 27617 20553 27629 20587
rect 27663 20584 27675 20587
rect 28994 20584 29000 20596
rect 27663 20556 29000 20584
rect 27663 20553 27675 20556
rect 27617 20547 27675 20553
rect 28994 20544 29000 20556
rect 29052 20544 29058 20596
rect 30834 20544 30840 20596
rect 30892 20584 30898 20596
rect 30929 20587 30987 20593
rect 30929 20584 30941 20587
rect 30892 20556 30941 20584
rect 30892 20544 30898 20556
rect 30929 20553 30941 20556
rect 30975 20553 30987 20587
rect 30929 20547 30987 20553
rect 27706 20516 27712 20528
rect 26528 20488 27712 20516
rect 27706 20476 27712 20488
rect 27764 20476 27770 20528
rect 30944 20516 30972 20547
rect 31754 20544 31760 20596
rect 31812 20544 31818 20596
rect 32125 20519 32183 20525
rect 32125 20516 32137 20519
rect 30944 20488 32137 20516
rect 32125 20485 32137 20488
rect 32171 20485 32183 20519
rect 32125 20479 32183 20485
rect 27246 20448 27252 20460
rect 25884 20420 27252 20448
rect 27246 20408 27252 20420
rect 27304 20408 27310 20460
rect 27525 20451 27583 20457
rect 27525 20417 27537 20451
rect 27571 20448 27583 20451
rect 27614 20448 27620 20460
rect 27571 20420 27620 20448
rect 27571 20417 27583 20420
rect 27525 20411 27583 20417
rect 27614 20408 27620 20420
rect 27672 20408 27678 20460
rect 27724 20448 27752 20476
rect 28350 20448 28356 20460
rect 27724 20420 28356 20448
rect 28350 20408 28356 20420
rect 28408 20408 28414 20460
rect 29730 20408 29736 20460
rect 29788 20408 29794 20460
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20448 31079 20451
rect 36906 20448 36912 20460
rect 31067 20420 36912 20448
rect 31067 20417 31079 20420
rect 31021 20411 31079 20417
rect 36906 20408 36912 20420
rect 36964 20408 36970 20460
rect 16899 20352 17356 20380
rect 17681 20383 17739 20389
rect 16899 20349 16911 20352
rect 16853 20343 16911 20349
rect 17681 20349 17693 20383
rect 17727 20380 17739 20383
rect 18782 20380 18788 20392
rect 17727 20352 18788 20380
rect 17727 20349 17739 20352
rect 17681 20343 17739 20349
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 18874 20340 18880 20392
rect 18932 20380 18938 20392
rect 18969 20383 19027 20389
rect 18969 20380 18981 20383
rect 18932 20352 18981 20380
rect 18932 20340 18938 20352
rect 18969 20349 18981 20352
rect 19015 20349 19027 20383
rect 18969 20343 19027 20349
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20349 19119 20383
rect 19061 20343 19119 20349
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20622 20380 20628 20392
rect 20027 20352 20628 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 15396 20284 16068 20312
rect 15396 20244 15424 20284
rect 13832 20216 15424 20244
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 16040 20244 16068 20284
rect 16114 20272 16120 20324
rect 16172 20312 16178 20324
rect 17037 20315 17095 20321
rect 17037 20312 17049 20315
rect 16172 20284 17049 20312
rect 16172 20272 16178 20284
rect 17037 20281 17049 20284
rect 17083 20281 17095 20315
rect 17037 20275 17095 20281
rect 17402 20272 17408 20324
rect 17460 20312 17466 20324
rect 19076 20312 19104 20343
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 24581 20383 24639 20389
rect 24581 20349 24593 20383
rect 24627 20380 24639 20383
rect 24670 20380 24676 20392
rect 24627 20352 24676 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 24670 20340 24676 20352
rect 24728 20340 24734 20392
rect 25958 20340 25964 20392
rect 26016 20380 26022 20392
rect 26053 20383 26111 20389
rect 26053 20380 26065 20383
rect 26016 20352 26065 20380
rect 26016 20340 26022 20352
rect 26053 20349 26065 20352
rect 26099 20380 26111 20383
rect 27709 20383 27767 20389
rect 26099 20352 27292 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 17460 20284 19104 20312
rect 17460 20272 17466 20284
rect 16574 20244 16580 20256
rect 16040 20216 16580 20244
rect 16574 20204 16580 20216
rect 16632 20204 16638 20256
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 18874 20244 18880 20256
rect 17184 20216 18880 20244
rect 17184 20204 17190 20216
rect 18874 20204 18880 20216
rect 18932 20204 18938 20256
rect 19076 20244 19104 20284
rect 22554 20272 22560 20324
rect 22612 20312 22618 20324
rect 27157 20315 27215 20321
rect 27157 20312 27169 20315
rect 22612 20284 24440 20312
rect 22612 20272 22618 20284
rect 21453 20247 21511 20253
rect 21453 20244 21465 20247
rect 19076 20216 21465 20244
rect 21453 20213 21465 20216
rect 21499 20213 21511 20247
rect 21453 20207 21511 20213
rect 21818 20204 21824 20256
rect 21876 20244 21882 20256
rect 22186 20244 22192 20256
rect 21876 20216 22192 20244
rect 21876 20204 21882 20216
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 24412 20244 24440 20284
rect 25608 20284 27169 20312
rect 25608 20244 25636 20284
rect 27157 20281 27169 20284
rect 27203 20281 27215 20315
rect 27264 20312 27292 20352
rect 27709 20349 27721 20383
rect 27755 20349 27767 20383
rect 27709 20343 27767 20349
rect 28629 20383 28687 20389
rect 28629 20349 28641 20383
rect 28675 20380 28687 20383
rect 30190 20380 30196 20392
rect 28675 20352 30196 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 27724 20312 27752 20343
rect 30190 20340 30196 20352
rect 30248 20340 30254 20392
rect 30282 20340 30288 20392
rect 30340 20380 30346 20392
rect 31113 20383 31171 20389
rect 31113 20380 31125 20383
rect 30340 20352 31125 20380
rect 30340 20340 30346 20352
rect 31113 20349 31125 20352
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 27264 20284 27752 20312
rect 27157 20275 27215 20281
rect 29638 20272 29644 20324
rect 29696 20312 29702 20324
rect 31573 20315 31631 20321
rect 31573 20312 31585 20315
rect 29696 20284 31585 20312
rect 29696 20272 29702 20284
rect 31573 20281 31585 20284
rect 31619 20281 31631 20315
rect 31573 20275 31631 20281
rect 24412 20216 25636 20244
rect 25682 20204 25688 20256
rect 25740 20244 25746 20256
rect 26421 20247 26479 20253
rect 26421 20244 26433 20247
rect 25740 20216 26433 20244
rect 25740 20204 25746 20216
rect 26421 20213 26433 20216
rect 26467 20244 26479 20247
rect 27246 20244 27252 20256
rect 26467 20216 27252 20244
rect 26467 20213 26479 20216
rect 26421 20207 26479 20213
rect 27246 20204 27252 20216
rect 27304 20204 27310 20256
rect 28810 20204 28816 20256
rect 28868 20244 28874 20256
rect 30101 20247 30159 20253
rect 30101 20244 30113 20247
rect 28868 20216 30113 20244
rect 28868 20204 28874 20216
rect 30101 20213 30113 20216
rect 30147 20213 30159 20247
rect 30101 20207 30159 20213
rect 30190 20204 30196 20256
rect 30248 20244 30254 20256
rect 30561 20247 30619 20253
rect 30561 20244 30573 20247
rect 30248 20216 30573 20244
rect 30248 20204 30254 20216
rect 30561 20213 30573 20216
rect 30607 20213 30619 20247
rect 30561 20207 30619 20213
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 5442 20040 5448 20052
rect 4540 20012 5448 20040
rect 4540 19913 4568 20012
rect 5442 20000 5448 20012
rect 5500 20040 5506 20052
rect 8846 20040 8852 20052
rect 5500 20012 8852 20040
rect 5500 20000 5506 20012
rect 6270 19932 6276 19984
rect 6328 19932 6334 19984
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19873 4583 19907
rect 4525 19867 4583 19873
rect 6733 19907 6791 19913
rect 6733 19873 6745 19907
rect 6779 19904 6791 19907
rect 6840 19904 6868 20012
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 9490 20000 9496 20052
rect 9548 20040 9554 20052
rect 10778 20040 10784 20052
rect 9548 20012 10784 20040
rect 9548 20000 9554 20012
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11256 20012 11744 20040
rect 11256 19972 11284 20012
rect 10796 19944 11284 19972
rect 11716 19972 11744 20012
rect 11790 20000 11796 20052
rect 11848 20000 11854 20052
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 12124 20012 14197 20040
rect 12124 20000 12130 20012
rect 14185 20009 14197 20012
rect 14231 20040 14243 20043
rect 17126 20040 17132 20052
rect 14231 20012 17132 20040
rect 14231 20009 14243 20012
rect 14185 20003 14243 20009
rect 17126 20000 17132 20012
rect 17184 20000 17190 20052
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19334 20040 19340 20052
rect 18739 20012 19340 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19576 20012 19717 20040
rect 19576 20000 19582 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 49234 20040 49240 20052
rect 19705 20003 19763 20009
rect 22066 20012 49240 20040
rect 13538 19972 13544 19984
rect 11716 19944 13544 19972
rect 6779 19876 6868 19904
rect 7009 19907 7067 19913
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 7009 19873 7021 19907
rect 7055 19904 7067 19907
rect 9030 19904 9036 19916
rect 7055 19876 9036 19904
rect 7055 19873 7067 19876
rect 7009 19867 7067 19873
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 10796 19904 10824 19944
rect 13538 19932 13544 19944
rect 13596 19972 13602 19984
rect 13722 19972 13728 19984
rect 13596 19944 13728 19972
rect 13596 19932 13602 19944
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 14090 19932 14096 19984
rect 14148 19972 14154 19984
rect 14550 19972 14556 19984
rect 14148 19944 14556 19972
rect 14148 19932 14154 19944
rect 14550 19932 14556 19944
rect 14608 19932 14614 19984
rect 16945 19975 17003 19981
rect 16945 19941 16957 19975
rect 16991 19972 17003 19975
rect 16991 19944 17816 19972
rect 16991 19941 17003 19944
rect 16945 19935 17003 19941
rect 9171 19876 10824 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 10870 19864 10876 19916
rect 10928 19864 10934 19916
rect 12345 19907 12403 19913
rect 12345 19873 12357 19907
rect 12391 19904 12403 19907
rect 13354 19904 13360 19916
rect 12391 19876 13360 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 13679 19876 14841 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14829 19873 14841 19876
rect 14875 19904 14887 19907
rect 15470 19904 15476 19916
rect 14875 19876 15476 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 16761 19907 16819 19913
rect 16761 19873 16773 19907
rect 16807 19904 16819 19907
rect 17494 19904 17500 19916
rect 16807 19876 17500 19904
rect 16807 19873 16819 19876
rect 16761 19867 16819 19873
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17678 19864 17684 19916
rect 17736 19864 17742 19916
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 4430 19836 4436 19848
rect 1811 19808 4436 19836
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 10778 19796 10784 19848
rect 10836 19836 10842 19848
rect 12253 19839 12311 19845
rect 10836 19808 11376 19836
rect 10836 19796 10842 19808
rect 2777 19771 2835 19777
rect 2777 19737 2789 19771
rect 2823 19768 2835 19771
rect 2866 19768 2872 19780
rect 2823 19740 2872 19768
rect 2823 19737 2835 19740
rect 2777 19731 2835 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 3605 19771 3663 19777
rect 3605 19737 3617 19771
rect 3651 19768 3663 19771
rect 4522 19768 4528 19780
rect 3651 19740 4528 19768
rect 3651 19737 3663 19740
rect 3605 19731 3663 19737
rect 4522 19728 4528 19740
rect 4580 19728 4586 19780
rect 4798 19728 4804 19780
rect 4856 19728 4862 19780
rect 6270 19768 6276 19780
rect 6026 19740 6276 19768
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 3881 19703 3939 19709
rect 3881 19700 3893 19703
rect 3467 19672 3893 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 3881 19669 3893 19672
rect 3927 19700 3939 19703
rect 4065 19703 4123 19709
rect 4065 19700 4077 19703
rect 3927 19672 4077 19700
rect 3927 19669 3939 19672
rect 3881 19663 3939 19669
rect 4065 19669 4077 19672
rect 4111 19700 4123 19703
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 4111 19672 4261 19700
rect 4111 19669 4123 19672
rect 4065 19663 4123 19669
rect 4249 19669 4261 19672
rect 4295 19700 4307 19703
rect 6104 19700 6132 19740
rect 6270 19728 6276 19740
rect 6328 19768 6334 19780
rect 8662 19768 8668 19780
rect 6328 19740 7498 19768
rect 8312 19740 8668 19768
rect 6328 19728 6334 19740
rect 4295 19672 6132 19700
rect 7392 19700 7420 19740
rect 8312 19712 8340 19740
rect 8662 19728 8668 19740
rect 8720 19728 8726 19780
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 9324 19740 9413 19768
rect 8294 19700 8300 19712
rect 7392 19672 8300 19700
rect 4295 19669 4307 19672
rect 4249 19663 4307 19669
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8846 19700 8852 19712
rect 8527 19672 8852 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9324 19700 9352 19740
rect 9401 19737 9413 19740
rect 9447 19737 9459 19771
rect 9401 19731 9459 19737
rect 9490 19728 9496 19780
rect 9548 19768 9554 19780
rect 9548 19740 9890 19768
rect 9548 19728 9554 19740
rect 11054 19728 11060 19780
rect 11112 19768 11118 19780
rect 11348 19777 11376 19808
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 14458 19836 14464 19848
rect 12299 19808 14464 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 17788 19836 17816 19944
rect 21542 19932 21548 19984
rect 21600 19972 21606 19984
rect 22066 19972 22094 20012
rect 49234 20000 49240 20012
rect 49292 20000 49298 20052
rect 21600 19944 22094 19972
rect 21600 19932 21606 19944
rect 22738 19932 22744 19984
rect 22796 19972 22802 19984
rect 27617 19975 27675 19981
rect 22796 19944 25084 19972
rect 22796 19932 22802 19944
rect 17865 19907 17923 19913
rect 17865 19873 17877 19907
rect 17911 19904 17923 19907
rect 17911 19876 18736 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 17788 19808 18552 19836
rect 11333 19771 11391 19777
rect 11112 19740 11284 19768
rect 11112 19728 11118 19740
rect 11146 19700 11152 19712
rect 9324 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11256 19700 11284 19740
rect 11333 19737 11345 19771
rect 11379 19768 11391 19771
rect 11517 19771 11575 19777
rect 11517 19768 11529 19771
rect 11379 19740 11529 19768
rect 11379 19737 11391 19740
rect 11333 19731 11391 19737
rect 11517 19737 11529 19740
rect 11563 19768 11575 19771
rect 13262 19768 13268 19780
rect 11563 19740 13268 19768
rect 11563 19737 11575 19740
rect 11517 19731 11575 19737
rect 13262 19728 13268 19740
rect 13320 19728 13326 19780
rect 13449 19771 13507 19777
rect 13449 19737 13461 19771
rect 13495 19768 13507 19771
rect 13495 19740 15240 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 12161 19703 12219 19709
rect 12161 19700 12173 19703
rect 11256 19672 12173 19700
rect 12161 19669 12173 19672
rect 12207 19669 12219 19703
rect 12161 19663 12219 19669
rect 12986 19660 12992 19712
rect 13044 19660 13050 19712
rect 13354 19660 13360 19712
rect 13412 19660 13418 19712
rect 13906 19660 13912 19712
rect 13964 19700 13970 19712
rect 14642 19700 14648 19712
rect 13964 19672 14648 19700
rect 13964 19660 13970 19672
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 15212 19700 15240 19740
rect 15286 19728 15292 19780
rect 15344 19728 15350 19780
rect 18322 19768 18328 19780
rect 16224 19740 18328 19768
rect 16224 19700 16252 19740
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 15212 19672 16252 19700
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 16390 19700 16396 19712
rect 16347 19672 16396 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 17586 19660 17592 19712
rect 17644 19660 17650 19712
rect 17678 19660 17684 19712
rect 17736 19700 17742 19712
rect 17862 19700 17868 19712
rect 17736 19672 17868 19700
rect 17736 19660 17742 19672
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 18414 19660 18420 19712
rect 18472 19660 18478 19712
rect 18524 19700 18552 19808
rect 18708 19768 18736 19876
rect 18782 19864 18788 19916
rect 18840 19904 18846 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 18840 19876 20545 19904
rect 18840 19864 18846 19876
rect 20533 19873 20545 19876
rect 20579 19904 20591 19907
rect 21174 19904 21180 19916
rect 20579 19876 21180 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 22005 19907 22063 19913
rect 22005 19904 22017 19907
rect 21560 19876 22017 19904
rect 21560 19848 21588 19876
rect 22005 19873 22017 19876
rect 22051 19904 22063 19907
rect 23842 19904 23848 19916
rect 22051 19876 23848 19904
rect 22051 19873 22063 19876
rect 22005 19867 22063 19873
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19058 19836 19064 19848
rect 18923 19808 19064 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19702 19796 19708 19848
rect 19760 19836 19766 19848
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 19760 19808 20269 19836
rect 19760 19796 19766 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 21542 19796 21548 19848
rect 21600 19796 21606 19848
rect 22278 19796 22284 19848
rect 22336 19836 22342 19848
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22336 19808 22569 19836
rect 22336 19796 22342 19808
rect 22557 19805 22569 19808
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 23750 19796 23756 19848
rect 23808 19796 23814 19848
rect 25056 19836 25084 19944
rect 27617 19941 27629 19975
rect 27663 19972 27675 19975
rect 27798 19972 27804 19984
rect 27663 19944 27804 19972
rect 27663 19941 27675 19944
rect 27617 19935 27675 19941
rect 27798 19932 27804 19944
rect 27856 19932 27862 19984
rect 29733 19975 29791 19981
rect 29733 19941 29745 19975
rect 29779 19972 29791 19975
rect 29779 19944 31432 19972
rect 29779 19941 29791 19944
rect 29733 19935 29791 19941
rect 25317 19907 25375 19913
rect 25317 19873 25329 19907
rect 25363 19904 25375 19907
rect 26142 19904 26148 19916
rect 25363 19876 26148 19904
rect 25363 19873 25375 19876
rect 25317 19867 25375 19873
rect 26142 19864 26148 19876
rect 26200 19864 26206 19916
rect 28626 19864 28632 19916
rect 28684 19864 28690 19916
rect 28994 19864 29000 19916
rect 29052 19904 29058 19916
rect 31297 19907 31355 19913
rect 31297 19904 31309 19907
rect 29052 19876 31309 19904
rect 29052 19864 29058 19876
rect 31297 19873 31309 19876
rect 31343 19873 31355 19907
rect 31404 19904 31432 19944
rect 31754 19932 31760 19984
rect 31812 19972 31818 19984
rect 46934 19972 46940 19984
rect 31812 19944 46940 19972
rect 31812 19932 31818 19944
rect 46934 19932 46940 19944
rect 46992 19932 46998 19984
rect 32030 19904 32036 19916
rect 31404 19876 32036 19904
rect 31297 19867 31355 19873
rect 32030 19864 32036 19876
rect 32088 19864 32094 19916
rect 25056 19808 25728 19836
rect 18966 19768 18972 19780
rect 18708 19740 18972 19768
rect 18966 19728 18972 19740
rect 19024 19768 19030 19780
rect 19334 19768 19340 19780
rect 19024 19740 19340 19768
rect 19024 19728 19030 19740
rect 19334 19728 19340 19740
rect 19392 19728 19398 19780
rect 19613 19771 19671 19777
rect 19613 19737 19625 19771
rect 19659 19768 19671 19771
rect 19886 19768 19892 19780
rect 19659 19740 19892 19768
rect 19659 19737 19671 19740
rect 19613 19731 19671 19737
rect 19628 19700 19656 19731
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 21910 19768 21916 19780
rect 21758 19740 21916 19768
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 22738 19728 22744 19780
rect 22796 19728 22802 19780
rect 25041 19771 25099 19777
rect 25041 19737 25053 19771
rect 25087 19768 25099 19771
rect 25590 19768 25596 19780
rect 25087 19740 25596 19768
rect 25087 19737 25099 19740
rect 25041 19731 25099 19737
rect 25590 19728 25596 19740
rect 25648 19728 25654 19780
rect 25700 19768 25728 19808
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25832 19808 25881 19836
rect 25832 19796 25838 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 27246 19796 27252 19848
rect 27304 19836 27310 19848
rect 27982 19836 27988 19848
rect 27304 19808 27988 19836
rect 27304 19796 27310 19808
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 28353 19839 28411 19845
rect 28353 19805 28365 19839
rect 28399 19836 28411 19839
rect 28442 19836 28448 19848
rect 28399 19808 28448 19836
rect 28399 19805 28411 19808
rect 28353 19799 28411 19805
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 29914 19796 29920 19848
rect 29972 19836 29978 19848
rect 30193 19839 30251 19845
rect 30193 19836 30205 19839
rect 29972 19808 30205 19836
rect 29972 19796 29978 19808
rect 30193 19805 30205 19808
rect 30239 19805 30251 19839
rect 30193 19799 30251 19805
rect 30374 19796 30380 19848
rect 30432 19836 30438 19848
rect 31113 19839 31171 19845
rect 31113 19836 31125 19839
rect 30432 19808 31125 19836
rect 30432 19796 30438 19808
rect 31113 19805 31125 19808
rect 31159 19836 31171 19839
rect 31662 19836 31668 19848
rect 31159 19808 31668 19836
rect 31159 19805 31171 19808
rect 31113 19799 31171 19805
rect 31662 19796 31668 19808
rect 31720 19796 31726 19848
rect 26145 19771 26203 19777
rect 26145 19768 26157 19771
rect 25700 19740 26157 19768
rect 26145 19737 26157 19740
rect 26191 19768 26203 19771
rect 26418 19768 26424 19780
rect 26191 19740 26424 19768
rect 26191 19737 26203 19740
rect 26145 19731 26203 19737
rect 26418 19728 26424 19740
rect 26476 19728 26482 19780
rect 27908 19740 30788 19768
rect 18524 19672 19656 19700
rect 23290 19660 23296 19712
rect 23348 19660 23354 19712
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 24673 19703 24731 19709
rect 24673 19700 24685 19703
rect 23808 19672 24685 19700
rect 23808 19660 23814 19672
rect 24673 19669 24685 19672
rect 24719 19669 24731 19703
rect 24673 19663 24731 19669
rect 25133 19703 25191 19709
rect 25133 19669 25145 19703
rect 25179 19700 25191 19703
rect 27908 19700 27936 19740
rect 25179 19672 27936 19700
rect 25179 19669 25191 19672
rect 25133 19663 25191 19669
rect 27982 19660 27988 19712
rect 28040 19700 28046 19712
rect 29730 19700 29736 19712
rect 28040 19672 29736 19700
rect 28040 19660 28046 19672
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 30374 19660 30380 19712
rect 30432 19660 30438 19712
rect 30760 19709 30788 19740
rect 30745 19703 30803 19709
rect 30745 19669 30757 19703
rect 30791 19669 30803 19703
rect 30745 19663 30803 19669
rect 31205 19703 31263 19709
rect 31205 19669 31217 19703
rect 31251 19700 31263 19703
rect 37182 19700 37188 19712
rect 31251 19672 37188 19700
rect 31251 19669 31263 19672
rect 31205 19663 31263 19669
rect 37182 19660 37188 19672
rect 37240 19660 37246 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 5258 19456 5264 19508
rect 5316 19456 5322 19508
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 6730 19496 6736 19508
rect 5767 19468 6736 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 6730 19456 6736 19468
rect 6788 19456 6794 19508
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 10686 19496 10692 19508
rect 7616 19468 10692 19496
rect 7616 19456 7622 19468
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 10873 19499 10931 19505
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 11882 19496 11888 19508
rect 10919 19468 11888 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 14090 19496 14096 19508
rect 11992 19468 14096 19496
rect 11992 19440 12020 19468
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 14369 19499 14427 19505
rect 14369 19465 14381 19499
rect 14415 19465 14427 19499
rect 14369 19459 14427 19465
rect 4154 19388 4160 19440
rect 4212 19428 4218 19440
rect 4341 19431 4399 19437
rect 4341 19428 4353 19431
rect 4212 19400 4353 19428
rect 4212 19388 4218 19400
rect 4341 19397 4353 19400
rect 4387 19397 4399 19431
rect 4341 19391 4399 19397
rect 5629 19431 5687 19437
rect 5629 19397 5641 19431
rect 5675 19428 5687 19431
rect 5675 19400 9076 19428
rect 5675 19397 5687 19400
rect 5629 19391 5687 19397
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19360 1823 19363
rect 2130 19360 2136 19372
rect 1811 19332 2136 19360
rect 1811 19329 1823 19332
rect 1765 19323 1823 19329
rect 2130 19320 2136 19332
rect 2188 19320 2194 19372
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 3602 19320 3608 19372
rect 3660 19320 3666 19372
rect 6641 19363 6699 19369
rect 6641 19329 6653 19363
rect 6687 19334 6699 19363
rect 6687 19329 6776 19334
rect 6641 19323 6776 19329
rect 6656 19306 6776 19323
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 8662 19360 8668 19372
rect 8619 19332 8668 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 9048 19360 9076 19400
rect 9122 19388 9128 19440
rect 9180 19428 9186 19440
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 9180 19400 9321 19428
rect 9180 19388 9186 19400
rect 9309 19397 9321 19400
rect 9355 19397 9367 19431
rect 11422 19428 11428 19440
rect 9309 19391 9367 19397
rect 10428 19400 11428 19428
rect 10318 19360 10324 19372
rect 9048 19332 10324 19360
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 4246 19252 4252 19304
rect 4304 19292 4310 19304
rect 5813 19295 5871 19301
rect 5813 19292 5825 19295
rect 4304 19264 5825 19292
rect 4304 19252 4310 19264
rect 5813 19261 5825 19264
rect 5859 19292 5871 19295
rect 6546 19292 6552 19304
rect 5859 19264 6552 19292
rect 5859 19261 5871 19264
rect 5813 19255 5871 19261
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 4982 19184 4988 19236
rect 5040 19224 5046 19236
rect 5350 19224 5356 19236
rect 5040 19196 5356 19224
rect 5040 19184 5046 19196
rect 5350 19184 5356 19196
rect 5408 19184 5414 19236
rect 5442 19184 5448 19236
rect 5500 19224 5506 19236
rect 6748 19224 6776 19306
rect 10134 19252 10140 19304
rect 10192 19252 10198 19304
rect 5500 19196 6776 19224
rect 5500 19184 5506 19196
rect 6914 19184 6920 19236
rect 6972 19224 6978 19236
rect 10226 19224 10232 19236
rect 6972 19196 10232 19224
rect 6972 19184 6978 19196
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 10428 19233 10456 19400
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 11974 19428 11980 19440
rect 11716 19400 11980 19428
rect 10778 19320 10784 19372
rect 10836 19320 10842 19372
rect 11606 19360 11612 19372
rect 11348 19332 11612 19360
rect 10962 19252 10968 19304
rect 11020 19252 11026 19304
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11348 19292 11376 19332
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 11716 19369 11744 19400
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 13262 19428 13268 19440
rect 13202 19400 13268 19428
rect 13262 19388 13268 19400
rect 13320 19428 13326 19440
rect 13814 19428 13820 19440
rect 13320 19400 13820 19428
rect 13320 19388 13326 19400
rect 13814 19388 13820 19400
rect 13872 19388 13878 19440
rect 13906 19388 13912 19440
rect 13964 19388 13970 19440
rect 14384 19428 14412 19459
rect 14642 19456 14648 19508
rect 14700 19496 14706 19508
rect 14829 19499 14887 19505
rect 14829 19496 14841 19499
rect 14700 19468 14841 19496
rect 14700 19456 14706 19468
rect 14829 19465 14841 19468
rect 14875 19465 14887 19499
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 14829 19459 14887 19465
rect 15120 19468 17877 19496
rect 14292 19400 14412 19428
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 14292 19360 14320 19400
rect 14458 19388 14464 19440
rect 14516 19428 14522 19440
rect 15120 19428 15148 19468
rect 17865 19465 17877 19468
rect 17911 19465 17923 19499
rect 17865 19459 17923 19465
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 18012 19468 18337 19496
rect 18012 19456 18018 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 18325 19459 18383 19465
rect 19058 19456 19064 19508
rect 19116 19456 19122 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 19392 19468 21465 19496
rect 19392 19456 19398 19468
rect 21453 19465 21465 19468
rect 21499 19465 21511 19499
rect 21453 19459 21511 19465
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 23290 19496 23296 19508
rect 22419 19468 23296 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 25682 19496 25688 19508
rect 23400 19468 25688 19496
rect 14516 19400 15148 19428
rect 16761 19431 16819 19437
rect 14516 19388 14522 19400
rect 16761 19397 16773 19431
rect 16807 19428 16819 19431
rect 17126 19428 17132 19440
rect 16807 19400 17132 19428
rect 16807 19397 16819 19400
rect 16761 19391 16819 19397
rect 17126 19388 17132 19400
rect 17184 19388 17190 19440
rect 19426 19428 19432 19440
rect 17236 19400 19432 19428
rect 13504 19332 14320 19360
rect 13504 19320 13510 19332
rect 14550 19320 14556 19372
rect 14608 19360 14614 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14608 19332 14749 19360
rect 14608 19320 14614 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 15286 19360 15292 19372
rect 14737 19323 14795 19329
rect 14844 19332 15292 19360
rect 11112 19264 11376 19292
rect 11977 19295 12035 19301
rect 11112 19252 11118 19264
rect 11977 19261 11989 19295
rect 12023 19292 12035 19295
rect 13722 19292 13728 19304
rect 12023 19264 13728 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 14844 19292 14872 19332
rect 15286 19320 15292 19332
rect 15344 19320 15350 19372
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 14016 19264 14872 19292
rect 10413 19227 10471 19233
rect 10413 19193 10425 19227
rect 10459 19193 10471 19227
rect 10413 19187 10471 19193
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 6086 19156 6092 19168
rect 4672 19128 6092 19156
rect 4672 19116 4678 19128
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 8478 19156 8484 19168
rect 6512 19128 8484 19156
rect 6512 19116 6518 19128
rect 8478 19116 8484 19128
rect 8536 19156 8542 19168
rect 9490 19156 9496 19168
rect 8536 19128 9496 19156
rect 8536 19116 8542 19128
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 10321 19159 10379 19165
rect 10321 19125 10333 19159
rect 10367 19156 10379 19159
rect 10778 19156 10784 19168
rect 10367 19128 10784 19156
rect 10367 19125 10379 19128
rect 10321 19119 10379 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 10980 19156 11008 19252
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 10980 19128 13461 19156
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14016 19165 14044 19264
rect 14918 19252 14924 19304
rect 14976 19252 14982 19304
rect 16942 19252 16948 19304
rect 17000 19252 17006 19304
rect 17236 19233 17264 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 22465 19431 22523 19437
rect 22465 19397 22477 19431
rect 22511 19428 22523 19431
rect 22646 19428 22652 19440
rect 22511 19400 22652 19428
rect 22511 19397 22523 19400
rect 22465 19391 22523 19397
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 23400 19428 23428 19468
rect 25682 19456 25688 19468
rect 25740 19456 25746 19508
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 26421 19499 26479 19505
rect 26421 19496 26433 19499
rect 26292 19468 26433 19496
rect 26292 19456 26298 19468
rect 26421 19465 26433 19468
rect 26467 19465 26479 19499
rect 26421 19459 26479 19465
rect 26786 19456 26792 19508
rect 26844 19496 26850 19508
rect 27246 19496 27252 19508
rect 26844 19468 27252 19496
rect 26844 19456 26850 19468
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 27706 19456 27712 19508
rect 27764 19456 27770 19508
rect 27798 19456 27804 19508
rect 27856 19496 27862 19508
rect 30374 19496 30380 19508
rect 27856 19468 30380 19496
rect 27856 19456 27862 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 30469 19499 30527 19505
rect 30469 19465 30481 19499
rect 30515 19496 30527 19499
rect 32122 19496 32128 19508
rect 30515 19468 32128 19496
rect 30515 19465 30527 19468
rect 30469 19459 30527 19465
rect 32122 19456 32128 19468
rect 32180 19456 32186 19508
rect 22756 19400 23428 19428
rect 17413 19363 17471 19369
rect 17413 19329 17425 19363
rect 17459 19360 17471 19363
rect 17678 19360 17684 19372
rect 17459 19332 17684 19360
rect 17459 19329 17471 19332
rect 17413 19323 17471 19329
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18233 19363 18291 19369
rect 18233 19360 18245 19363
rect 17828 19332 18245 19360
rect 17828 19320 17834 19332
rect 18233 19329 18245 19332
rect 18279 19360 18291 19363
rect 18506 19360 18512 19372
rect 18279 19332 18512 19360
rect 18279 19329 18291 19332
rect 18233 19323 18291 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 19116 19332 19257 19360
rect 19116 19320 19122 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 21910 19360 21916 19372
rect 21114 19332 21916 19360
rect 19245 19323 19303 19329
rect 21910 19320 21916 19332
rect 21968 19360 21974 19372
rect 22756 19360 22784 19400
rect 25314 19388 25320 19440
rect 25372 19428 25378 19440
rect 28537 19431 28595 19437
rect 28537 19428 28549 19431
rect 25372 19400 28549 19428
rect 25372 19388 25378 19400
rect 28537 19397 28549 19400
rect 28583 19428 28595 19431
rect 28810 19428 28816 19440
rect 28583 19400 28816 19428
rect 28583 19397 28595 19400
rect 28537 19391 28595 19397
rect 28810 19388 28816 19400
rect 28868 19388 28874 19440
rect 21968 19332 22784 19360
rect 21968 19320 21974 19332
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 17368 19264 18429 19292
rect 17368 19252 17374 19264
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19812 19264 19993 19292
rect 17221 19227 17279 19233
rect 17221 19193 17233 19227
rect 17267 19193 17279 19227
rect 17221 19187 17279 19193
rect 17678 19184 17684 19236
rect 17736 19224 17742 19236
rect 19720 19224 19748 19252
rect 17736 19196 19748 19224
rect 17736 19184 17742 19196
rect 14001 19159 14059 19165
rect 14001 19156 14013 19159
rect 13872 19128 14013 19156
rect 13872 19116 13878 19128
rect 14001 19125 14013 19128
rect 14047 19125 14059 19159
rect 14001 19119 14059 19125
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 15749 19159 15807 19165
rect 15749 19156 15761 19159
rect 14516 19128 15761 19156
rect 14516 19116 14522 19128
rect 15749 19125 15761 19128
rect 15795 19125 15807 19159
rect 15749 19119 15807 19125
rect 16022 19116 16028 19168
rect 16080 19156 16086 19168
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 16080 19128 16221 19156
rect 16080 19116 16086 19128
rect 16209 19125 16221 19128
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 16485 19159 16543 19165
rect 16485 19125 16497 19159
rect 16531 19156 16543 19159
rect 17770 19156 17776 19168
rect 16531 19128 17776 19156
rect 16531 19125 16543 19128
rect 16485 19119 16543 19125
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18690 19116 18696 19168
rect 18748 19156 18754 19168
rect 19812 19156 19840 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 22554 19292 22560 19304
rect 20680 19264 22560 19292
rect 20680 19252 20686 19264
rect 22554 19252 22560 19264
rect 22612 19252 22618 19304
rect 22664 19292 22692 19332
rect 22830 19320 22836 19372
rect 22888 19360 22894 19372
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 22888 19332 24041 19360
rect 22888 19320 22894 19332
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 24121 19363 24179 19369
rect 24121 19329 24133 19363
rect 24167 19360 24179 19363
rect 24486 19360 24492 19372
rect 24167 19332 24492 19360
rect 24167 19329 24179 19332
rect 24121 19323 24179 19329
rect 24486 19320 24492 19332
rect 24544 19320 24550 19372
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19360 25007 19363
rect 25038 19360 25044 19372
rect 24995 19332 25044 19360
rect 24995 19329 25007 19332
rect 24949 19323 25007 19329
rect 23017 19295 23075 19301
rect 23017 19292 23029 19295
rect 22664 19264 23029 19292
rect 23017 19261 23029 19264
rect 23063 19261 23075 19295
rect 23017 19255 23075 19261
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24854 19292 24860 19304
rect 24351 19264 24860 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 22002 19184 22008 19236
rect 22060 19184 22066 19236
rect 22094 19184 22100 19236
rect 22152 19224 22158 19236
rect 23385 19227 23443 19233
rect 23385 19224 23397 19227
rect 22152 19196 23397 19224
rect 22152 19184 22158 19196
rect 23385 19193 23397 19196
rect 23431 19224 23443 19227
rect 24964 19224 24992 19323
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 29638 19320 29644 19372
rect 29696 19320 29702 19372
rect 30650 19320 30656 19372
rect 30708 19360 30714 19372
rect 31113 19363 31171 19369
rect 31113 19360 31125 19363
rect 30708 19332 31125 19360
rect 30708 19320 30714 19332
rect 31113 19329 31125 19332
rect 31159 19329 31171 19363
rect 31846 19360 31852 19372
rect 31113 19323 31171 19329
rect 31772 19332 31852 19360
rect 25774 19252 25780 19304
rect 25832 19252 25838 19304
rect 26878 19252 26884 19304
rect 26936 19292 26942 19304
rect 26973 19295 27031 19301
rect 26973 19292 26985 19295
rect 26936 19264 26985 19292
rect 26936 19252 26942 19264
rect 26973 19261 26985 19264
rect 27019 19261 27031 19295
rect 26973 19255 27031 19261
rect 27430 19252 27436 19304
rect 27488 19252 27494 19304
rect 28258 19252 28264 19304
rect 28316 19252 28322 19304
rect 30926 19292 30932 19304
rect 28368 19264 30932 19292
rect 28368 19224 28396 19264
rect 30926 19252 30932 19264
rect 30984 19252 30990 19304
rect 31021 19295 31079 19301
rect 31021 19261 31033 19295
rect 31067 19292 31079 19295
rect 31772 19292 31800 19332
rect 31846 19320 31852 19332
rect 31904 19320 31910 19372
rect 31067 19264 31800 19292
rect 31067 19261 31079 19264
rect 31021 19255 31079 19261
rect 23431 19196 24992 19224
rect 25424 19196 28396 19224
rect 23431 19193 23443 19196
rect 23385 19187 23443 19193
rect 23474 19156 23480 19168
rect 18748 19128 23480 19156
rect 18748 19116 18754 19128
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 23566 19116 23572 19168
rect 23624 19156 23630 19168
rect 23661 19159 23719 19165
rect 23661 19156 23673 19159
rect 23624 19128 23673 19156
rect 23624 19116 23630 19128
rect 23661 19125 23673 19128
rect 23707 19125 23719 19159
rect 23661 19119 23719 19125
rect 24118 19116 24124 19168
rect 24176 19156 24182 19168
rect 25424 19156 25452 19196
rect 24176 19128 25452 19156
rect 24176 19116 24182 19128
rect 27798 19116 27804 19168
rect 27856 19156 27862 19168
rect 27893 19159 27951 19165
rect 27893 19156 27905 19159
rect 27856 19128 27905 19156
rect 27856 19116 27862 19128
rect 27893 19125 27905 19128
rect 27939 19125 27951 19159
rect 27893 19119 27951 19125
rect 28626 19116 28632 19168
rect 28684 19156 28690 19168
rect 30009 19159 30067 19165
rect 30009 19156 30021 19159
rect 28684 19128 30021 19156
rect 28684 19116 28690 19128
rect 30009 19125 30021 19128
rect 30055 19156 30067 19159
rect 30282 19156 30288 19168
rect 30055 19128 30288 19156
rect 30055 19125 30067 19128
rect 30009 19119 30067 19125
rect 30282 19116 30288 19128
rect 30340 19116 30346 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 15010 18952 15016 18964
rect 3927 18924 15016 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 3988 18825 4016 18924
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 22002 18952 22008 18964
rect 15120 18924 22008 18952
rect 8570 18844 8576 18896
rect 8628 18844 8634 18896
rect 9646 18856 9812 18884
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1452 18788 2053 18816
rect 1452 18776 1458 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 3973 18819 4031 18825
rect 3973 18785 3985 18819
rect 4019 18785 4031 18819
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 3973 18779 4031 18785
rect 4632 18788 6837 18816
rect 4632 18760 4660 18788
rect 6825 18785 6837 18788
rect 6871 18816 6883 18819
rect 8478 18816 8484 18828
rect 6871 18788 8484 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 4522 18748 4528 18760
rect 1811 18720 4528 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 8202 18708 8208 18760
rect 8260 18708 8266 18760
rect 8588 18748 8616 18844
rect 9122 18776 9128 18828
rect 9180 18816 9186 18828
rect 9646 18816 9674 18856
rect 9180 18788 9674 18816
rect 9180 18776 9186 18788
rect 9784 18757 9812 18856
rect 9858 18844 9864 18896
rect 9916 18884 9922 18896
rect 11609 18887 11667 18893
rect 11609 18884 11621 18887
rect 9916 18856 11621 18884
rect 9916 18844 9922 18856
rect 11609 18853 11621 18856
rect 11655 18853 11667 18887
rect 14737 18887 14795 18893
rect 14737 18884 14749 18887
rect 11609 18847 11667 18853
rect 12268 18856 14749 18884
rect 9950 18776 9956 18828
rect 10008 18776 10014 18828
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10502 18816 10508 18828
rect 10376 18788 10508 18816
rect 10376 18776 10382 18788
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11204 18788 12173 18816
rect 11204 18776 11210 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 9769 18751 9827 18757
rect 8588 18720 9674 18748
rect 4893 18683 4951 18689
rect 4893 18680 4905 18683
rect 4724 18652 4905 18680
rect 4724 18624 4752 18652
rect 4893 18649 4905 18652
rect 4939 18649 4951 18683
rect 6270 18680 6276 18692
rect 6118 18652 6276 18680
rect 4893 18643 4951 18649
rect 6270 18640 6276 18652
rect 6328 18640 6334 18692
rect 6730 18640 6736 18692
rect 6788 18680 6794 18692
rect 7101 18683 7159 18689
rect 7101 18680 7113 18683
rect 6788 18652 7113 18680
rect 6788 18640 6794 18652
rect 7101 18649 7113 18652
rect 7147 18649 7159 18683
rect 8754 18680 8760 18692
rect 7101 18643 7159 18649
rect 8404 18652 8760 18680
rect 2498 18572 2504 18624
rect 2556 18612 2562 18624
rect 3329 18615 3387 18621
rect 3329 18612 3341 18615
rect 2556 18584 3341 18612
rect 2556 18572 2562 18584
rect 3329 18581 3341 18584
rect 3375 18581 3387 18615
rect 3329 18575 3387 18581
rect 3418 18572 3424 18624
rect 3476 18612 3482 18624
rect 3513 18615 3571 18621
rect 3513 18612 3525 18615
rect 3476 18584 3525 18612
rect 3476 18572 3482 18584
rect 3513 18581 3525 18584
rect 3559 18581 3571 18615
rect 3513 18575 3571 18581
rect 4706 18572 4712 18624
rect 4764 18572 4770 18624
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 6365 18615 6423 18621
rect 6365 18612 6377 18615
rect 4856 18584 6377 18612
rect 4856 18572 4862 18584
rect 6365 18581 6377 18584
rect 6411 18612 6423 18615
rect 8404 18612 8432 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 8938 18640 8944 18692
rect 8996 18680 9002 18692
rect 9646 18680 9674 18720
rect 9769 18717 9781 18751
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 9858 18708 9864 18760
rect 9916 18708 9922 18760
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18748 10655 18751
rect 11238 18748 11244 18760
rect 10643 18720 11244 18748
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 12268 18748 12296 18856
rect 14737 18853 14749 18856
rect 14783 18853 14795 18887
rect 14737 18847 14795 18853
rect 13538 18776 13544 18828
rect 13596 18776 13602 18828
rect 11624 18720 12296 18748
rect 10042 18680 10048 18692
rect 8996 18652 9536 18680
rect 9646 18652 10048 18680
rect 8996 18640 9002 18652
rect 6411 18584 8432 18612
rect 6411 18581 6423 18584
rect 6365 18575 6423 18581
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 9033 18615 9091 18621
rect 9033 18612 9045 18615
rect 8628 18584 9045 18612
rect 8628 18572 8634 18584
rect 9033 18581 9045 18584
rect 9079 18612 9091 18615
rect 9122 18612 9128 18624
rect 9079 18584 9128 18612
rect 9079 18581 9091 18584
rect 9033 18575 9091 18581
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 9401 18615 9459 18621
rect 9401 18612 9413 18615
rect 9272 18584 9413 18612
rect 9272 18572 9278 18584
rect 9401 18581 9413 18584
rect 9447 18581 9459 18615
rect 9508 18612 9536 18652
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10965 18683 11023 18689
rect 10965 18680 10977 18683
rect 10284 18652 10977 18680
rect 10284 18640 10290 18652
rect 10965 18649 10977 18652
rect 11011 18680 11023 18683
rect 11624 18680 11652 18720
rect 11011 18652 11652 18680
rect 11011 18649 11023 18652
rect 10965 18643 11023 18649
rect 11698 18640 11704 18692
rect 11756 18680 11762 18692
rect 12069 18683 12127 18689
rect 12069 18680 12081 18683
rect 11756 18652 12081 18680
rect 11756 18640 11762 18652
rect 12069 18649 12081 18652
rect 12115 18649 12127 18683
rect 12069 18643 12127 18649
rect 12802 18640 12808 18692
rect 12860 18640 12866 18692
rect 14553 18683 14611 18689
rect 14553 18649 14565 18683
rect 14599 18680 14611 18683
rect 15120 18680 15148 18924
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22554 18912 22560 18964
rect 22612 18952 22618 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22612 18924 22937 18952
rect 22612 18912 22618 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 30742 18952 30748 18964
rect 22925 18915 22983 18921
rect 23584 18924 30748 18952
rect 17218 18844 17224 18896
rect 17276 18884 17282 18896
rect 18141 18887 18199 18893
rect 17276 18856 17632 18884
rect 17276 18844 17282 18856
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 16206 18816 16212 18828
rect 15243 18788 16212 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 16206 18776 16212 18788
rect 16264 18776 16270 18828
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 16816 18788 17509 18816
rect 16816 18776 16822 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17604 18816 17632 18856
rect 18141 18853 18153 18887
rect 18187 18884 18199 18887
rect 18322 18884 18328 18896
rect 18187 18856 18328 18884
rect 18187 18853 18199 18856
rect 18141 18847 18199 18853
rect 18322 18844 18328 18856
rect 18380 18844 18386 18896
rect 20901 18887 20959 18893
rect 20901 18853 20913 18887
rect 20947 18884 20959 18887
rect 21082 18884 21088 18896
rect 20947 18856 21088 18884
rect 20947 18853 20959 18856
rect 20901 18847 20959 18853
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 17604 18788 18705 18816
rect 17497 18779 17555 18785
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 19760 18788 20361 18816
rect 19760 18776 19766 18788
rect 20349 18785 20361 18788
rect 20395 18816 20407 18819
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 20395 18788 21189 18816
rect 20395 18785 20407 18788
rect 20349 18779 20407 18785
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 21542 18776 21548 18828
rect 21600 18816 21606 18828
rect 23584 18816 23612 18924
rect 30742 18912 30748 18924
rect 30800 18912 30806 18964
rect 48498 18952 48504 18964
rect 35866 18924 48504 18952
rect 29730 18844 29736 18896
rect 29788 18884 29794 18896
rect 30837 18887 30895 18893
rect 30837 18884 30849 18887
rect 29788 18856 30849 18884
rect 29788 18844 29794 18856
rect 30837 18853 30849 18856
rect 30883 18853 30895 18887
rect 30837 18847 30895 18853
rect 30926 18844 30932 18896
rect 30984 18884 30990 18896
rect 35866 18884 35894 18924
rect 48498 18912 48504 18924
rect 48556 18912 48562 18964
rect 30984 18856 35894 18884
rect 30984 18844 30990 18856
rect 21600 18788 23612 18816
rect 21600 18776 21606 18788
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 23716 18788 24593 18816
rect 23716 18776 23722 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25774 18816 25780 18828
rect 25455 18788 25780 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 26418 18776 26424 18828
rect 26476 18816 26482 18828
rect 27157 18819 27215 18825
rect 27157 18816 27169 18819
rect 26476 18788 27169 18816
rect 26476 18776 26482 18788
rect 27157 18785 27169 18788
rect 27203 18785 27215 18819
rect 27157 18779 27215 18785
rect 30190 18776 30196 18828
rect 30248 18776 30254 18828
rect 30285 18819 30343 18825
rect 30285 18785 30297 18819
rect 30331 18785 30343 18819
rect 46842 18816 46848 18828
rect 30285 18779 30343 18785
rect 35866 18788 46848 18816
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 17000 18720 18521 18748
rect 17000 18708 17006 18720
rect 18509 18717 18521 18720
rect 18555 18748 18567 18751
rect 18598 18748 18604 18760
rect 18555 18720 18604 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19659 18720 21220 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 14599 18652 15148 18680
rect 14599 18649 14611 18652
rect 14553 18643 14611 18649
rect 15470 18640 15476 18692
rect 15528 18640 15534 18692
rect 15930 18640 15936 18692
rect 15988 18640 15994 18692
rect 19702 18680 19708 18692
rect 16776 18652 19708 18680
rect 11057 18615 11115 18621
rect 11057 18612 11069 18615
rect 9508 18584 11069 18612
rect 9401 18575 9459 18581
rect 11057 18581 11069 18584
rect 11103 18581 11115 18615
rect 11057 18575 11115 18581
rect 11238 18572 11244 18624
rect 11296 18612 11302 18624
rect 11606 18612 11612 18624
rect 11296 18584 11612 18612
rect 11296 18572 11302 18584
rect 11606 18572 11612 18584
rect 11664 18612 11670 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11664 18584 11989 18612
rect 11664 18572 11670 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 12768 18584 14197 18612
rect 12768 18572 12774 18584
rect 14185 18581 14197 18584
rect 14231 18612 14243 18615
rect 15378 18612 15384 18624
rect 14231 18584 15384 18612
rect 14231 18581 14243 18584
rect 14185 18575 14243 18581
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 15488 18612 15516 18640
rect 16390 18612 16396 18624
rect 15488 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18612 16454 18624
rect 16776 18612 16804 18652
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 21192 18680 21220 18720
rect 23566 18708 23572 18760
rect 23624 18708 23630 18760
rect 24118 18748 24124 18760
rect 23676 18720 24124 18748
rect 21192 18652 21864 18680
rect 22678 18652 22784 18680
rect 16448 18584 16804 18612
rect 16945 18615 17003 18621
rect 16448 18572 16454 18584
rect 16945 18581 16957 18615
rect 16991 18612 17003 18615
rect 17034 18612 17040 18624
rect 16991 18584 17040 18612
rect 16991 18581 17003 18584
rect 16945 18575 17003 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 18049 18615 18107 18621
rect 18049 18612 18061 18615
rect 17184 18584 18061 18612
rect 17184 18572 17190 18584
rect 18049 18581 18061 18584
rect 18095 18612 18107 18615
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18095 18584 18613 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 18601 18581 18613 18584
rect 18647 18612 18659 18615
rect 18690 18612 18696 18624
rect 18647 18584 18696 18612
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 19337 18615 19395 18621
rect 19337 18581 19349 18615
rect 19383 18612 19395 18615
rect 20254 18612 20260 18624
rect 19383 18584 20260 18612
rect 19383 18581 19395 18584
rect 19337 18575 19395 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 21836 18612 21864 18652
rect 22094 18612 22100 18624
rect 21836 18584 22100 18612
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 22756 18612 22784 18652
rect 22922 18640 22928 18692
rect 22980 18680 22986 18692
rect 23676 18680 23704 18720
rect 24118 18708 24124 18720
rect 24176 18708 24182 18760
rect 26786 18708 26792 18760
rect 26844 18708 26850 18760
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 26988 18720 27629 18748
rect 22980 18652 23704 18680
rect 22980 18640 22986 18652
rect 23842 18640 23848 18692
rect 23900 18680 23906 18692
rect 24029 18683 24087 18689
rect 24029 18680 24041 18683
rect 23900 18652 24041 18680
rect 23900 18640 23906 18652
rect 24029 18649 24041 18652
rect 24075 18680 24087 18683
rect 25685 18683 25743 18689
rect 24075 18652 25084 18680
rect 24075 18649 24087 18652
rect 24029 18643 24087 18649
rect 23014 18612 23020 18624
rect 22756 18584 23020 18612
rect 23014 18572 23020 18584
rect 23072 18572 23078 18624
rect 23382 18572 23388 18624
rect 23440 18572 23446 18624
rect 23658 18572 23664 18624
rect 23716 18612 23722 18624
rect 25056 18621 25084 18652
rect 25685 18649 25697 18683
rect 25731 18680 25743 18683
rect 25958 18680 25964 18692
rect 25731 18652 25964 18680
rect 25731 18649 25743 18652
rect 25685 18643 25743 18649
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 24121 18615 24179 18621
rect 24121 18612 24133 18615
rect 23716 18584 24133 18612
rect 23716 18572 23722 18584
rect 24121 18581 24133 18584
rect 24167 18581 24179 18615
rect 24121 18575 24179 18581
rect 25041 18615 25099 18621
rect 25041 18581 25053 18615
rect 25087 18581 25099 18615
rect 25041 18575 25099 18581
rect 25130 18572 25136 18624
rect 25188 18612 25194 18624
rect 26988 18612 27016 18720
rect 27617 18717 27629 18720
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 27893 18751 27951 18757
rect 27893 18748 27905 18751
rect 27764 18720 27905 18748
rect 27764 18708 27770 18720
rect 27893 18717 27905 18720
rect 27939 18717 27951 18751
rect 27893 18711 27951 18717
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 30300 18748 30328 18779
rect 29880 18720 30328 18748
rect 29880 18708 29886 18720
rect 27062 18640 27068 18692
rect 27120 18680 27126 18692
rect 35866 18680 35894 18788
rect 46842 18776 46848 18788
rect 46900 18776 46906 18828
rect 27120 18652 35894 18680
rect 27120 18640 27126 18652
rect 25188 18584 27016 18612
rect 25188 18572 25194 18584
rect 29730 18572 29736 18624
rect 29788 18572 29794 18624
rect 30098 18572 30104 18624
rect 30156 18572 30162 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 5902 18408 5908 18420
rect 2746 18380 5908 18408
rect 2746 18340 2774 18380
rect 5902 18368 5908 18380
rect 5960 18368 5966 18420
rect 6730 18368 6736 18420
rect 6788 18408 6794 18420
rect 6788 18380 7236 18408
rect 6788 18368 6794 18380
rect 1780 18312 2774 18340
rect 7208 18340 7236 18380
rect 7282 18368 7288 18420
rect 7340 18408 7346 18420
rect 8938 18408 8944 18420
rect 7340 18380 8944 18408
rect 7340 18368 7346 18380
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 10134 18408 10140 18420
rect 9784 18380 10140 18408
rect 7926 18340 7932 18352
rect 7208 18312 7932 18340
rect 1780 18281 1808 18312
rect 7926 18300 7932 18312
rect 7984 18300 7990 18352
rect 9122 18300 9128 18352
rect 9180 18340 9186 18352
rect 9784 18340 9812 18380
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10413 18411 10471 18417
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 13354 18408 13360 18420
rect 10459 18380 13360 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 15010 18368 15016 18420
rect 15068 18368 15074 18420
rect 16853 18411 16911 18417
rect 16853 18377 16865 18411
rect 16899 18408 16911 18411
rect 17678 18408 17684 18420
rect 16899 18380 17684 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 21450 18408 21456 18420
rect 18156 18380 21456 18408
rect 9180 18312 9812 18340
rect 9953 18343 10011 18349
rect 9180 18300 9186 18312
rect 9953 18309 9965 18343
rect 9999 18340 10011 18343
rect 12802 18340 12808 18352
rect 9999 18312 12808 18340
rect 9999 18309 10011 18312
rect 9953 18303 10011 18309
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 4246 18272 4252 18284
rect 3651 18244 4252 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 5626 18232 5632 18284
rect 5684 18232 5690 18284
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 6454 18272 6460 18284
rect 5767 18244 6460 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 6454 18232 6460 18244
rect 6512 18232 6518 18284
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 3694 18164 3700 18216
rect 3752 18204 3758 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3752 18176 3893 18204
rect 3752 18164 3758 18176
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 5902 18164 5908 18216
rect 5960 18204 5966 18216
rect 6086 18204 6092 18216
rect 5960 18176 6092 18204
rect 5960 18164 5966 18176
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 4706 18096 4712 18148
rect 4764 18136 4770 18148
rect 6748 18136 6776 18235
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 8444 18244 8493 18272
rect 8444 18232 8450 18244
rect 8481 18241 8493 18244
rect 8527 18272 8539 18275
rect 9968 18272 9996 18303
rect 12802 18300 12808 18312
rect 12860 18340 12866 18352
rect 12860 18312 13216 18340
rect 12860 18300 12866 18312
rect 8527 18244 9996 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 10226 18232 10232 18284
rect 10284 18272 10290 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10284 18244 10793 18272
rect 10284 18232 10290 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 12342 18232 12348 18284
rect 12400 18232 12406 18284
rect 7190 18164 7196 18216
rect 7248 18164 7254 18216
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 8628 18176 9229 18204
rect 8628 18164 8634 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 9548 18176 10885 18204
rect 9548 18164 9554 18176
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 11057 18207 11115 18213
rect 11057 18173 11069 18207
rect 11103 18204 11115 18207
rect 12066 18204 12072 18216
rect 11103 18176 12072 18204
rect 11103 18173 11115 18176
rect 11057 18167 11115 18173
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 12434 18164 12440 18216
rect 12492 18164 12498 18216
rect 12618 18164 12624 18216
rect 12676 18164 12682 18216
rect 13188 18213 13216 18312
rect 14090 18300 14096 18352
rect 14148 18340 14154 18352
rect 14369 18343 14427 18349
rect 14369 18340 14381 18343
rect 14148 18312 14381 18340
rect 14148 18300 14154 18312
rect 14369 18309 14381 18312
rect 14415 18309 14427 18343
rect 14369 18303 14427 18309
rect 14642 18300 14648 18352
rect 14700 18340 14706 18352
rect 18156 18349 18184 18380
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 22557 18411 22615 18417
rect 22557 18377 22569 18411
rect 22603 18408 22615 18411
rect 22646 18408 22652 18420
rect 22603 18380 22652 18408
rect 22603 18377 22615 18380
rect 22557 18371 22615 18377
rect 15381 18343 15439 18349
rect 15381 18340 15393 18343
rect 14700 18312 15393 18340
rect 14700 18300 14706 18312
rect 15381 18309 15393 18312
rect 15427 18309 15439 18343
rect 15381 18303 15439 18309
rect 15473 18343 15531 18349
rect 15473 18309 15485 18343
rect 15519 18340 15531 18343
rect 18141 18343 18199 18349
rect 15519 18312 17540 18340
rect 15519 18309 15531 18312
rect 15473 18303 15531 18309
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 13679 18244 13713 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18204 13231 18207
rect 13648 18204 13676 18235
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16209 18275 16267 18281
rect 16209 18272 16221 18275
rect 15988 18244 16221 18272
rect 15988 18232 15994 18244
rect 16209 18241 16221 18244
rect 16255 18241 16267 18275
rect 16209 18235 16267 18241
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16632 18244 17233 18272
rect 16632 18232 16638 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 15102 18204 15108 18216
rect 13219 18176 15108 18204
rect 13219 18173 13231 18176
rect 13173 18167 13231 18173
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16942 18204 16948 18216
rect 15703 18176 16948 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17313 18207 17371 18213
rect 17313 18173 17325 18207
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 11977 18139 12035 18145
rect 4764 18108 5580 18136
rect 6748 18108 11928 18136
rect 4764 18096 4770 18108
rect 3418 18028 3424 18080
rect 3476 18068 3482 18080
rect 3694 18068 3700 18080
rect 3476 18040 3700 18068
rect 3476 18028 3482 18040
rect 3694 18028 3700 18040
rect 3752 18028 3758 18080
rect 5261 18071 5319 18077
rect 5261 18037 5273 18071
rect 5307 18068 5319 18071
rect 5442 18068 5448 18080
rect 5307 18040 5448 18068
rect 5307 18037 5319 18040
rect 5261 18031 5319 18037
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 5552 18068 5580 18108
rect 9582 18068 9588 18080
rect 5552 18040 9588 18068
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 9674 18028 9680 18080
rect 9732 18028 9738 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9916 18040 10057 18068
rect 9916 18028 9922 18040
rect 10045 18037 10057 18040
rect 10091 18068 10103 18071
rect 10410 18068 10416 18080
rect 10091 18040 10416 18068
rect 10091 18037 10103 18040
rect 10045 18031 10103 18037
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 11698 18028 11704 18080
rect 11756 18028 11762 18080
rect 11900 18068 11928 18108
rect 11977 18105 11989 18139
rect 12023 18136 12035 18139
rect 12158 18136 12164 18148
rect 12023 18108 12164 18136
rect 12023 18105 12035 18108
rect 11977 18099 12035 18105
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 16390 18136 16396 18148
rect 12268 18108 16396 18136
rect 12268 18068 12296 18108
rect 16390 18096 16396 18108
rect 16448 18096 16454 18148
rect 16850 18096 16856 18148
rect 16908 18136 16914 18148
rect 17126 18136 17132 18148
rect 16908 18108 17132 18136
rect 16908 18096 16914 18108
rect 17126 18096 17132 18108
rect 17184 18096 17190 18148
rect 17328 18136 17356 18167
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 17512 18204 17540 18312
rect 18141 18309 18153 18343
rect 18187 18309 18199 18343
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 18141 18303 18199 18309
rect 19306 18312 22017 18340
rect 17586 18232 17592 18284
rect 17644 18272 17650 18284
rect 19306 18272 19334 18312
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22005 18303 22063 18309
rect 17644 18244 19334 18272
rect 19889 18275 19947 18281
rect 17644 18232 17650 18244
rect 19889 18241 19901 18275
rect 19935 18272 19947 18275
rect 20254 18272 20260 18284
rect 19935 18244 20260 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 22572 18272 22600 18371
rect 22646 18368 22652 18380
rect 22704 18408 22710 18420
rect 22833 18411 22891 18417
rect 22833 18408 22845 18411
rect 22704 18380 22845 18408
rect 22704 18368 22710 18380
rect 22833 18377 22845 18380
rect 22879 18408 22891 18411
rect 22922 18408 22928 18420
rect 22879 18380 22928 18408
rect 22879 18377 22891 18380
rect 22833 18371 22891 18377
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 23474 18368 23480 18420
rect 23532 18408 23538 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 23532 18380 24869 18408
rect 23532 18368 23538 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 26786 18368 26792 18420
rect 26844 18368 26850 18420
rect 27157 18411 27215 18417
rect 27157 18377 27169 18411
rect 27203 18408 27215 18411
rect 30098 18408 30104 18420
rect 27203 18380 30104 18408
rect 27203 18377 27215 18380
rect 27157 18371 27215 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 30742 18368 30748 18420
rect 30800 18408 30806 18420
rect 31481 18411 31539 18417
rect 31481 18408 31493 18411
rect 30800 18380 31493 18408
rect 30800 18368 30806 18380
rect 31481 18377 31493 18380
rect 31527 18408 31539 18411
rect 31527 18380 35894 18408
rect 31527 18377 31539 18380
rect 31481 18371 31539 18377
rect 23014 18300 23020 18352
rect 23072 18340 23078 18352
rect 23842 18340 23848 18352
rect 23072 18312 23848 18340
rect 23072 18300 23078 18312
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 26050 18300 26056 18352
rect 26108 18300 26114 18352
rect 28258 18340 28264 18352
rect 28092 18312 28264 18340
rect 21140 18244 22600 18272
rect 21140 18232 21146 18244
rect 25038 18232 25044 18284
rect 25096 18272 25102 18284
rect 28092 18281 28120 18312
rect 28258 18300 28264 18312
rect 28316 18300 28322 18352
rect 28353 18343 28411 18349
rect 28353 18309 28365 18343
rect 28399 18340 28411 18343
rect 28626 18340 28632 18352
rect 28399 18312 28632 18340
rect 28399 18309 28411 18312
rect 28353 18303 28411 18309
rect 28626 18300 28632 18312
rect 28684 18300 28690 18352
rect 29638 18340 29644 18352
rect 29578 18312 29644 18340
rect 29638 18300 29644 18312
rect 29696 18300 29702 18352
rect 30650 18300 30656 18352
rect 30708 18340 30714 18352
rect 31294 18340 31300 18352
rect 30708 18312 31300 18340
rect 30708 18300 30714 18312
rect 31294 18300 31300 18312
rect 31352 18300 31358 18352
rect 25317 18275 25375 18281
rect 25317 18272 25329 18275
rect 25096 18244 25329 18272
rect 25096 18232 25102 18244
rect 25317 18241 25329 18244
rect 25363 18272 25375 18275
rect 26513 18275 26571 18281
rect 26513 18272 26525 18275
rect 25363 18244 26525 18272
rect 25363 18241 25375 18244
rect 25317 18235 25375 18241
rect 26513 18241 26525 18244
rect 26559 18241 26571 18275
rect 26513 18235 26571 18241
rect 28077 18275 28135 18281
rect 28077 18241 28089 18275
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 18138 18204 18144 18216
rect 17512 18176 18144 18204
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 18248 18176 18828 18204
rect 18248 18136 18276 18176
rect 17328 18108 18276 18136
rect 18800 18136 18828 18176
rect 18874 18164 18880 18216
rect 18932 18164 18938 18216
rect 18966 18164 18972 18216
rect 19024 18204 19030 18216
rect 19794 18204 19800 18216
rect 19024 18176 19800 18204
rect 19024 18164 19030 18176
rect 19794 18164 19800 18176
rect 19852 18204 19858 18216
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 19852 18176 19993 18204
rect 19852 18164 19858 18176
rect 19981 18173 19993 18176
rect 20027 18173 20039 18207
rect 19981 18167 20039 18173
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 18800 18108 19656 18136
rect 11900 18040 12296 18068
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13265 18071 13323 18077
rect 13265 18068 13277 18071
rect 12768 18040 13277 18068
rect 12768 18028 12774 18040
rect 13265 18037 13277 18040
rect 13311 18068 13323 18071
rect 13814 18068 13820 18080
rect 13311 18040 13820 18068
rect 13311 18037 13323 18040
rect 13265 18031 13323 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15712 18040 16037 18068
rect 15712 18028 15718 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 16482 18028 16488 18080
rect 16540 18028 16546 18080
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 18233 18071 18291 18077
rect 18233 18068 18245 18071
rect 16816 18040 18245 18068
rect 16816 18028 16822 18040
rect 18233 18037 18245 18040
rect 18279 18037 18291 18071
rect 18233 18031 18291 18037
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 19521 18071 19579 18077
rect 19521 18068 19533 18071
rect 18380 18040 19533 18068
rect 18380 18028 18386 18040
rect 19521 18037 19533 18040
rect 19567 18037 19579 18071
rect 19628 18068 19656 18108
rect 19702 18096 19708 18148
rect 19760 18136 19766 18148
rect 20180 18136 20208 18167
rect 21174 18164 21180 18216
rect 21232 18164 21238 18216
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 23109 18207 23167 18213
rect 23109 18173 23121 18207
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 26234 18204 26240 18216
rect 23431 18176 26240 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 19760 18108 20208 18136
rect 20717 18139 20775 18145
rect 19760 18096 19766 18108
rect 20717 18105 20729 18139
rect 20763 18105 20775 18139
rect 20717 18099 20775 18105
rect 20732 18068 20760 18099
rect 20990 18096 20996 18148
rect 21048 18136 21054 18148
rect 21284 18136 21312 18167
rect 21048 18108 21312 18136
rect 21048 18096 21054 18108
rect 19628 18040 20760 18068
rect 23124 18068 23152 18167
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 27062 18164 27068 18216
rect 27120 18204 27126 18216
rect 30837 18207 30895 18213
rect 27120 18176 30328 18204
rect 27120 18164 27126 18176
rect 30300 18145 30328 18176
rect 30837 18173 30849 18207
rect 30883 18204 30895 18207
rect 34606 18204 34612 18216
rect 30883 18176 34612 18204
rect 30883 18173 30895 18176
rect 30837 18167 30895 18173
rect 30285 18139 30343 18145
rect 30285 18105 30297 18139
rect 30331 18105 30343 18139
rect 30285 18099 30343 18105
rect 30374 18096 30380 18148
rect 30432 18136 30438 18148
rect 30852 18136 30880 18167
rect 34606 18164 34612 18176
rect 34664 18164 34670 18216
rect 30432 18108 30880 18136
rect 35866 18136 35894 18380
rect 41414 18136 41420 18148
rect 35866 18108 41420 18136
rect 30432 18096 30438 18108
rect 41414 18096 41420 18108
rect 41472 18096 41478 18148
rect 24670 18068 24676 18080
rect 23124 18040 24676 18068
rect 19521 18031 19579 18037
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 27338 18028 27344 18080
rect 27396 18068 27402 18080
rect 29822 18068 29828 18080
rect 27396 18040 29828 18068
rect 27396 18028 27402 18040
rect 29822 18028 29828 18040
rect 29880 18028 29886 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 3418 17824 3424 17876
rect 3476 17824 3482 17876
rect 3605 17867 3663 17873
rect 3605 17833 3617 17867
rect 3651 17864 3663 17867
rect 8386 17864 8392 17876
rect 3651 17836 8392 17864
rect 3651 17833 3663 17836
rect 3605 17827 3663 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 10594 17824 10600 17876
rect 10652 17824 10658 17876
rect 13446 17864 13452 17876
rect 11716 17836 13452 17864
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 4433 17799 4491 17805
rect 4433 17796 4445 17799
rect 1912 17768 4445 17796
rect 1912 17756 1918 17768
rect 4433 17765 4445 17768
rect 4479 17765 4491 17799
rect 4433 17759 4491 17765
rect 6178 17756 6184 17808
rect 6236 17796 6242 17808
rect 6641 17799 6699 17805
rect 6641 17796 6653 17799
rect 6236 17768 6653 17796
rect 6236 17756 6242 17768
rect 6641 17765 6653 17768
rect 6687 17765 6699 17799
rect 6641 17759 6699 17765
rect 7834 17756 7840 17808
rect 7892 17756 7898 17808
rect 8018 17756 8024 17808
rect 8076 17796 8082 17808
rect 8846 17796 8852 17808
rect 8076 17768 8852 17796
rect 8076 17756 8082 17768
rect 8846 17756 8852 17768
rect 8904 17756 8910 17808
rect 10318 17756 10324 17808
rect 10376 17796 10382 17808
rect 11514 17796 11520 17808
rect 10376 17768 11520 17796
rect 10376 17756 10382 17768
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 1780 17700 7389 17728
rect 1780 17669 1808 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 7926 17688 7932 17740
rect 7984 17728 7990 17740
rect 8481 17731 8539 17737
rect 8481 17728 8493 17731
rect 7984 17700 8493 17728
rect 7984 17688 7990 17700
rect 8481 17697 8493 17700
rect 8527 17728 8539 17731
rect 8527 17700 9260 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17629 1823 17663
rect 1765 17623 1823 17629
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4614 17660 4620 17672
rect 4212 17632 4620 17660
rect 4212 17620 4218 17632
rect 4614 17620 4620 17632
rect 4672 17660 4678 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4672 17632 4905 17660
rect 4672 17620 4678 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 6270 17620 6276 17672
rect 6328 17620 6334 17672
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 7650 17620 7656 17672
rect 7708 17660 7714 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7708 17632 8217 17660
rect 7708 17620 7714 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 8386 17620 8392 17672
rect 8444 17660 8450 17672
rect 8570 17660 8576 17672
rect 8444 17632 8576 17660
rect 8444 17620 8450 17632
rect 8570 17620 8576 17632
rect 8628 17660 8634 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 8628 17632 9137 17660
rect 8628 17620 8634 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9232 17660 9260 17700
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9456 17700 9873 17728
rect 9456 17688 9462 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10100 17700 11161 17728
rect 10100 17688 10106 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11480 17700 11621 17728
rect 11480 17688 11486 17700
rect 11609 17697 11621 17700
rect 11655 17697 11667 17731
rect 11609 17691 11667 17697
rect 10870 17660 10876 17672
rect 9232 17632 10876 17660
rect 9125 17623 9183 17629
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11716 17660 11744 17836
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 13722 17824 13728 17876
rect 13780 17824 13786 17876
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 16206 17864 16212 17876
rect 15896 17836 16212 17864
rect 15896 17824 15902 17836
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 16390 17824 16396 17876
rect 16448 17864 16454 17876
rect 20717 17867 20775 17873
rect 20717 17864 20729 17867
rect 16448 17836 20729 17864
rect 16448 17824 16454 17836
rect 20717 17833 20729 17836
rect 20763 17833 20775 17867
rect 30929 17867 30987 17873
rect 30929 17864 30941 17867
rect 20717 17827 20775 17833
rect 21192 17836 30941 17864
rect 13262 17756 13268 17808
rect 13320 17796 13326 17808
rect 14918 17796 14924 17808
rect 13320 17768 14924 17796
rect 13320 17756 13326 17768
rect 14918 17756 14924 17768
rect 14976 17756 14982 17808
rect 18325 17799 18383 17805
rect 18325 17796 18337 17799
rect 17696 17768 18337 17796
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12618 17728 12624 17740
rect 12299 17700 12624 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 14553 17731 14611 17737
rect 14553 17728 14565 17731
rect 12860 17700 14565 17728
rect 12860 17688 12866 17700
rect 14553 17697 14565 17700
rect 14599 17697 14611 17731
rect 14553 17691 14611 17697
rect 16298 17688 16304 17740
rect 16356 17688 16362 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16942 17728 16948 17740
rect 16623 17700 16948 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 11011 17632 11744 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 15010 17660 15016 17672
rect 14415 17632 15016 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 934 17552 940 17604
rect 992 17592 998 17604
rect 2501 17595 2559 17601
rect 2501 17592 2513 17595
rect 992 17564 2513 17592
rect 992 17552 998 17564
rect 2501 17561 2513 17564
rect 2547 17561 2559 17595
rect 2501 17555 2559 17561
rect 4246 17552 4252 17604
rect 4304 17552 4310 17604
rect 5169 17595 5227 17601
rect 5169 17561 5181 17595
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 2130 17484 2136 17536
rect 2188 17524 2194 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 2188 17496 3801 17524
rect 2188 17484 2194 17496
rect 3789 17493 3801 17496
rect 3835 17524 3847 17527
rect 4798 17524 4804 17536
rect 3835 17496 4804 17524
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 5184 17524 5212 17555
rect 7466 17552 7472 17604
rect 7524 17592 7530 17604
rect 8297 17595 8355 17601
rect 7524 17564 8156 17592
rect 7524 17552 7530 17564
rect 8018 17524 8024 17536
rect 5184 17496 8024 17524
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 8128 17524 8156 17564
rect 8297 17561 8309 17595
rect 8343 17592 8355 17595
rect 9214 17592 9220 17604
rect 8343 17564 9220 17592
rect 8343 17561 8355 17564
rect 8297 17555 8355 17561
rect 9214 17552 9220 17564
rect 9272 17552 9278 17604
rect 9398 17552 9404 17604
rect 9456 17592 9462 17604
rect 11057 17595 11115 17601
rect 11057 17592 11069 17595
rect 9456 17564 11069 17592
rect 9456 17552 9462 17564
rect 11057 17561 11069 17564
rect 11103 17561 11115 17595
rect 11057 17555 11115 17561
rect 12250 17552 12256 17604
rect 12308 17592 12314 17604
rect 12710 17592 12716 17604
rect 12308 17564 12716 17592
rect 12308 17552 12314 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 13814 17552 13820 17604
rect 13872 17592 13878 17604
rect 14918 17592 14924 17604
rect 13872 17564 14924 17592
rect 13872 17552 13878 17564
rect 14918 17552 14924 17564
rect 14976 17552 14982 17604
rect 15286 17552 15292 17604
rect 15344 17592 15350 17604
rect 15344 17564 15976 17592
rect 15344 17552 15350 17564
rect 15948 17536 15976 17564
rect 12066 17524 12072 17536
rect 8128 17496 12072 17524
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 14829 17527 14887 17533
rect 14829 17493 14841 17527
rect 14875 17524 14887 17527
rect 15010 17524 15016 17536
rect 14875 17496 15016 17524
rect 14875 17493 14887 17496
rect 14829 17487 14887 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 15102 17484 15108 17536
rect 15160 17484 15166 17536
rect 15194 17484 15200 17536
rect 15252 17524 15258 17536
rect 15381 17527 15439 17533
rect 15381 17524 15393 17527
rect 15252 17496 15393 17524
rect 15252 17484 15258 17496
rect 15381 17493 15393 17496
rect 15427 17493 15439 17527
rect 15381 17487 15439 17493
rect 15930 17484 15936 17536
rect 15988 17524 15994 17536
rect 16025 17527 16083 17533
rect 16025 17524 16037 17527
rect 15988 17496 16037 17524
rect 15988 17484 15994 17496
rect 16025 17493 16037 17496
rect 16071 17524 16083 17527
rect 16298 17524 16304 17536
rect 16071 17496 16304 17524
rect 16071 17493 16083 17496
rect 16025 17487 16083 17493
rect 16298 17484 16304 17496
rect 16356 17524 16362 17536
rect 17696 17524 17724 17768
rect 18325 17765 18337 17768
rect 18371 17765 18383 17799
rect 21082 17796 21088 17808
rect 18325 17759 18383 17765
rect 19306 17768 21088 17796
rect 17770 17688 17776 17740
rect 17828 17728 17834 17740
rect 19306 17728 19334 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 17828 17700 19334 17728
rect 17828 17688 17834 17700
rect 19426 17688 19432 17740
rect 19484 17688 19490 17740
rect 20990 17728 20996 17740
rect 19536 17700 20996 17728
rect 19536 17660 19564 17700
rect 20990 17688 20996 17700
rect 21048 17688 21054 17740
rect 21192 17737 21220 17836
rect 30929 17833 30941 17836
rect 30975 17833 30987 17867
rect 30929 17827 30987 17833
rect 22005 17799 22063 17805
rect 22005 17765 22017 17799
rect 22051 17796 22063 17799
rect 22278 17796 22284 17808
rect 22051 17768 22284 17796
rect 22051 17765 22063 17768
rect 22005 17759 22063 17765
rect 22278 17756 22284 17768
rect 22336 17756 22342 17808
rect 26234 17756 26240 17808
rect 26292 17796 26298 17808
rect 26605 17799 26663 17805
rect 26605 17796 26617 17799
rect 26292 17768 26617 17796
rect 26292 17756 26298 17768
rect 26605 17765 26617 17768
rect 26651 17765 26663 17799
rect 26605 17759 26663 17765
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 29733 17799 29791 17805
rect 29733 17796 29745 17799
rect 28500 17768 29745 17796
rect 28500 17756 28506 17768
rect 29733 17765 29745 17768
rect 29779 17765 29791 17799
rect 29733 17759 29791 17765
rect 21177 17731 21235 17737
rect 21177 17697 21189 17731
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 21269 17731 21327 17737
rect 21269 17697 21281 17731
rect 21315 17728 21327 17731
rect 24578 17728 24584 17740
rect 21315 17700 24584 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 18340 17632 19564 17660
rect 18340 17536 18368 17632
rect 19702 17620 19708 17672
rect 19760 17620 19766 17672
rect 20438 17620 20444 17672
rect 20496 17660 20502 17672
rect 21284 17660 21312 17691
rect 24578 17688 24584 17700
rect 24636 17688 24642 17740
rect 24670 17688 24676 17740
rect 24728 17728 24734 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24728 17700 24869 17728
rect 24728 17688 24734 17700
rect 24857 17697 24869 17700
rect 24903 17728 24915 17731
rect 25774 17728 25780 17740
rect 24903 17700 25780 17728
rect 24903 17697 24915 17700
rect 24857 17691 24915 17697
rect 25774 17688 25780 17700
rect 25832 17728 25838 17740
rect 27065 17731 27123 17737
rect 27065 17728 27077 17731
rect 25832 17700 27077 17728
rect 25832 17688 25838 17700
rect 27065 17697 27077 17700
rect 27111 17728 27123 17731
rect 28350 17728 28356 17740
rect 27111 17700 28356 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 28350 17688 28356 17700
rect 28408 17688 28414 17740
rect 29181 17731 29239 17737
rect 29181 17728 29193 17731
rect 28460 17700 29193 17728
rect 20496 17632 21312 17660
rect 20496 17620 20502 17632
rect 22002 17620 22008 17672
rect 22060 17660 22066 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22060 17632 22293 17660
rect 22060 17620 22066 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 28460 17646 28488 17700
rect 29181 17697 29193 17700
rect 29227 17728 29239 17731
rect 29638 17728 29644 17740
rect 29227 17700 29644 17728
rect 29227 17697 29239 17700
rect 29181 17691 29239 17697
rect 29638 17688 29644 17700
rect 29696 17688 29702 17740
rect 30282 17688 30288 17740
rect 30340 17688 30346 17740
rect 31481 17731 31539 17737
rect 31481 17728 31493 17731
rect 30392 17700 31493 17728
rect 22281 17623 22339 17629
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 30392 17660 30420 17700
rect 31481 17697 31493 17700
rect 31527 17697 31539 17731
rect 31481 17691 31539 17697
rect 28868 17632 30420 17660
rect 28868 17620 28874 17632
rect 31018 17620 31024 17672
rect 31076 17660 31082 17672
rect 31297 17663 31355 17669
rect 31297 17660 31309 17663
rect 31076 17632 31309 17660
rect 31076 17620 31082 17632
rect 31297 17629 31309 17632
rect 31343 17629 31355 17663
rect 31297 17623 31355 17629
rect 31389 17663 31447 17669
rect 31389 17629 31401 17663
rect 31435 17660 31447 17663
rect 34514 17660 34520 17672
rect 31435 17632 34520 17660
rect 31435 17629 31447 17632
rect 31389 17623 31447 17629
rect 34514 17620 34520 17632
rect 34572 17620 34578 17672
rect 18874 17552 18880 17604
rect 18932 17592 18938 17604
rect 21085 17595 21143 17601
rect 21085 17592 21097 17595
rect 18932 17564 21097 17592
rect 18932 17552 18938 17564
rect 21085 17561 21097 17564
rect 21131 17561 21143 17595
rect 22557 17595 22615 17601
rect 22557 17592 22569 17595
rect 21085 17555 21143 17561
rect 21192 17564 22569 17592
rect 16356 17496 17724 17524
rect 18049 17527 18107 17533
rect 16356 17484 16362 17496
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18322 17524 18328 17536
rect 18095 17496 18328 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 18690 17484 18696 17536
rect 18748 17484 18754 17536
rect 19886 17484 19892 17536
rect 19944 17524 19950 17536
rect 21192 17524 21220 17564
rect 22557 17561 22569 17564
rect 22603 17561 22615 17595
rect 23842 17592 23848 17604
rect 23782 17564 23848 17592
rect 22557 17555 22615 17561
rect 23842 17552 23848 17564
rect 23900 17552 23906 17604
rect 25130 17592 25136 17604
rect 24044 17564 25136 17592
rect 19944 17496 21220 17524
rect 21821 17527 21879 17533
rect 19944 17484 19950 17496
rect 21821 17493 21833 17527
rect 21867 17524 21879 17527
rect 21910 17524 21916 17536
rect 21867 17496 21916 17524
rect 21867 17493 21879 17496
rect 21821 17487 21879 17493
rect 21910 17484 21916 17496
rect 21968 17524 21974 17536
rect 23474 17524 23480 17536
rect 21968 17496 23480 17524
rect 21968 17484 21974 17496
rect 23474 17484 23480 17496
rect 23532 17524 23538 17536
rect 23860 17524 23888 17552
rect 24044 17533 24072 17564
rect 25130 17552 25136 17564
rect 25188 17552 25194 17604
rect 26786 17592 26792 17604
rect 26358 17564 26792 17592
rect 26786 17552 26792 17564
rect 26844 17552 26850 17604
rect 27338 17552 27344 17604
rect 27396 17552 27402 17604
rect 30101 17595 30159 17601
rect 30101 17592 30113 17595
rect 28644 17564 30113 17592
rect 23532 17496 23888 17524
rect 24029 17527 24087 17533
rect 23532 17484 23538 17496
rect 24029 17493 24041 17527
rect 24075 17493 24087 17527
rect 24029 17487 24087 17493
rect 24394 17484 24400 17536
rect 24452 17524 24458 17536
rect 28644 17524 28672 17564
rect 30101 17561 30113 17564
rect 30147 17592 30159 17595
rect 30926 17592 30932 17604
rect 30147 17564 30932 17592
rect 30147 17561 30159 17564
rect 30101 17555 30159 17561
rect 30926 17552 30932 17564
rect 30984 17552 30990 17604
rect 24452 17496 28672 17524
rect 24452 17484 24458 17496
rect 28810 17484 28816 17536
rect 28868 17484 28874 17536
rect 30190 17484 30196 17536
rect 30248 17484 30254 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 5261 17323 5319 17329
rect 3528 17292 5212 17320
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 3528 17184 3556 17292
rect 4617 17255 4675 17261
rect 4617 17221 4629 17255
rect 4663 17252 4675 17255
rect 5074 17252 5080 17264
rect 4663 17224 5080 17252
rect 4663 17221 4675 17224
rect 4617 17215 4675 17221
rect 5074 17212 5080 17224
rect 5132 17212 5138 17264
rect 5184 17252 5212 17292
rect 5261 17289 5273 17323
rect 5307 17320 5319 17323
rect 7285 17323 7343 17329
rect 7285 17320 7297 17323
rect 5307 17292 7297 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 7285 17289 7297 17292
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7800 17292 8033 17320
rect 7800 17280 7806 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 9122 17320 9128 17332
rect 8021 17283 8079 17289
rect 8128 17292 9128 17320
rect 8128 17252 8156 17292
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 9548 17292 9965 17320
rect 9548 17280 9554 17292
rect 9953 17289 9965 17292
rect 9999 17320 10011 17323
rect 9999 17292 12434 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 5184 17224 8156 17252
rect 8386 17212 8392 17264
rect 8444 17212 8450 17264
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 9646 17224 10977 17252
rect 1811 17156 3556 17184
rect 3605 17187 3663 17193
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 3786 17184 3792 17196
rect 3651 17156 3792 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5184 17156 5641 17184
rect 1118 17076 1124 17128
rect 1176 17116 1182 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1176 17088 2053 17116
rect 1176 17076 1182 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 4430 17076 4436 17128
rect 4488 17116 4494 17128
rect 5184 17125 5212 17156
rect 5629 17153 5641 17156
rect 5675 17184 5687 17187
rect 6086 17184 6092 17196
rect 5675 17156 6092 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 8570 17144 8576 17196
rect 8628 17144 8634 17196
rect 9490 17144 9496 17196
rect 9548 17184 9554 17196
rect 9646 17184 9674 17224
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11480 17224 11805 17252
rect 11480 17212 11486 17224
rect 11793 17221 11805 17224
rect 11839 17221 11851 17255
rect 11793 17215 11851 17221
rect 9548 17156 9674 17184
rect 9548 17144 9554 17156
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17153 10839 17187
rect 12406 17184 12434 17292
rect 12526 17280 12532 17332
rect 12584 17280 12590 17332
rect 13725 17323 13783 17329
rect 13725 17289 13737 17323
rect 13771 17320 13783 17323
rect 14642 17320 14648 17332
rect 13771 17292 14648 17320
rect 13771 17289 13783 17292
rect 13725 17283 13783 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 16853 17323 16911 17329
rect 16853 17320 16865 17323
rect 14884 17292 16865 17320
rect 14884 17280 14890 17292
rect 16853 17289 16865 17292
rect 16899 17289 16911 17323
rect 16853 17283 16911 17289
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17770 17320 17776 17332
rect 17092 17292 17776 17320
rect 17092 17280 17098 17292
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 22005 17323 22063 17329
rect 22005 17320 22017 17323
rect 17920 17292 22017 17320
rect 17920 17280 17926 17292
rect 22005 17289 22017 17292
rect 22051 17289 22063 17323
rect 23934 17320 23940 17332
rect 22005 17283 22063 17289
rect 22204 17292 23940 17320
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 13814 17252 13820 17264
rect 13035 17224 13820 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 14274 17212 14280 17264
rect 14332 17252 14338 17264
rect 18322 17252 18328 17264
rect 14332 17224 18328 17252
rect 14332 17212 14338 17224
rect 18322 17212 18328 17224
rect 18380 17252 18386 17264
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 18380 17224 18429 17252
rect 18380 17212 18386 17224
rect 18417 17221 18429 17224
rect 18463 17221 18475 17255
rect 18417 17215 18475 17221
rect 20070 17212 20076 17264
rect 20128 17252 20134 17264
rect 20165 17255 20223 17261
rect 20165 17252 20177 17255
rect 20128 17224 20177 17252
rect 20128 17212 20134 17224
rect 20165 17221 20177 17224
rect 20211 17221 20223 17255
rect 20165 17215 20223 17221
rect 12526 17184 12532 17196
rect 12406 17156 12532 17184
rect 10781 17147 10839 17153
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4488 17088 4997 17116
rect 4488 17076 4494 17088
rect 4985 17085 4997 17088
rect 5031 17116 5043 17119
rect 5169 17119 5227 17125
rect 5169 17116 5181 17119
rect 5031 17088 5181 17116
rect 5031 17085 5043 17088
rect 4985 17079 5043 17085
rect 5169 17085 5181 17088
rect 5215 17085 5227 17119
rect 5169 17079 5227 17085
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 2498 17008 2504 17060
rect 2556 17048 2562 17060
rect 2556 17020 5580 17048
rect 2556 17008 2562 17020
rect 5166 16940 5172 16992
rect 5224 16980 5230 16992
rect 5350 16980 5356 16992
rect 5224 16952 5356 16980
rect 5224 16940 5230 16952
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5552 16980 5580 17020
rect 5626 17008 5632 17060
rect 5684 17048 5690 17060
rect 5736 17048 5764 17079
rect 5810 17076 5816 17128
rect 5868 17076 5874 17128
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7834 17116 7840 17128
rect 7515 17088 7840 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 8202 17076 8208 17128
rect 8260 17116 8266 17128
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 8260 17088 8493 17116
rect 8260 17076 8266 17088
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 8588 17060 8616 17144
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 8754 17116 8760 17128
rect 8711 17088 8760 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 9398 17076 9404 17128
rect 9456 17116 9462 17128
rect 9766 17116 9772 17128
rect 9456 17088 9772 17116
rect 9456 17076 9462 17088
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 10134 17076 10140 17128
rect 10192 17116 10198 17128
rect 10686 17116 10692 17128
rect 10192 17088 10692 17116
rect 10192 17076 10198 17088
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 10796 17116 10824 17147
rect 12526 17144 12532 17156
rect 12584 17184 12590 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12584 17156 12909 17184
rect 12584 17144 12590 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 13906 17184 13912 17196
rect 12897 17147 12955 17153
rect 13096 17156 13912 17184
rect 13096 17116 13124 17156
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 14090 17144 14096 17196
rect 14148 17144 14154 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14200 17156 14749 17184
rect 14200 17128 14228 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 14918 17144 14924 17196
rect 14976 17144 14982 17196
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17184 15255 17187
rect 15286 17184 15292 17196
rect 15243 17156 15292 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17184 15715 17187
rect 15838 17184 15844 17196
rect 15703 17156 15844 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 17126 17184 17132 17196
rect 16347 17156 17132 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 17218 17144 17224 17196
rect 17276 17144 17282 17196
rect 20180 17184 20208 17215
rect 20898 17212 20904 17264
rect 20956 17252 20962 17264
rect 22204 17252 22232 17292
rect 23934 17280 23940 17292
rect 23992 17280 23998 17332
rect 24210 17280 24216 17332
rect 24268 17320 24274 17332
rect 24305 17323 24363 17329
rect 24305 17320 24317 17323
rect 24268 17292 24317 17320
rect 24268 17280 24274 17292
rect 24305 17289 24317 17292
rect 24351 17289 24363 17323
rect 28810 17320 28816 17332
rect 24305 17283 24363 17289
rect 24964 17292 28816 17320
rect 20956 17224 22232 17252
rect 20956 17212 20962 17224
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 22465 17255 22523 17261
rect 22465 17252 22477 17255
rect 22336 17224 22477 17252
rect 22336 17212 22342 17224
rect 22465 17221 22477 17224
rect 22511 17252 22523 17255
rect 23106 17252 23112 17264
rect 22511 17224 23112 17252
rect 22511 17221 22523 17224
rect 22465 17215 22523 17221
rect 23106 17212 23112 17224
rect 23164 17212 23170 17264
rect 24964 17261 24992 17292
rect 28810 17280 28816 17292
rect 28868 17280 28874 17332
rect 29638 17280 29644 17332
rect 29696 17320 29702 17332
rect 29825 17323 29883 17329
rect 29825 17320 29837 17323
rect 29696 17292 29837 17320
rect 29696 17280 29702 17292
rect 29825 17289 29837 17292
rect 29871 17289 29883 17323
rect 29825 17283 29883 17289
rect 30190 17280 30196 17332
rect 30248 17320 30254 17332
rect 30561 17323 30619 17329
rect 30561 17320 30573 17323
rect 30248 17292 30573 17320
rect 30248 17280 30254 17292
rect 30561 17289 30573 17292
rect 30607 17289 30619 17323
rect 30561 17283 30619 17289
rect 30926 17280 30932 17332
rect 30984 17320 30990 17332
rect 30984 17292 31754 17320
rect 30984 17280 30990 17292
rect 24949 17255 25007 17261
rect 24949 17221 24961 17255
rect 24995 17221 25007 17255
rect 26234 17252 26240 17264
rect 26174 17224 26240 17252
rect 24949 17215 25007 17221
rect 26234 17212 26240 17224
rect 26292 17252 26298 17264
rect 26786 17252 26792 17264
rect 26292 17224 26792 17252
rect 26292 17212 26298 17224
rect 26786 17212 26792 17224
rect 26844 17212 26850 17264
rect 28350 17252 28356 17264
rect 27816 17224 28356 17252
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 10796 17088 13124 17116
rect 13173 17119 13231 17125
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13722 17116 13728 17128
rect 13219 17088 13728 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 14182 17076 14188 17128
rect 14240 17076 14246 17128
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 15470 17116 15476 17128
rect 14415 17088 15476 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 15930 17076 15936 17128
rect 15988 17116 15994 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 15988 17088 17325 17116
rect 15988 17076 15994 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 5684 17020 5764 17048
rect 6012 17020 6592 17048
rect 5684 17008 5690 17020
rect 6012 16980 6040 17020
rect 5552 16952 6040 16980
rect 6454 16940 6460 16992
rect 6512 16940 6518 16992
rect 6564 16980 6592 17020
rect 6638 17008 6644 17060
rect 6696 17048 6702 17060
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 6696 17020 6837 17048
rect 6696 17008 6702 17020
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 8570 17008 8576 17060
rect 8628 17008 8634 17060
rect 11977 17051 12035 17057
rect 11977 17048 11989 17051
rect 9692 17020 11989 17048
rect 9125 16983 9183 16989
rect 9125 16980 9137 16983
rect 6564 16952 9137 16980
rect 9125 16949 9137 16952
rect 9171 16980 9183 16983
rect 9398 16980 9404 16992
rect 9171 16952 9404 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 9490 16940 9496 16992
rect 9548 16940 9554 16992
rect 9582 16940 9588 16992
rect 9640 16980 9646 16992
rect 9692 16980 9720 17020
rect 11977 17017 11989 17020
rect 12023 17017 12035 17051
rect 11977 17011 12035 17017
rect 12066 17008 12072 17060
rect 12124 17048 12130 17060
rect 16117 17051 16175 17057
rect 16117 17048 16129 17051
rect 12124 17020 16129 17048
rect 12124 17008 12130 17020
rect 16117 17017 16129 17020
rect 16163 17017 16175 17051
rect 16117 17011 16175 17017
rect 17420 16992 17448 17079
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17828 17088 18153 17116
rect 17828 17076 17834 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18966 17116 18972 17128
rect 18141 17079 18199 17085
rect 18248 17088 18972 17116
rect 17954 17008 17960 17060
rect 18012 17048 18018 17060
rect 18248 17048 18276 17088
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 18012 17020 18276 17048
rect 19536 17048 19564 17170
rect 20180 17156 21097 17184
rect 21085 17153 21097 17156
rect 21131 17184 21143 17187
rect 22296 17184 22324 17212
rect 21131 17156 22324 17184
rect 22373 17187 22431 17193
rect 21131 17153 21143 17156
rect 21085 17147 21143 17153
rect 22373 17153 22385 17187
rect 22419 17184 22431 17187
rect 22646 17184 22652 17196
rect 22419 17156 22652 17184
rect 22419 17153 22431 17156
rect 22373 17147 22431 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17184 23719 17187
rect 24394 17184 24400 17196
rect 23707 17156 24400 17184
rect 23707 17153 23719 17156
rect 23661 17147 23719 17153
rect 20346 17076 20352 17128
rect 20404 17116 20410 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 20404 17088 21189 17116
rect 20404 17076 20410 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17085 21419 17119
rect 21361 17079 21419 17085
rect 21082 17048 21088 17060
rect 19536 17020 21088 17048
rect 18012 17008 18018 17020
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 9640 16952 9720 16980
rect 11333 16983 11391 16989
rect 9640 16940 9646 16952
rect 11333 16949 11345 16983
rect 11379 16980 11391 16983
rect 11606 16980 11612 16992
rect 11379 16952 11612 16980
rect 11379 16949 11391 16952
rect 11333 16943 11391 16949
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 12768 16952 15485 16980
rect 12768 16940 12774 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 15746 16940 15752 16992
rect 15804 16980 15810 16992
rect 16482 16980 16488 16992
rect 15804 16952 16488 16980
rect 15804 16940 15810 16952
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 17402 16940 17408 16992
rect 17460 16940 17466 16992
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 19886 16980 19892 16992
rect 17552 16952 19892 16980
rect 17552 16940 17558 16952
rect 19886 16940 19892 16952
rect 19944 16940 19950 16992
rect 20346 16940 20352 16992
rect 20404 16940 20410 16992
rect 20714 16940 20720 16992
rect 20772 16940 20778 16992
rect 21192 16980 21220 17079
rect 21376 17048 21404 17079
rect 21910 17076 21916 17128
rect 21968 17116 21974 17128
rect 21968 17088 22508 17116
rect 21968 17076 21974 17088
rect 21818 17048 21824 17060
rect 21376 17020 21824 17048
rect 21818 17008 21824 17020
rect 21876 17008 21882 17060
rect 22480 17048 22508 17088
rect 22554 17076 22560 17128
rect 22612 17076 22618 17128
rect 23676 17048 23704 17147
rect 24394 17144 24400 17156
rect 24452 17144 24458 17196
rect 24670 17144 24676 17196
rect 24728 17144 24734 17196
rect 27816 17193 27844 17224
rect 28350 17212 28356 17224
rect 28408 17212 28414 17264
rect 29656 17252 29684 17280
rect 29302 17224 29684 17252
rect 30837 17255 30895 17261
rect 30837 17221 30849 17255
rect 30883 17252 30895 17255
rect 31018 17252 31024 17264
rect 30883 17224 31024 17252
rect 30883 17221 30895 17224
rect 30837 17215 30895 17221
rect 31018 17212 31024 17224
rect 31076 17212 31082 17264
rect 27801 17187 27859 17193
rect 27801 17153 27813 17187
rect 27847 17153 27859 17187
rect 27801 17147 27859 17153
rect 23750 17076 23756 17128
rect 23808 17076 23814 17128
rect 23842 17076 23848 17128
rect 23900 17076 23906 17128
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 26421 17119 26479 17125
rect 26421 17116 26433 17119
rect 24636 17088 26433 17116
rect 24636 17076 24642 17088
rect 26421 17085 26433 17088
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27614 17116 27620 17128
rect 27203 17088 27620 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17116 28135 17119
rect 30282 17116 30288 17128
rect 28123 17088 30288 17116
rect 28123 17085 28135 17088
rect 28077 17079 28135 17085
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 22480 17020 23704 17048
rect 30190 17008 30196 17060
rect 30248 17048 30254 17060
rect 31726 17048 31754 17292
rect 34514 17212 34520 17264
rect 34572 17252 34578 17264
rect 48314 17252 48320 17264
rect 34572 17224 48320 17252
rect 34572 17212 34578 17224
rect 48314 17212 48320 17224
rect 48372 17212 48378 17264
rect 47210 17048 47216 17060
rect 30248 17020 30880 17048
rect 31726 17020 47216 17048
rect 30248 17008 30254 17020
rect 21542 16980 21548 16992
rect 21192 16952 21548 16980
rect 21542 16940 21548 16952
rect 21600 16980 21606 16992
rect 21726 16980 21732 16992
rect 21600 16952 21732 16980
rect 21600 16940 21606 16952
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 23290 16940 23296 16992
rect 23348 16940 23354 16992
rect 24578 16940 24584 16992
rect 24636 16980 24642 16992
rect 25038 16980 25044 16992
rect 24636 16952 25044 16980
rect 24636 16940 24642 16952
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 25130 16940 25136 16992
rect 25188 16980 25194 16992
rect 25958 16980 25964 16992
rect 25188 16952 25964 16980
rect 25188 16940 25194 16952
rect 25958 16940 25964 16952
rect 26016 16940 26022 16992
rect 27246 16940 27252 16992
rect 27304 16980 27310 16992
rect 29549 16983 29607 16989
rect 29549 16980 29561 16983
rect 27304 16952 29561 16980
rect 27304 16940 27310 16952
rect 29549 16949 29561 16952
rect 29595 16949 29607 16983
rect 30852 16980 30880 17020
rect 47210 17008 47216 17020
rect 47268 17008 47274 17060
rect 47026 16980 47032 16992
rect 30852 16952 47032 16980
rect 29549 16943 29607 16949
rect 47026 16940 47032 16952
rect 47084 16940 47090 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 3605 16779 3663 16785
rect 3605 16745 3617 16779
rect 3651 16776 3663 16779
rect 5074 16776 5080 16788
rect 3651 16748 5080 16776
rect 3651 16745 3663 16748
rect 3605 16739 3663 16745
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 5718 16736 5724 16788
rect 5776 16776 5782 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5776 16748 6009 16776
rect 5776 16736 5782 16748
rect 5997 16745 6009 16748
rect 6043 16745 6055 16779
rect 5997 16739 6055 16745
rect 7837 16779 7895 16785
rect 7837 16745 7849 16779
rect 7883 16776 7895 16779
rect 7883 16748 9168 16776
rect 7883 16745 7895 16748
rect 7837 16739 7895 16745
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 6178 16708 6184 16720
rect 2648 16680 6184 16708
rect 2648 16668 2654 16680
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 9140 16708 9168 16748
rect 9214 16736 9220 16788
rect 9272 16776 9278 16788
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 9272 16748 9781 16776
rect 9272 16736 9278 16748
rect 9769 16745 9781 16748
rect 9815 16776 9827 16779
rect 10410 16776 10416 16788
rect 9815 16748 10416 16776
rect 9815 16745 9827 16748
rect 9769 16739 9827 16745
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 11882 16776 11888 16788
rect 11572 16748 11888 16776
rect 11572 16736 11578 16748
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12526 16736 12532 16788
rect 12584 16736 12590 16788
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 13722 16776 13728 16788
rect 12676 16748 13728 16776
rect 12676 16736 12682 16748
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 18874 16776 18880 16788
rect 13832 16748 18880 16776
rect 9306 16708 9312 16720
rect 8128 16680 8524 16708
rect 9140 16680 9312 16708
rect 3418 16600 3424 16652
rect 3476 16600 3482 16652
rect 3988 16612 4200 16640
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 3988 16572 4016 16612
rect 1811 16544 4016 16572
rect 4065 16575 4123 16581
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4172 16572 4200 16612
rect 6822 16600 6828 16652
rect 6880 16640 6886 16652
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 6880 16612 7113 16640
rect 6880 16600 6886 16612
rect 7101 16609 7113 16612
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 8128 16640 8156 16680
rect 7331 16612 8156 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 8496 16649 8524 16680
rect 9306 16668 9312 16680
rect 9364 16668 9370 16720
rect 9398 16668 9404 16720
rect 9456 16708 9462 16720
rect 13832 16708 13860 16748
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 19702 16776 19708 16788
rect 19076 16748 19708 16776
rect 9456 16680 13860 16708
rect 14369 16711 14427 16717
rect 9456 16668 9462 16680
rect 10520 16649 10548 16680
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 14550 16708 14556 16720
rect 14415 16680 14556 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 14550 16668 14556 16680
rect 14608 16668 14614 16720
rect 15010 16668 15016 16720
rect 15068 16668 15074 16720
rect 15562 16668 15568 16720
rect 15620 16708 15626 16720
rect 19076 16708 19104 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 20128 16748 20760 16776
rect 20128 16736 20134 16748
rect 15620 16680 19104 16708
rect 20732 16708 20760 16748
rect 23750 16736 23756 16788
rect 23808 16776 23814 16788
rect 30190 16776 30196 16788
rect 23808 16748 30196 16776
rect 23808 16736 23814 16748
rect 30190 16736 30196 16748
rect 30248 16736 30254 16788
rect 22002 16708 22008 16720
rect 20732 16680 22008 16708
rect 15620 16668 15626 16680
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 25682 16708 25688 16720
rect 25148 16680 25688 16708
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 8260 16612 8309 16640
rect 8260 16600 8266 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 10505 16643 10563 16649
rect 8527 16612 10364 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 4172 16544 4844 16572
rect 4065 16535 4123 16541
rect 1210 16464 1216 16516
rect 1268 16504 1274 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1268 16476 2513 16504
rect 1268 16464 1274 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 2501 16467 2559 16473
rect 4080 16436 4108 16535
rect 4816 16504 4844 16544
rect 4890 16532 4896 16584
rect 4948 16532 4954 16584
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 5000 16544 9413 16572
rect 5000 16504 5028 16544
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9401 16535 9459 16541
rect 4816 16476 5028 16504
rect 5718 16464 5724 16516
rect 5776 16504 5782 16516
rect 5905 16507 5963 16513
rect 5905 16504 5917 16507
rect 5776 16476 5917 16504
rect 5776 16464 5782 16476
rect 5905 16473 5917 16476
rect 5951 16473 5963 16507
rect 7282 16504 7288 16516
rect 5905 16467 5963 16473
rect 6012 16476 7288 16504
rect 6012 16436 6040 16476
rect 7282 16464 7288 16476
rect 7340 16464 7346 16516
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 7800 16476 8432 16504
rect 7800 16464 7806 16476
rect 4080 16408 6040 16436
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 6730 16436 6736 16448
rect 6687 16408 6736 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6972 16408 7021 16436
rect 6972 16396 6978 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7009 16399 7067 16405
rect 8202 16396 8208 16448
rect 8260 16396 8266 16448
rect 8404 16436 8432 16476
rect 9214 16464 9220 16516
rect 9272 16464 9278 16516
rect 10336 16504 10364 16612
rect 10505 16609 10517 16643
rect 10551 16609 10563 16643
rect 10505 16603 10563 16609
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 10410 16532 10416 16584
rect 10468 16532 10474 16584
rect 10704 16572 10732 16603
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 11701 16643 11759 16649
rect 11701 16640 11713 16643
rect 11664 16612 11713 16640
rect 11664 16600 11670 16612
rect 11701 16609 11713 16612
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 10962 16572 10968 16584
rect 10704 16544 10968 16572
rect 10704 16504 10732 16544
rect 10962 16532 10968 16544
rect 11020 16572 11026 16584
rect 11900 16572 11928 16603
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 12584 16612 12725 16640
rect 12584 16600 12590 16612
rect 12713 16609 12725 16612
rect 12759 16640 12771 16643
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 12759 16612 13461 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 13449 16609 13461 16612
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16640 13691 16643
rect 14274 16640 14280 16652
rect 13679 16612 14280 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 14516 16612 15485 16640
rect 14516 16600 14522 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 15746 16640 15752 16652
rect 15703 16612 15752 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 16393 16643 16451 16649
rect 16393 16640 16405 16643
rect 16356 16612 16405 16640
rect 16356 16600 16362 16612
rect 16393 16609 16405 16612
rect 16439 16609 16451 16643
rect 16393 16603 16451 16609
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16640 16819 16643
rect 17218 16640 17224 16652
rect 16807 16612 17224 16640
rect 16807 16609 16819 16612
rect 16761 16603 16819 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 18693 16643 18751 16649
rect 18693 16640 18705 16643
rect 17328 16612 18705 16640
rect 11020 16544 11928 16572
rect 11020 16532 11026 16544
rect 9324 16476 10088 16504
rect 10336 16476 10732 16504
rect 11609 16507 11667 16513
rect 9324 16436 9352 16476
rect 10060 16445 10088 16476
rect 11609 16473 11621 16507
rect 11655 16504 11667 16507
rect 11790 16504 11796 16516
rect 11655 16476 11796 16504
rect 11655 16473 11667 16476
rect 11609 16467 11667 16473
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 11900 16504 11928 16544
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 15286 16572 15292 16584
rect 14599 16544 15292 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 15378 16532 15384 16584
rect 15436 16532 15442 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 17328 16572 17356 16612
rect 18693 16609 18705 16612
rect 18739 16609 18751 16643
rect 18693 16603 18751 16609
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20438 16640 20444 16652
rect 19751 16612 20444 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 20772 16612 22477 16640
rect 20772 16600 20778 16612
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22646 16600 22652 16652
rect 22704 16600 22710 16652
rect 23750 16600 23756 16652
rect 23808 16600 23814 16652
rect 25038 16600 25044 16652
rect 25096 16640 25102 16652
rect 25148 16649 25176 16680
rect 25682 16668 25688 16680
rect 25740 16668 25746 16720
rect 25958 16668 25964 16720
rect 26016 16708 26022 16720
rect 26016 16680 28488 16708
rect 26016 16668 26022 16680
rect 25133 16643 25191 16649
rect 25133 16640 25145 16643
rect 25096 16612 25145 16640
rect 25096 16600 25102 16612
rect 25133 16609 25145 16612
rect 25179 16609 25191 16643
rect 25133 16603 25191 16609
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16640 25375 16643
rect 25774 16640 25780 16652
rect 25363 16612 25780 16640
rect 25363 16609 25375 16612
rect 25317 16603 25375 16609
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 25866 16600 25872 16652
rect 25924 16640 25930 16652
rect 26970 16640 26976 16652
rect 25924 16612 26976 16640
rect 25924 16600 25930 16612
rect 26970 16600 26976 16612
rect 27028 16600 27034 16652
rect 27062 16600 27068 16652
rect 27120 16600 27126 16652
rect 27246 16600 27252 16652
rect 27304 16600 27310 16652
rect 27798 16600 27804 16652
rect 27856 16640 27862 16652
rect 28258 16640 28264 16652
rect 27856 16612 28264 16640
rect 27856 16600 27862 16612
rect 28258 16600 28264 16612
rect 28316 16600 28322 16652
rect 28460 16649 28488 16680
rect 28445 16643 28503 16649
rect 28445 16609 28457 16643
rect 28491 16640 28503 16643
rect 28994 16640 29000 16652
rect 28491 16612 29000 16640
rect 28491 16609 28503 16612
rect 28445 16603 28503 16609
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 15620 16544 17356 16572
rect 17589 16575 17647 16581
rect 15620 16532 15626 16544
rect 17589 16541 17601 16575
rect 17635 16572 17647 16575
rect 17770 16572 17776 16584
rect 17635 16544 17776 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18230 16532 18236 16584
rect 18288 16532 18294 16584
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16572 22431 16575
rect 23290 16572 23296 16584
rect 22419 16544 23296 16572
rect 22419 16541 22431 16544
rect 22373 16535 22431 16541
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 23658 16572 23664 16584
rect 23615 16544 23664 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 23658 16532 23664 16544
rect 23716 16572 23722 16584
rect 24210 16572 24216 16584
rect 23716 16544 24216 16572
rect 23716 16532 23722 16544
rect 24210 16532 24216 16544
rect 24268 16532 24274 16584
rect 24486 16532 24492 16584
rect 24544 16572 24550 16584
rect 24544 16544 25452 16572
rect 24544 16532 24550 16544
rect 17954 16504 17960 16516
rect 11900 16476 17960 16504
rect 17954 16464 17960 16476
rect 18012 16464 18018 16516
rect 19978 16504 19984 16516
rect 18708 16476 19984 16504
rect 8404 16408 9352 16436
rect 10045 16439 10103 16445
rect 10045 16405 10057 16439
rect 10091 16405 10103 16439
rect 10045 16399 10103 16405
rect 10502 16396 10508 16448
rect 10560 16436 10566 16448
rect 11241 16439 11299 16445
rect 11241 16436 11253 16439
rect 10560 16408 11253 16436
rect 10560 16396 10566 16408
rect 11241 16405 11253 16408
rect 11287 16405 11299 16439
rect 11808 16436 11836 16464
rect 12253 16439 12311 16445
rect 12253 16436 12265 16439
rect 11808 16408 12265 16436
rect 11241 16399 11299 16405
rect 12253 16405 12265 16408
rect 12299 16405 12311 16439
rect 12253 16399 12311 16405
rect 12989 16439 13047 16445
rect 12989 16405 13001 16439
rect 13035 16436 13047 16439
rect 13170 16436 13176 16448
rect 13035 16408 13176 16436
rect 13035 16405 13047 16408
rect 12989 16399 13047 16405
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 13354 16396 13360 16448
rect 13412 16396 13418 16448
rect 14366 16396 14372 16448
rect 14424 16436 14430 16448
rect 15562 16436 15568 16448
rect 14424 16408 15568 16436
rect 14424 16396 14430 16408
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 16117 16439 16175 16445
rect 16117 16405 16129 16439
rect 16163 16436 16175 16439
rect 16206 16436 16212 16448
rect 16163 16408 16212 16436
rect 16163 16405 16175 16408
rect 16117 16399 16175 16405
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 16301 16439 16359 16445
rect 16301 16405 16313 16439
rect 16347 16436 16359 16439
rect 16482 16436 16488 16448
rect 16347 16408 16488 16436
rect 16347 16405 16359 16408
rect 16301 16399 16359 16405
rect 16482 16396 16488 16408
rect 16540 16396 16546 16448
rect 16758 16396 16764 16448
rect 16816 16436 16822 16448
rect 17405 16439 17463 16445
rect 17405 16436 17417 16439
rect 16816 16408 17417 16436
rect 16816 16396 16822 16408
rect 17405 16405 17417 16408
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18049 16439 18107 16445
rect 18049 16405 18061 16439
rect 18095 16436 18107 16439
rect 18708 16436 18736 16476
rect 19978 16464 19984 16476
rect 20036 16464 20042 16516
rect 21082 16504 21088 16516
rect 20930 16476 21088 16504
rect 21082 16464 21088 16476
rect 21140 16464 21146 16516
rect 21453 16507 21511 16513
rect 21453 16473 21465 16507
rect 21499 16473 21511 16507
rect 21453 16467 21511 16473
rect 18095 16408 18736 16436
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 18966 16396 18972 16448
rect 19024 16436 19030 16448
rect 21468 16436 21496 16467
rect 23382 16464 23388 16516
rect 23440 16504 23446 16516
rect 25424 16504 25452 16544
rect 25590 16532 25596 16584
rect 25648 16572 25654 16584
rect 25648 16544 26740 16572
rect 25648 16532 25654 16544
rect 23440 16476 24716 16504
rect 25424 16476 26648 16504
rect 23440 16464 23446 16476
rect 19024 16408 21496 16436
rect 19024 16396 19030 16408
rect 21542 16396 21548 16448
rect 21600 16436 21606 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 21600 16408 22017 16436
rect 21600 16396 21606 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 22462 16396 22468 16448
rect 22520 16436 22526 16448
rect 23201 16439 23259 16445
rect 23201 16436 23213 16439
rect 22520 16408 23213 16436
rect 22520 16396 22526 16408
rect 23201 16405 23213 16408
rect 23247 16405 23259 16439
rect 23201 16399 23259 16405
rect 23661 16439 23719 16445
rect 23661 16405 23673 16439
rect 23707 16436 23719 16439
rect 23842 16436 23848 16448
rect 23707 16408 23848 16436
rect 23707 16405 23719 16408
rect 23661 16399 23719 16405
rect 23842 16396 23848 16408
rect 23900 16436 23906 16448
rect 24578 16436 24584 16448
rect 23900 16408 24584 16436
rect 23900 16396 23906 16408
rect 24578 16396 24584 16408
rect 24636 16396 24642 16448
rect 24688 16445 24716 16476
rect 24673 16439 24731 16445
rect 24673 16405 24685 16439
rect 24719 16405 24731 16439
rect 24673 16399 24731 16405
rect 25041 16439 25099 16445
rect 25041 16405 25053 16439
rect 25087 16436 25099 16439
rect 25130 16436 25136 16448
rect 25087 16408 25136 16436
rect 25087 16405 25099 16408
rect 25041 16399 25099 16405
rect 25130 16396 25136 16408
rect 25188 16436 25194 16448
rect 25866 16436 25872 16448
rect 25188 16408 25872 16436
rect 25188 16396 25194 16408
rect 25866 16396 25872 16408
rect 25924 16396 25930 16448
rect 26620 16445 26648 16476
rect 26605 16439 26663 16445
rect 26605 16405 26617 16439
rect 26651 16405 26663 16439
rect 26712 16436 26740 16544
rect 27614 16532 27620 16584
rect 27672 16572 27678 16584
rect 28169 16575 28227 16581
rect 28169 16572 28181 16575
rect 27672 16544 28181 16572
rect 27672 16532 27678 16544
rect 28169 16541 28181 16544
rect 28215 16541 28227 16575
rect 28169 16535 28227 16541
rect 26973 16507 27031 16513
rect 26973 16473 26985 16507
rect 27019 16504 27031 16507
rect 28442 16504 28448 16516
rect 27019 16476 28448 16504
rect 27019 16473 27031 16476
rect 26973 16467 27031 16473
rect 28442 16464 28448 16476
rect 28500 16464 28506 16516
rect 27801 16439 27859 16445
rect 27801 16436 27813 16439
rect 26712 16408 27813 16436
rect 26605 16399 26663 16405
rect 27801 16405 27813 16408
rect 27847 16405 27859 16439
rect 27801 16399 27859 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 3878 16192 3884 16244
rect 3936 16232 3942 16244
rect 4890 16232 4896 16244
rect 3936 16204 4896 16232
rect 3936 16192 3942 16204
rect 4890 16192 4896 16204
rect 4948 16232 4954 16244
rect 5626 16232 5632 16244
rect 4948 16204 5632 16232
rect 4948 16192 4954 16204
rect 5626 16192 5632 16204
rect 5684 16192 5690 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 5994 16232 6000 16244
rect 5767 16204 6000 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 7374 16232 7380 16244
rect 7331 16204 7380 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 12526 16232 12532 16244
rect 7852 16204 12532 16232
rect 4338 16124 4344 16176
rect 4396 16124 4402 16176
rect 5442 16124 5448 16176
rect 5500 16164 5506 16176
rect 6638 16164 6644 16176
rect 5500 16136 6644 16164
rect 5500 16124 5506 16136
rect 6638 16124 6644 16136
rect 6696 16124 6702 16176
rect 7098 16124 7104 16176
rect 7156 16164 7162 16176
rect 7745 16167 7803 16173
rect 7745 16164 7757 16167
rect 7156 16136 7757 16164
rect 7156 16124 7162 16136
rect 7745 16133 7757 16136
rect 7791 16133 7803 16167
rect 7745 16127 7803 16133
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 1854 16096 1860 16108
rect 1811 16068 1860 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 5626 16056 5632 16108
rect 5684 16056 5690 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 7064 16068 7665 16096
rect 7064 16056 7070 16068
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7852 16096 7880 16204
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 13722 16192 13728 16244
rect 13780 16192 13786 16244
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16356 16204 16773 16232
rect 16356 16192 16362 16204
rect 8754 16164 8760 16176
rect 7653 16059 7711 16065
rect 7760 16068 7880 16096
rect 8036 16136 8760 16164
rect 1118 15988 1124 16040
rect 1176 16028 1182 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1176 16000 2053 16028
rect 1176 15988 1182 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 6086 16028 6092 16040
rect 5951 16000 6092 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6086 15988 6092 16000
rect 6144 16028 6150 16040
rect 6362 16028 6368 16040
rect 6144 16000 6368 16028
rect 6144 15988 6150 16000
rect 6362 15988 6368 16000
rect 6420 15988 6426 16040
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 7558 16028 7564 16040
rect 6687 16000 7564 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 7558 15988 7564 16000
rect 7616 15988 7622 16040
rect 7760 16028 7788 16068
rect 7668 16000 7788 16028
rect 7929 16031 7987 16037
rect 4430 15920 4436 15972
rect 4488 15960 4494 15972
rect 7668 15960 7696 16000
rect 7929 15997 7941 16031
rect 7975 16028 7987 16031
rect 8036 16028 8064 16136
rect 8754 16124 8760 16136
rect 8812 16124 8818 16176
rect 10042 16164 10048 16176
rect 9982 16136 10048 16164
rect 10042 16124 10048 16136
rect 10100 16164 10106 16176
rect 12250 16164 12256 16176
rect 10100 16136 12256 16164
rect 10100 16124 10106 16136
rect 12250 16124 12256 16136
rect 12308 16164 12314 16176
rect 14645 16167 14703 16173
rect 12308 16136 12742 16164
rect 12308 16124 12314 16136
rect 14645 16133 14657 16167
rect 14691 16164 14703 16167
rect 16482 16164 16488 16176
rect 14691 16136 16488 16164
rect 14691 16133 14703 16136
rect 14645 16127 14703 16133
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 8478 16056 8484 16108
rect 8536 16056 8542 16108
rect 10594 16056 10600 16108
rect 10652 16056 10658 16108
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 11149 16099 11207 16105
rect 11020 16068 11100 16096
rect 11020 16056 11026 16068
rect 8202 16028 8208 16040
rect 7975 16000 8064 16028
rect 8128 16000 8208 16028
rect 7975 15997 7987 16000
rect 7929 15991 7987 15997
rect 8128 15960 8156 16000
rect 8202 15988 8208 16000
rect 8260 16028 8266 16040
rect 8757 16031 8815 16037
rect 8757 16028 8769 16031
rect 8260 16000 8769 16028
rect 8260 15988 8266 16000
rect 8757 15997 8769 16000
rect 8803 16028 8815 16031
rect 9950 16028 9956 16040
rect 8803 16000 9956 16028
rect 8803 15997 8815 16000
rect 8757 15991 8815 15997
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 10229 16031 10287 16037
rect 10229 16028 10241 16031
rect 10192 16000 10241 16028
rect 10192 15988 10198 16000
rect 10229 15997 10241 16000
rect 10275 16028 10287 16031
rect 10870 16028 10876 16040
rect 10275 16000 10876 16028
rect 10275 15997 10287 16000
rect 10229 15991 10287 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 11072 16028 11100 16068
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11790 16096 11796 16108
rect 11195 16068 11796 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11790 16056 11796 16068
rect 11848 16056 11854 16108
rect 11974 16056 11980 16108
rect 12032 16056 12038 16108
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 14918 16096 14924 16108
rect 14783 16068 14924 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 14918 16056 14924 16068
rect 14976 16056 14982 16108
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16390 16096 16396 16108
rect 16347 16068 16396 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16592 16096 16620 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 16761 16195 16819 16201
rect 17126 16192 17132 16244
rect 17184 16192 17190 16244
rect 17405 16235 17463 16241
rect 17405 16201 17417 16235
rect 17451 16232 17463 16235
rect 17586 16232 17592 16244
rect 17451 16204 17592 16232
rect 17451 16201 17463 16204
rect 17405 16195 17463 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 17862 16192 17868 16244
rect 17920 16192 17926 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 20441 16235 20499 16241
rect 20441 16232 20453 16235
rect 18748 16204 20453 16232
rect 18748 16192 18754 16204
rect 20441 16201 20453 16204
rect 20487 16201 20499 16235
rect 20441 16195 20499 16201
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 21450 16232 21456 16244
rect 21232 16204 21456 16232
rect 21232 16192 21238 16204
rect 21450 16192 21456 16204
rect 21508 16232 21514 16244
rect 21508 16204 24900 16232
rect 21508 16192 21514 16204
rect 16666 16124 16672 16176
rect 16724 16164 16730 16176
rect 16724 16136 18092 16164
rect 16724 16124 16730 16136
rect 17586 16096 17592 16108
rect 16592 16068 17592 16096
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 11238 16028 11244 16040
rect 11072 16000 11244 16028
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 11422 15988 11428 16040
rect 11480 16028 11486 16040
rect 11698 16028 11704 16040
rect 11480 16000 11704 16028
rect 11480 15988 11486 16000
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 12250 15988 12256 16040
rect 12308 15988 12314 16040
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 14829 16031 14887 16037
rect 12676 16000 14412 16028
rect 12676 15988 12682 16000
rect 4488 15932 7696 15960
rect 7760 15932 8156 15960
rect 9968 15960 9996 15988
rect 10778 15960 10784 15972
rect 9968 15932 10784 15960
rect 4488 15920 4494 15932
rect 5258 15852 5264 15904
rect 5316 15852 5322 15904
rect 5810 15852 5816 15904
rect 5868 15892 5874 15904
rect 7760 15892 7788 15932
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 10962 15920 10968 15972
rect 11020 15920 11026 15972
rect 14277 15963 14335 15969
rect 14277 15960 14289 15963
rect 13372 15932 14289 15960
rect 5868 15864 7788 15892
rect 5868 15852 5874 15864
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 9858 15892 9864 15904
rect 8812 15864 9864 15892
rect 8812 15852 8818 15864
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 13372 15892 13400 15932
rect 14277 15929 14289 15932
rect 14323 15929 14335 15963
rect 14384 15960 14412 16000
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14936 16028 14964 16056
rect 14936 16000 15056 16028
rect 14829 15991 14887 15997
rect 14844 15960 14872 15991
rect 14384 15932 14872 15960
rect 15028 15960 15056 16000
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 15562 15988 15568 16040
rect 15620 16028 15626 16040
rect 17788 16028 17816 16059
rect 15620 16000 17816 16028
rect 17957 16031 18015 16037
rect 15620 15988 15626 16000
rect 17957 15997 17969 16031
rect 18003 15997 18015 16031
rect 18064 16028 18092 16136
rect 18874 16124 18880 16176
rect 18932 16164 18938 16176
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 18932 16136 19717 16164
rect 18932 16124 18938 16136
rect 19705 16133 19717 16136
rect 19751 16164 19763 16167
rect 20533 16167 20591 16173
rect 20533 16164 20545 16167
rect 19751 16136 20545 16164
rect 19751 16133 19763 16136
rect 19705 16127 19763 16133
rect 20533 16133 20545 16136
rect 20579 16133 20591 16167
rect 24872 16164 24900 16204
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 26605 16235 26663 16241
rect 26605 16232 26617 16235
rect 25004 16204 26617 16232
rect 25004 16192 25010 16204
rect 26605 16201 26617 16204
rect 26651 16201 26663 16235
rect 26605 16195 26663 16201
rect 27614 16192 27620 16244
rect 27672 16232 27678 16244
rect 27709 16235 27767 16241
rect 27709 16232 27721 16235
rect 27672 16204 27721 16232
rect 27672 16192 27678 16204
rect 27709 16201 27721 16204
rect 27755 16232 27767 16235
rect 27798 16232 27804 16244
rect 27755 16204 27804 16232
rect 27755 16201 27767 16204
rect 27709 16195 27767 16201
rect 27798 16192 27804 16204
rect 27856 16192 27862 16244
rect 25406 16164 25412 16176
rect 20533 16127 20591 16133
rect 20640 16136 24808 16164
rect 24872 16136 25412 16164
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16096 18659 16099
rect 19150 16096 19156 16108
rect 18647 16068 19156 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 20070 16096 20076 16108
rect 19484 16068 20076 16096
rect 19484 16056 19490 16068
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 20640 16037 20668 16136
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16096 21511 16099
rect 22281 16099 22339 16105
rect 21499 16068 22232 16096
rect 21499 16065 21511 16068
rect 21453 16059 21511 16065
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18064 16000 18889 16028
rect 17957 15991 18015 15997
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 15028 15932 16988 15960
rect 14277 15923 14335 15929
rect 11756 15864 13400 15892
rect 11756 15852 11762 15864
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 16960 15901 16988 15932
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 17972 15960 18000 15991
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 21692 16000 22017 16028
rect 21692 15988 21698 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22204 16028 22232 16068
rect 22281 16065 22293 16099
rect 22327 16096 22339 16099
rect 22370 16096 22376 16108
rect 22327 16068 22376 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 23658 16056 23664 16108
rect 23716 16096 23722 16108
rect 24305 16099 24363 16105
rect 24305 16096 24317 16099
rect 23716 16068 24317 16096
rect 23716 16056 23722 16068
rect 24305 16065 24317 16068
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 24578 16056 24584 16108
rect 24636 16056 24642 16108
rect 23753 16031 23811 16037
rect 22204 16000 22968 16028
rect 22005 15991 22063 15997
rect 17552 15932 18000 15960
rect 20073 15963 20131 15969
rect 17552 15920 17558 15932
rect 20073 15929 20085 15963
rect 20119 15960 20131 15963
rect 22830 15960 22836 15972
rect 20119 15932 22836 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 22830 15920 22836 15932
rect 22888 15920 22894 15972
rect 22940 15960 22968 16000
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 23842 16028 23848 16040
rect 23799 16000 23848 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 23937 16031 23995 16037
rect 23937 15997 23949 16031
rect 23983 16028 23995 16031
rect 24026 16028 24032 16040
rect 23983 16000 24032 16028
rect 23983 15997 23995 16000
rect 23937 15991 23995 15997
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24780 16028 24808 16136
rect 25406 16124 25412 16136
rect 25464 16124 25470 16176
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 26234 16056 26240 16108
rect 26292 16096 26298 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26292 16068 26985 16096
rect 26292 16056 26298 16068
rect 26973 16065 26985 16068
rect 27019 16096 27031 16099
rect 27062 16096 27068 16108
rect 27019 16068 27068 16096
rect 27019 16065 27031 16068
rect 26973 16059 27031 16065
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24780 16000 25145 16028
rect 25133 15997 25145 16000
rect 25179 16028 25191 16031
rect 27246 16028 27252 16040
rect 25179 16000 27252 16028
rect 25179 15997 25191 16000
rect 25133 15991 25191 15997
rect 27246 15988 27252 16000
rect 27304 15988 27310 16040
rect 22940 15932 24624 15960
rect 16117 15895 16175 15901
rect 16117 15892 16129 15895
rect 14056 15864 16129 15892
rect 14056 15852 14062 15864
rect 16117 15861 16129 15864
rect 16163 15861 16175 15895
rect 16117 15855 16175 15861
rect 16945 15895 17003 15901
rect 16945 15861 16957 15895
rect 16991 15892 17003 15895
rect 20162 15892 20168 15904
rect 16991 15864 20168 15892
rect 16991 15861 17003 15864
rect 16945 15855 17003 15861
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 23293 15895 23351 15901
rect 23293 15892 23305 15895
rect 22244 15864 23305 15892
rect 22244 15852 22250 15864
rect 23293 15861 23305 15864
rect 23339 15861 23351 15895
rect 24596 15892 24624 15932
rect 25222 15892 25228 15904
rect 24596 15864 25228 15892
rect 23293 15855 23351 15861
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 6270 15688 6276 15700
rect 5500 15660 6276 15688
rect 5500 15648 5506 15660
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7248 15660 7849 15688
rect 7248 15648 7254 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8260 15660 8432 15688
rect 8260 15648 8266 15660
rect 3421 15623 3479 15629
rect 3421 15589 3433 15623
rect 3467 15620 3479 15623
rect 3786 15620 3792 15632
rect 3467 15592 3792 15620
rect 3467 15589 3479 15592
rect 3421 15583 3479 15589
rect 3786 15580 3792 15592
rect 3844 15620 3850 15632
rect 3844 15592 7052 15620
rect 3844 15580 3850 15592
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 3418 15484 3424 15496
rect 1811 15456 3424 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 4062 15484 4068 15496
rect 3651 15456 4068 15484
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4632 15484 4660 15515
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5592 15524 5641 15552
rect 5592 15512 5598 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15521 5779 15555
rect 5721 15515 5779 15521
rect 5736 15484 5764 15515
rect 5810 15512 5816 15564
rect 5868 15552 5874 15564
rect 6917 15555 6975 15561
rect 6917 15552 6929 15555
rect 5868 15524 6929 15552
rect 5868 15512 5874 15524
rect 6917 15521 6929 15524
rect 6963 15521 6975 15555
rect 7024 15552 7052 15592
rect 8404 15561 8432 15660
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8720 15660 9321 15688
rect 8720 15648 8726 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 9309 15651 9367 15657
rect 9769 15691 9827 15697
rect 9769 15657 9781 15691
rect 9815 15688 9827 15691
rect 10042 15688 10048 15700
rect 9815 15660 10048 15688
rect 9815 15657 9827 15660
rect 9769 15651 9827 15657
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 13354 15688 13360 15700
rect 10468 15660 13360 15688
rect 10468 15648 10474 15660
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 14734 15688 14740 15700
rect 14608 15660 14740 15688
rect 14608 15648 14614 15660
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 15841 15691 15899 15697
rect 15841 15657 15853 15691
rect 15887 15688 15899 15691
rect 15930 15688 15936 15700
rect 15887 15660 15936 15688
rect 15887 15657 15899 15660
rect 15841 15651 15899 15657
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 17828 15660 21588 15688
rect 17828 15648 17834 15660
rect 8570 15580 8576 15632
rect 8628 15620 8634 15632
rect 9122 15620 9128 15632
rect 8628 15592 9128 15620
rect 8628 15580 8634 15592
rect 9122 15580 9128 15592
rect 9180 15580 9186 15632
rect 9214 15580 9220 15632
rect 9272 15620 9278 15632
rect 9272 15592 11652 15620
rect 9272 15580 9278 15592
rect 8297 15555 8355 15561
rect 8297 15552 8309 15555
rect 7024 15524 8309 15552
rect 6917 15515 6975 15521
rect 8297 15521 8309 15524
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 9398 15552 9404 15564
rect 8536 15524 9404 15552
rect 8536 15512 8542 15524
rect 9398 15512 9404 15524
rect 9456 15512 9462 15564
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 10410 15552 10416 15564
rect 10275 15524 10416 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 10410 15512 10416 15524
rect 10468 15512 10474 15564
rect 10778 15512 10784 15564
rect 10836 15552 10842 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 10836 15524 11437 15552
rect 10836 15512 10842 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11624 15552 11652 15592
rect 12066 15580 12072 15632
rect 12124 15580 12130 15632
rect 13541 15623 13599 15629
rect 13541 15620 13553 15623
rect 12176 15592 13553 15620
rect 12176 15552 12204 15592
rect 13541 15589 13553 15592
rect 13587 15589 13599 15623
rect 13541 15583 13599 15589
rect 13630 15580 13636 15632
rect 13688 15620 13694 15632
rect 14461 15623 14519 15629
rect 14461 15620 14473 15623
rect 13688 15592 14473 15620
rect 13688 15580 13694 15592
rect 14461 15589 14473 15592
rect 14507 15589 14519 15623
rect 14461 15583 14519 15589
rect 19886 15580 19892 15632
rect 19944 15580 19950 15632
rect 21560 15620 21588 15660
rect 21634 15648 21640 15700
rect 21692 15688 21698 15700
rect 22465 15691 22523 15697
rect 22465 15688 22477 15691
rect 21692 15660 22477 15688
rect 21692 15648 21698 15660
rect 22465 15657 22477 15660
rect 22511 15657 22523 15691
rect 22465 15651 22523 15657
rect 24489 15691 24547 15697
rect 24489 15657 24501 15691
rect 24535 15688 24547 15691
rect 24578 15688 24584 15700
rect 24535 15660 24584 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 29730 15688 29736 15700
rect 25516 15660 29736 15688
rect 25516 15620 25544 15660
rect 29730 15648 29736 15660
rect 29788 15648 29794 15700
rect 26329 15623 26387 15629
rect 26329 15620 26341 15623
rect 21560 15592 25544 15620
rect 25608 15592 26341 15620
rect 11624 15524 12204 15552
rect 12713 15555 12771 15561
rect 11425 15515 11483 15521
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12802 15552 12808 15564
rect 12759 15524 12808 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 14366 15512 14372 15564
rect 14424 15552 14430 15564
rect 15013 15555 15071 15561
rect 15013 15552 15025 15555
rect 14424 15524 15025 15552
rect 14424 15512 14430 15524
rect 15013 15521 15025 15524
rect 15059 15521 15071 15555
rect 15013 15515 15071 15521
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 4632 15456 5672 15484
rect 5736 15456 6500 15484
rect 5537 15419 5595 15425
rect 5537 15416 5549 15419
rect 3988 15388 5549 15416
rect 3988 15357 4016 15388
rect 5537 15385 5549 15388
rect 5583 15385 5595 15419
rect 5537 15379 5595 15385
rect 3973 15351 4031 15357
rect 3973 15317 3985 15351
rect 4019 15317 4031 15351
rect 3973 15311 4031 15317
rect 4338 15308 4344 15360
rect 4396 15308 4402 15360
rect 5166 15308 5172 15360
rect 5224 15308 5230 15360
rect 5644 15348 5672 15456
rect 6086 15348 6092 15360
rect 5644 15320 6092 15348
rect 6086 15308 6092 15320
rect 6144 15308 6150 15360
rect 6362 15308 6368 15360
rect 6420 15308 6426 15360
rect 6472 15348 6500 15456
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6696 15456 6837 15484
rect 6696 15444 6702 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7374 15444 7380 15496
rect 7432 15484 7438 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 7432 15456 7481 15484
rect 7432 15444 7438 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 8110 15444 8116 15496
rect 8168 15484 8174 15496
rect 12437 15487 12495 15493
rect 12437 15484 12449 15487
rect 8168 15456 12449 15484
rect 8168 15444 8174 15456
rect 12437 15453 12449 15456
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13722 15484 13728 15496
rect 13311 15456 13728 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 15470 15484 15476 15496
rect 14875 15456 15476 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 6733 15419 6791 15425
rect 6733 15385 6745 15419
rect 6779 15416 6791 15419
rect 8478 15416 8484 15428
rect 6779 15388 8484 15416
rect 6779 15385 6791 15388
rect 6733 15379 6791 15385
rect 8478 15376 8484 15388
rect 8536 15376 8542 15428
rect 9214 15376 9220 15428
rect 9272 15376 9278 15428
rect 11330 15416 11336 15428
rect 9876 15388 11336 15416
rect 9876 15360 9904 15388
rect 11330 15376 11336 15388
rect 11388 15376 11394 15428
rect 14921 15419 14979 15425
rect 14921 15416 14933 15419
rect 13740 15388 14933 15416
rect 13740 15360 13768 15388
rect 14921 15385 14933 15388
rect 14967 15385 14979 15419
rect 14921 15379 14979 15385
rect 16022 15376 16028 15428
rect 16080 15416 16086 15428
rect 16500 15416 16528 15515
rect 20070 15512 20076 15564
rect 20128 15552 20134 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 20128 15524 20269 15552
rect 20128 15512 20134 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21140 15524 21680 15552
rect 21140 15512 21146 15524
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 19610 15444 19616 15496
rect 19668 15444 19674 15496
rect 21652 15484 21680 15524
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22741 15555 22799 15561
rect 22741 15552 22753 15555
rect 22152 15524 22753 15552
rect 22152 15512 22158 15524
rect 22741 15521 22753 15524
rect 22787 15552 22799 15555
rect 22787 15524 23152 15552
rect 22787 15521 22799 15524
rect 22741 15515 22799 15521
rect 22370 15484 22376 15496
rect 21652 15470 22376 15484
rect 21666 15456 22376 15470
rect 22370 15444 22376 15456
rect 22428 15444 22434 15496
rect 23124 15493 23152 15524
rect 25608 15496 25636 15592
rect 26329 15589 26341 15592
rect 26375 15620 26387 15623
rect 26970 15620 26976 15632
rect 26375 15592 26976 15620
rect 26375 15589 26387 15592
rect 26329 15583 26387 15589
rect 26970 15580 26976 15592
rect 27028 15620 27034 15632
rect 34514 15620 34520 15632
rect 27028 15592 34520 15620
rect 27028 15580 27034 15592
rect 34514 15580 34520 15592
rect 34572 15580 34578 15632
rect 25774 15512 25780 15564
rect 25832 15512 25838 15564
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15484 23167 15487
rect 23290 15484 23296 15496
rect 23155 15456 23296 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 25590 15444 25596 15496
rect 25648 15444 25654 15496
rect 17310 15416 17316 15428
rect 16080 15388 16344 15416
rect 16500 15388 17316 15416
rect 16080 15376 16086 15388
rect 7374 15348 7380 15360
rect 6472 15320 7380 15348
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 7466 15308 7472 15360
rect 7524 15348 7530 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 7524 15320 8217 15348
rect 7524 15308 7530 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8205 15311 8263 15317
rect 8570 15308 8576 15360
rect 8628 15348 8634 15360
rect 9582 15348 9588 15360
rect 8628 15320 9588 15348
rect 8628 15308 8634 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 10870 15308 10876 15360
rect 10928 15308 10934 15360
rect 11241 15351 11299 15357
rect 11241 15317 11253 15351
rect 11287 15348 11299 15351
rect 11422 15348 11428 15360
rect 11287 15320 11428 15348
rect 11287 15317 11299 15320
rect 11241 15311 11299 15317
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 13722 15308 13728 15360
rect 13780 15308 13786 15360
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 13964 15320 14105 15348
rect 13964 15308 13970 15320
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 16316 15357 16344 15388
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17586 15376 17592 15428
rect 17644 15416 17650 15428
rect 17644 15388 17802 15416
rect 17644 15376 17650 15388
rect 20254 15376 20260 15428
rect 20312 15416 20318 15428
rect 20533 15419 20591 15425
rect 20533 15416 20545 15419
rect 20312 15388 20545 15416
rect 20312 15376 20318 15388
rect 20533 15385 20545 15388
rect 20579 15385 20591 15419
rect 22646 15416 22652 15428
rect 20533 15379 20591 15385
rect 21836 15388 22652 15416
rect 16209 15351 16267 15357
rect 16209 15348 16221 15351
rect 15528 15320 16221 15348
rect 15528 15308 15534 15320
rect 16209 15317 16221 15320
rect 16255 15317 16267 15351
rect 16209 15311 16267 15317
rect 16301 15351 16359 15357
rect 16301 15317 16313 15351
rect 16347 15348 16359 15351
rect 16390 15348 16396 15360
rect 16347 15320 16396 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 17460 15320 18797 15348
rect 17460 15308 17466 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 19392 15320 19441 15348
rect 19392 15308 19398 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 20548 15348 20576 15379
rect 21836 15348 21864 15388
rect 22646 15376 22652 15388
rect 22704 15416 22710 15428
rect 23566 15416 23572 15428
rect 22704 15388 23572 15416
rect 22704 15376 22710 15388
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 23934 15376 23940 15428
rect 23992 15376 23998 15428
rect 25406 15376 25412 15428
rect 25464 15416 25470 15428
rect 25685 15419 25743 15425
rect 25685 15416 25697 15419
rect 25464 15388 25697 15416
rect 25464 15376 25470 15388
rect 25685 15385 25697 15388
rect 25731 15416 25743 15419
rect 26326 15416 26332 15428
rect 25731 15388 26332 15416
rect 25731 15385 25743 15388
rect 25685 15379 25743 15385
rect 26326 15376 26332 15388
rect 26384 15416 26390 15428
rect 26421 15419 26479 15425
rect 26421 15416 26433 15419
rect 26384 15388 26433 15416
rect 26384 15376 26390 15388
rect 26421 15385 26433 15388
rect 26467 15416 26479 15419
rect 26467 15388 31754 15416
rect 26467 15385 26479 15388
rect 26421 15379 26479 15385
rect 20548 15320 21864 15348
rect 19429 15311 19487 15317
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21968 15320 22017 15348
rect 21968 15308 21974 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22005 15311 22063 15317
rect 22370 15308 22376 15360
rect 22428 15348 22434 15360
rect 23474 15348 23480 15360
rect 22428 15320 23480 15348
rect 22428 15308 22434 15320
rect 23474 15308 23480 15320
rect 23532 15348 23538 15360
rect 23842 15348 23848 15360
rect 23532 15320 23848 15348
rect 23532 15308 23538 15320
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 25222 15308 25228 15360
rect 25280 15308 25286 15360
rect 31726 15348 31754 15388
rect 40770 15348 40776 15360
rect 31726 15320 40776 15348
rect 40770 15308 40776 15320
rect 40828 15308 40834 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 3510 15104 3516 15156
rect 3568 15104 3574 15156
rect 4798 15104 4804 15156
rect 4856 15144 4862 15156
rect 5902 15144 5908 15156
rect 4856 15116 5908 15144
rect 4856 15104 4862 15116
rect 5902 15104 5908 15116
rect 5960 15104 5966 15156
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 6236 15116 8677 15144
rect 6236 15104 6242 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8665 15107 8723 15113
rect 9217 15147 9275 15153
rect 9217 15113 9229 15147
rect 9263 15113 9275 15147
rect 9217 15107 9275 15113
rect 4706 15076 4712 15088
rect 1780 15048 4712 15076
rect 1780 15017 1808 15048
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 5442 15036 5448 15088
rect 5500 15036 5506 15088
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 7653 15079 7711 15085
rect 7653 15076 7665 15079
rect 5776 15048 7665 15076
rect 5776 15036 5782 15048
rect 7653 15045 7665 15048
rect 7699 15045 7711 15079
rect 7653 15039 7711 15045
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 3694 14968 3700 15020
rect 3752 14968 3758 15020
rect 4154 14968 4160 15020
rect 4212 14968 4218 15020
rect 5902 14968 5908 15020
rect 5960 15008 5966 15020
rect 6638 15008 6644 15020
rect 5960 14980 6644 15008
rect 5960 14968 5966 14980
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 7668 15008 7696 15039
rect 7926 15008 7932 15020
rect 7668 14980 7932 15008
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8570 14968 8576 15020
rect 8628 14968 8634 15020
rect 9232 15008 9260 15107
rect 9306 15104 9312 15156
rect 9364 15104 9370 15156
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 9548 15116 10364 15144
rect 9548 15104 9554 15116
rect 9324 15076 9352 15104
rect 9677 15079 9735 15085
rect 9677 15076 9689 15079
rect 9324 15048 9689 15076
rect 9677 15045 9689 15048
rect 9723 15045 9735 15079
rect 9677 15039 9735 15045
rect 9306 15008 9312 15020
rect 9232 14980 9312 15008
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 10336 15008 10364 15116
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12492 15116 13001 15144
rect 12492 15104 12498 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 14826 15144 14832 15156
rect 12989 15107 13047 15113
rect 13096 15116 14832 15144
rect 10594 15036 10600 15088
rect 10652 15076 10658 15088
rect 10781 15079 10839 15085
rect 10781 15076 10793 15079
rect 10652 15048 10793 15076
rect 10652 15036 10658 15048
rect 10781 15045 10793 15048
rect 10827 15045 10839 15079
rect 10781 15039 10839 15045
rect 10873 15079 10931 15085
rect 10873 15045 10885 15079
rect 10919 15076 10931 15079
rect 10962 15076 10968 15088
rect 10919 15048 10968 15076
rect 10919 15045 10931 15048
rect 10873 15039 10931 15045
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11882 15008 11888 15020
rect 9631 14980 10272 15008
rect 10336 14980 11888 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 1118 14900 1124 14952
rect 1176 14940 1182 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1176 14912 2053 14940
rect 1176 14900 1182 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14940 4491 14943
rect 4798 14940 4804 14952
rect 4479 14912 4804 14940
rect 4479 14909 4491 14912
rect 4433 14903 4491 14909
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 5718 14900 5724 14952
rect 5776 14940 5782 14952
rect 6086 14940 6092 14952
rect 5776 14912 6092 14940
rect 5776 14900 5782 14912
rect 6086 14900 6092 14912
rect 6144 14900 6150 14952
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 7745 14943 7803 14949
rect 7745 14940 7757 14943
rect 6512 14912 7757 14940
rect 6512 14900 6518 14912
rect 7745 14909 7757 14912
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 6825 14875 6883 14881
rect 6825 14872 6837 14875
rect 5460 14844 6837 14872
rect 1854 14764 1860 14816
rect 1912 14804 1918 14816
rect 5460 14804 5488 14844
rect 6825 14841 6837 14844
rect 6871 14841 6883 14875
rect 7558 14872 7564 14884
rect 6825 14835 6883 14841
rect 7208 14844 7564 14872
rect 1912 14776 5488 14804
rect 1912 14764 1918 14776
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 5905 14807 5963 14813
rect 5905 14804 5917 14807
rect 5868 14776 5917 14804
rect 5868 14764 5874 14776
rect 5905 14773 5917 14776
rect 5951 14773 5963 14807
rect 5905 14767 5963 14773
rect 6086 14764 6092 14816
rect 6144 14804 6150 14816
rect 7208 14804 7236 14844
rect 7558 14832 7564 14844
rect 7616 14872 7622 14884
rect 7760 14872 7788 14903
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 8938 14900 8944 14952
rect 8996 14940 9002 14952
rect 9674 14940 9680 14952
rect 8996 14912 9680 14940
rect 8996 14900 9002 14912
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 9861 14943 9919 14949
rect 9861 14909 9873 14943
rect 9907 14909 9919 14943
rect 10244 14940 10272 14980
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 11974 14968 11980 15020
rect 12032 14968 12038 15020
rect 13096 15008 13124 15116
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 16850 15144 16856 15156
rect 14936 15116 16856 15144
rect 14182 15076 14188 15088
rect 12406 14980 13124 15008
rect 13188 15048 14188 15076
rect 10410 14940 10416 14952
rect 10244 14912 10416 14940
rect 9861 14903 9919 14909
rect 9876 14872 9904 14903
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10962 14900 10968 14952
rect 11020 14900 11026 14952
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14940 11759 14943
rect 12406 14940 12434 14980
rect 13188 14940 13216 15048
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 14734 15036 14740 15088
rect 14792 15076 14798 15088
rect 14936 15076 14964 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 22094 15144 22100 15156
rect 19306 15116 22100 15144
rect 16298 15076 16304 15088
rect 14792 15048 14964 15076
rect 16054 15048 16304 15076
rect 14792 15036 14798 15048
rect 16298 15036 16304 15048
rect 16356 15076 16362 15088
rect 16574 15076 16580 15088
rect 16356 15048 16580 15076
rect 16356 15036 16362 15048
rect 16574 15036 16580 15048
rect 16632 15036 16638 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 18322 15076 18328 15088
rect 16816 15048 18328 15076
rect 16816 15036 16822 15048
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 13814 15008 13820 15020
rect 13648 14980 13820 15008
rect 13648 14949 13676 14980
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 18414 14968 18420 15020
rect 18472 15008 18478 15020
rect 18874 15008 18880 15020
rect 18472 14980 18880 15008
rect 18472 14968 18478 14980
rect 18874 14968 18880 14980
rect 18932 15008 18938 15020
rect 19306 15008 19334 15116
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 23566 15104 23572 15156
rect 23624 15144 23630 15156
rect 23753 15147 23811 15153
rect 23753 15144 23765 15147
rect 23624 15116 23765 15144
rect 23624 15104 23630 15116
rect 23753 15113 23765 15116
rect 23799 15113 23811 15147
rect 23753 15107 23811 15113
rect 23842 15104 23848 15156
rect 23900 15144 23906 15156
rect 24029 15147 24087 15153
rect 24029 15144 24041 15147
rect 23900 15116 24041 15144
rect 23900 15104 23906 15116
rect 24029 15113 24041 15116
rect 24075 15144 24087 15147
rect 24213 15147 24271 15153
rect 24213 15144 24225 15147
rect 24075 15116 24225 15144
rect 24075 15113 24087 15116
rect 24029 15107 24087 15113
rect 24213 15113 24225 15116
rect 24259 15113 24271 15147
rect 24213 15107 24271 15113
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 27062 15104 27068 15156
rect 27120 15104 27126 15156
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 21542 15076 21548 15088
rect 20211 15048 21548 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 21542 15036 21548 15048
rect 21600 15036 21606 15088
rect 21818 15036 21824 15088
rect 21876 15076 21882 15088
rect 22281 15079 22339 15085
rect 22281 15076 22293 15079
rect 21876 15048 22293 15076
rect 21876 15036 21882 15048
rect 22281 15045 22293 15048
rect 22327 15045 22339 15079
rect 23860 15076 23888 15104
rect 23506 15048 23888 15076
rect 24964 15076 24992 15104
rect 25133 15079 25191 15085
rect 25133 15076 25145 15079
rect 24964 15048 25145 15076
rect 22281 15039 22339 15045
rect 25133 15045 25145 15048
rect 25179 15045 25191 15079
rect 27080 15076 27108 15104
rect 26358 15048 27108 15076
rect 25133 15039 25191 15045
rect 18932 14980 19334 15008
rect 18932 14968 18938 14980
rect 19702 14968 19708 15020
rect 19760 15008 19766 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19760 14980 20085 15008
rect 19760 14968 19766 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 15008 20867 15011
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 20855 14980 20913 15008
rect 20855 14977 20867 14980
rect 20809 14971 20867 14977
rect 20901 14977 20913 14980
rect 20947 15008 20959 15011
rect 20990 15008 20996 15020
rect 20947 14980 20996 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 22002 14968 22008 15020
rect 22060 14968 22066 15020
rect 23934 14968 23940 15020
rect 23992 15008 23998 15020
rect 24857 15011 24915 15017
rect 24857 15008 24869 15011
rect 23992 14980 24869 15008
rect 23992 14968 23998 14980
rect 24857 14977 24869 14980
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 11747 14912 12434 14940
rect 12544 14912 13216 14940
rect 13449 14943 13507 14949
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 10502 14872 10508 14884
rect 7616 14844 7696 14872
rect 7760 14844 8800 14872
rect 9876 14844 10508 14872
rect 7616 14832 7622 14844
rect 6144 14776 7236 14804
rect 6144 14764 6150 14776
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 7668 14804 7696 14844
rect 7834 14804 7840 14816
rect 7668 14776 7840 14804
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 8772 14804 8800 14844
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 10778 14832 10784 14884
rect 10836 14872 10842 14884
rect 12544 14872 12572 14912
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 13633 14903 13691 14909
rect 10836 14844 12572 14872
rect 13464 14872 13492 14903
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 14332 14912 14565 14940
rect 14332 14900 14338 14912
rect 14553 14909 14565 14912
rect 14599 14909 14611 14943
rect 14553 14903 14611 14909
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 14918 14940 14924 14952
rect 14875 14912 14924 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 16390 14900 16396 14952
rect 16448 14940 16454 14952
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16448 14912 16773 14940
rect 16448 14900 16454 14912
rect 16761 14909 16773 14912
rect 16807 14940 16819 14943
rect 20162 14940 20168 14952
rect 16807 14912 20168 14940
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 20349 14943 20407 14949
rect 20349 14909 20361 14943
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 14001 14875 14059 14881
rect 14001 14872 14013 14875
rect 13464 14844 14013 14872
rect 10836 14832 10842 14844
rect 14001 14841 14013 14844
rect 14047 14841 14059 14875
rect 14001 14835 14059 14841
rect 16224 14844 17172 14872
rect 9582 14804 9588 14816
rect 8772 14776 9588 14804
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 10413 14807 10471 14813
rect 10413 14804 10425 14807
rect 9732 14776 10425 14804
rect 9732 14764 9738 14776
rect 10413 14773 10425 14776
rect 10459 14773 10471 14807
rect 14016 14804 14044 14835
rect 16224 14804 16252 14844
rect 14016 14776 16252 14804
rect 10413 14767 10471 14773
rect 16298 14764 16304 14816
rect 16356 14764 16362 14816
rect 17144 14804 17172 14844
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 19978 14872 19984 14884
rect 17276 14844 19984 14872
rect 17276 14832 17282 14844
rect 19978 14832 19984 14844
rect 20036 14832 20042 14884
rect 20364 14872 20392 14903
rect 26142 14900 26148 14952
rect 26200 14940 26206 14952
rect 30558 14940 30564 14952
rect 26200 14912 30564 14940
rect 26200 14900 26206 14912
rect 30558 14900 30564 14912
rect 30616 14900 30622 14952
rect 21910 14872 21916 14884
rect 20364 14844 20668 14872
rect 18598 14804 18604 14816
rect 17144 14776 18604 14804
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 19150 14764 19156 14816
rect 19208 14764 19214 14816
rect 19334 14764 19340 14816
rect 19392 14764 19398 14816
rect 19705 14807 19763 14813
rect 19705 14773 19717 14807
rect 19751 14804 19763 14807
rect 20530 14804 20536 14816
rect 19751 14776 20536 14804
rect 19751 14773 19763 14776
rect 19705 14767 19763 14773
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 20640 14804 20668 14844
rect 20824 14844 21916 14872
rect 20824 14804 20852 14844
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 20640 14776 20852 14804
rect 26602 14764 26608 14816
rect 26660 14764 26666 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 5902 14600 5908 14612
rect 4019 14572 5908 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 6086 14560 6092 14612
rect 6144 14600 6150 14612
rect 6144 14572 9352 14600
rect 6144 14560 6150 14572
rect 5442 14532 5448 14544
rect 2746 14504 5448 14532
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 2746 14396 2774 14504
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 7193 14535 7251 14541
rect 7193 14501 7205 14535
rect 7239 14532 7251 14535
rect 7466 14532 7472 14544
rect 7239 14504 7472 14532
rect 7239 14501 7251 14504
rect 7193 14495 7251 14501
rect 7466 14492 7472 14504
rect 7524 14532 7530 14544
rect 7650 14532 7656 14544
rect 7524 14504 7656 14532
rect 7524 14492 7530 14504
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 9324 14532 9352 14572
rect 9398 14560 9404 14612
rect 9456 14560 9462 14612
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 9640 14572 11621 14600
rect 9640 14560 9646 14572
rect 11609 14569 11621 14572
rect 11655 14600 11667 14603
rect 13354 14600 13360 14612
rect 11655 14572 13360 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13725 14603 13783 14609
rect 13725 14600 13737 14603
rect 13596 14572 13737 14600
rect 13596 14560 13602 14572
rect 13725 14569 13737 14572
rect 13771 14600 13783 14603
rect 13814 14600 13820 14612
rect 13771 14572 13820 14600
rect 13771 14569 13783 14572
rect 13725 14563 13783 14569
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 14369 14603 14427 14609
rect 14369 14569 14381 14603
rect 14415 14600 14427 14603
rect 14734 14600 14740 14612
rect 14415 14572 14740 14600
rect 14415 14569 14427 14572
rect 14369 14563 14427 14569
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 14976 14572 18613 14600
rect 14976 14560 14982 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 18601 14563 18659 14569
rect 19429 14603 19487 14609
rect 19429 14569 19441 14603
rect 19475 14600 19487 14603
rect 26878 14600 26884 14612
rect 19475 14572 26884 14600
rect 19475 14569 19487 14572
rect 19429 14563 19487 14569
rect 26878 14560 26884 14572
rect 26936 14560 26942 14612
rect 26970 14560 26976 14612
rect 27028 14560 27034 14612
rect 10778 14532 10784 14544
rect 7984 14504 8340 14532
rect 9324 14504 10784 14532
rect 7984 14492 7990 14504
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 4893 14467 4951 14473
rect 4893 14464 4905 14467
rect 4488 14436 4905 14464
rect 4488 14424 4494 14436
rect 4893 14433 4905 14436
rect 4939 14464 4951 14467
rect 5810 14464 5816 14476
rect 4939 14436 5816 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 6730 14424 6736 14476
rect 6788 14464 6794 14476
rect 6788 14436 8248 14464
rect 6788 14424 6794 14436
rect 1811 14368 2774 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 4246 14356 4252 14408
rect 4304 14396 4310 14408
rect 4304 14368 4844 14396
rect 4304 14356 4310 14368
rect 2682 14288 2688 14340
rect 2740 14328 2746 14340
rect 4617 14331 4675 14337
rect 4617 14328 4629 14331
rect 2740 14300 4629 14328
rect 2740 14288 2746 14300
rect 4617 14297 4629 14300
rect 4663 14297 4675 14331
rect 4617 14291 4675 14297
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14260 3479 14263
rect 3510 14260 3516 14272
rect 3467 14232 3516 14260
rect 3467 14229 3479 14232
rect 3421 14223 3479 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 4249 14263 4307 14269
rect 4249 14229 4261 14263
rect 4295 14260 4307 14263
rect 4522 14260 4528 14272
rect 4295 14232 4528 14260
rect 4295 14229 4307 14232
rect 4249 14223 4307 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 4706 14220 4712 14272
rect 4764 14220 4770 14272
rect 4816 14260 4844 14368
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 8220 14405 8248 14436
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 5224 14368 5457 14396
rect 5224 14356 5230 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14365 8263 14399
rect 8312 14396 8340 14504
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 21358 14492 21364 14544
rect 21416 14532 21422 14544
rect 21545 14535 21603 14541
rect 21545 14532 21557 14535
rect 21416 14504 21557 14532
rect 21416 14492 21422 14504
rect 21545 14501 21557 14504
rect 21591 14501 21603 14535
rect 21545 14495 21603 14501
rect 21726 14492 21732 14544
rect 21784 14492 21790 14544
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 24029 14535 24087 14541
rect 24029 14532 24041 14535
rect 23716 14504 24041 14532
rect 23716 14492 23722 14504
rect 24029 14501 24041 14504
rect 24075 14532 24087 14535
rect 25774 14532 25780 14544
rect 24075 14504 25780 14532
rect 24075 14501 24087 14504
rect 24029 14495 24087 14501
rect 25774 14492 25780 14504
rect 25832 14492 25838 14544
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 9766 14464 9772 14476
rect 8527 14436 9772 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 9861 14467 9919 14473
rect 9861 14433 9873 14467
rect 9907 14464 9919 14467
rect 10045 14467 10103 14473
rect 9907 14436 9996 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 9968 14396 9996 14436
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10134 14464 10140 14476
rect 10091 14436 10140 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10744 14436 11161 14464
rect 10744 14424 10750 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 12253 14467 12311 14473
rect 12253 14433 12265 14467
rect 12299 14464 12311 14467
rect 12802 14464 12808 14476
rect 12299 14436 12808 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 15930 14464 15936 14476
rect 14967 14436 15936 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 15930 14424 15936 14436
rect 15988 14464 15994 14476
rect 16298 14464 16304 14476
rect 15988 14436 16304 14464
rect 15988 14424 15994 14436
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14464 16911 14467
rect 17126 14464 17132 14476
rect 16899 14436 17132 14464
rect 16899 14433 16911 14436
rect 16853 14427 16911 14433
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17586 14424 17592 14476
rect 17644 14464 17650 14476
rect 18877 14467 18935 14473
rect 18877 14464 18889 14467
rect 17644 14436 18889 14464
rect 17644 14424 17650 14436
rect 18877 14433 18889 14436
rect 18923 14464 18935 14467
rect 19150 14464 19156 14476
rect 18923 14436 19156 14464
rect 18923 14433 18935 14436
rect 18877 14427 18935 14433
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 19852 14436 21097 14464
rect 19852 14424 19858 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 10870 14396 10876 14408
rect 8312 14368 9904 14396
rect 9968 14368 10876 14396
rect 8205 14359 8263 14365
rect 5718 14288 5724 14340
rect 5776 14288 5782 14340
rect 6270 14288 6276 14340
rect 6328 14288 6334 14340
rect 7742 14288 7748 14340
rect 7800 14328 7806 14340
rect 8297 14331 8355 14337
rect 8297 14328 8309 14331
rect 7800 14300 8309 14328
rect 7800 14288 7806 14300
rect 8297 14297 8309 14300
rect 8343 14297 8355 14331
rect 8297 14291 8355 14297
rect 7374 14260 7380 14272
rect 4816 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 8938 14220 8944 14272
rect 8996 14260 9002 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8996 14232 9045 14260
rect 8996 14220 9002 14232
rect 9033 14229 9045 14232
rect 9079 14229 9091 14263
rect 9033 14223 9091 14229
rect 9766 14220 9772 14272
rect 9824 14220 9830 14272
rect 9876 14260 9904 14368
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11054 14396 11060 14408
rect 11011 14368 11060 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11974 14356 11980 14408
rect 12032 14356 12038 14408
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 14332 14368 14657 14396
rect 14332 14356 14338 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 16574 14396 16580 14408
rect 16054 14368 16580 14396
rect 14645 14359 14703 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 18432 14368 19625 14396
rect 17129 14331 17187 14337
rect 13478 14300 13952 14328
rect 13924 14272 13952 14300
rect 16316 14300 17080 14328
rect 10502 14260 10508 14272
rect 9876 14232 10508 14260
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 10836 14232 11069 14260
rect 10836 14220 10842 14232
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 11057 14223 11115 14229
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 13964 14232 14105 14260
rect 13964 14220 13970 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 15010 14220 15016 14272
rect 15068 14260 15074 14272
rect 16316 14260 16344 14300
rect 15068 14232 16344 14260
rect 15068 14220 15074 14232
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 17052 14260 17080 14300
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17402 14328 17408 14340
rect 17175 14300 17408 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 17586 14288 17592 14340
rect 17644 14288 17650 14340
rect 18432 14260 18460 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14396 21051 14399
rect 21744 14396 21772 14492
rect 22002 14424 22008 14476
rect 22060 14464 22066 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22060 14436 22293 14464
rect 22060 14424 22066 14436
rect 22281 14433 22293 14436
rect 22327 14464 22339 14467
rect 23934 14464 23940 14476
rect 22327 14436 23940 14464
rect 22327 14433 22339 14436
rect 22281 14427 22339 14433
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 25038 14424 25044 14476
rect 25096 14424 25102 14476
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14464 25191 14467
rect 26329 14467 26387 14473
rect 26329 14464 26341 14467
rect 25179 14436 26341 14464
rect 25179 14433 25191 14436
rect 25133 14427 25191 14433
rect 26329 14433 26341 14436
rect 26375 14464 26387 14467
rect 26602 14464 26608 14476
rect 26375 14436 26608 14464
rect 26375 14433 26387 14436
rect 26329 14427 26387 14433
rect 25148 14396 25176 14427
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 21039 14368 21772 14396
rect 23952 14368 25176 14396
rect 26145 14399 26203 14405
rect 21039 14365 21051 14368
rect 20993 14359 21051 14365
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 19484 14300 21864 14328
rect 19484 14288 19490 14300
rect 17052 14232 18460 14260
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 21358 14260 21364 14272
rect 20947 14232 21364 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 21836 14260 21864 14300
rect 21910 14288 21916 14340
rect 21968 14328 21974 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 21968 14300 22569 14328
rect 21968 14288 21974 14300
rect 22557 14297 22569 14300
rect 22603 14297 22615 14331
rect 23842 14328 23848 14340
rect 23782 14300 23848 14328
rect 22557 14291 22615 14297
rect 23842 14288 23848 14300
rect 23900 14288 23906 14340
rect 22646 14260 22652 14272
rect 21836 14232 22652 14260
rect 22646 14220 22652 14232
rect 22704 14220 22710 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23952 14260 23980 14368
rect 26145 14365 26157 14399
rect 26191 14396 26203 14399
rect 26970 14396 26976 14408
rect 26191 14368 26976 14396
rect 26191 14365 26203 14368
rect 26145 14359 26203 14365
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 24949 14331 25007 14337
rect 24949 14297 24961 14331
rect 24995 14328 25007 14331
rect 25130 14328 25136 14340
rect 24995 14300 25136 14328
rect 24995 14297 25007 14300
rect 24949 14291 25007 14297
rect 25130 14288 25136 14300
rect 25188 14328 25194 14340
rect 25866 14328 25872 14340
rect 25188 14300 25872 14328
rect 25188 14288 25194 14300
rect 25866 14288 25872 14300
rect 25924 14288 25930 14340
rect 26237 14331 26295 14337
rect 26237 14297 26249 14331
rect 26283 14328 26295 14331
rect 26326 14328 26332 14340
rect 26283 14300 26332 14328
rect 26283 14297 26295 14300
rect 26237 14291 26295 14297
rect 26326 14288 26332 14300
rect 26384 14328 26390 14340
rect 26789 14331 26847 14337
rect 26789 14328 26801 14331
rect 26384 14300 26801 14328
rect 26384 14288 26390 14300
rect 26789 14297 26801 14300
rect 26835 14297 26847 14331
rect 26789 14291 26847 14297
rect 22796 14232 23980 14260
rect 22796 14220 22802 14232
rect 24578 14220 24584 14272
rect 24636 14220 24642 14272
rect 25774 14220 25780 14272
rect 25832 14220 25838 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 4706 14056 4712 14068
rect 4111 14028 4712 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 6362 14056 6368 14068
rect 5675 14028 6368 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 4525 13991 4583 13997
rect 4525 13988 4537 13991
rect 2372 13960 4537 13988
rect 2372 13948 2378 13960
rect 4525 13957 4537 13960
rect 4571 13957 4583 13991
rect 4525 13951 4583 13957
rect 5718 13948 5724 14000
rect 5776 13948 5782 14000
rect 6932 13988 6960 14019
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 9582 14056 9588 14068
rect 8159 14028 9588 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 9692 14028 10916 14056
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 6932 13960 8493 13988
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 9692 13988 9720 14028
rect 8680 13960 9720 13988
rect 10888 13988 10916 14028
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11112 14028 11989 14056
rect 11112 14016 11118 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 12124 14028 13645 14056
rect 12124 14016 12130 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14240 14028 14749 14056
rect 14240 14016 14246 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 14826 14016 14832 14068
rect 14884 14016 14890 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16758 14056 16764 14068
rect 15611 14028 16764 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 17368 14028 18889 14056
rect 17368 14016 17374 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 20622 14056 20628 14068
rect 19475 14028 20628 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 21140 14028 23397 14056
rect 21140 14016 21146 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 24949 14059 25007 14065
rect 24949 14025 24961 14059
rect 24995 14056 25007 14059
rect 25774 14056 25780 14068
rect 24995 14028 25780 14056
rect 24995 14025 25007 14028
rect 24949 14019 25007 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 25866 14016 25872 14068
rect 25924 14016 25930 14068
rect 26878 14016 26884 14068
rect 26936 14056 26942 14068
rect 35066 14056 35072 14068
rect 26936 14028 35072 14056
rect 26936 14016 26942 14028
rect 35066 14016 35072 14028
rect 35124 14016 35130 14068
rect 13998 13988 14004 14000
rect 10888 13960 14004 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 1854 13920 1860 13932
rect 1811 13892 1860 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 3620 13852 3648 13883
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 4304 13892 4445 13920
rect 4304 13880 4310 13892
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 4540 13892 5212 13920
rect 4540 13852 4568 13892
rect 3620 13824 4568 13852
rect 4617 13855 4675 13861
rect 2041 13815 2099 13821
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 4798 13852 4804 13864
rect 4663 13824 4804 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 4632 13784 4660 13815
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5184 13852 5212 13892
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 5316 13892 7389 13920
rect 5316 13880 5322 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 8680 13920 8708 13960
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 16632 13960 16681 13988
rect 16632 13948 16638 13960
rect 16669 13957 16681 13960
rect 16715 13988 16727 13991
rect 16715 13960 17894 13988
rect 16715 13957 16727 13960
rect 16669 13951 16727 13957
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 21821 13991 21879 13997
rect 21821 13988 21833 13991
rect 21416 13960 21833 13988
rect 21416 13948 21422 13960
rect 21821 13957 21833 13960
rect 21867 13957 21879 13991
rect 23753 13991 23811 13997
rect 23753 13988 23765 13991
rect 21821 13951 21879 13957
rect 22756 13960 23765 13988
rect 10870 13920 10876 13932
rect 7377 13883 7435 13889
rect 7576 13892 8708 13920
rect 10718 13892 10876 13920
rect 5718 13852 5724 13864
rect 5184 13824 5724 13852
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 3476 13756 4660 13784
rect 5828 13784 5856 13815
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 6144 13824 6377 13852
rect 6144 13812 6150 13824
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 6365 13815 6423 13821
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 6696 13824 7420 13852
rect 6696 13812 6702 13824
rect 5902 13784 5908 13796
rect 5828 13756 5908 13784
rect 3476 13744 3482 13756
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 6454 13744 6460 13796
rect 6512 13784 6518 13796
rect 6549 13787 6607 13793
rect 6549 13784 6561 13787
rect 6512 13756 6561 13784
rect 6512 13744 6518 13756
rect 6549 13753 6561 13756
rect 6595 13753 6607 13787
rect 7392 13784 7420 13824
rect 7466 13812 7472 13864
rect 7524 13812 7530 13864
rect 7576 13784 7604 13892
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 11330 13880 11336 13932
rect 11388 13920 11394 13932
rect 11609 13923 11667 13929
rect 11609 13920 11621 13923
rect 11388 13892 11621 13920
rect 11388 13880 11394 13892
rect 11609 13889 11621 13892
rect 11655 13920 11667 13923
rect 12066 13920 12072 13932
rect 11655 13892 12072 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 12176 13892 12357 13920
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 7392 13756 7604 13784
rect 6549 13747 6607 13753
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 8680 13784 8708 13815
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 9631 13824 10916 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 7708 13756 8708 13784
rect 10888 13784 10916 13824
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 11020 13824 11069 13852
rect 11020 13812 11026 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 12176 13852 12204 13892
rect 12345 13889 12357 13892
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 13538 13880 13544 13932
rect 13596 13880 13602 13932
rect 15562 13920 15568 13932
rect 13740 13892 15568 13920
rect 11572 13824 12204 13852
rect 11572 13812 11578 13824
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12308 13824 12449 13852
rect 12308 13812 12314 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 13740 13852 13768 13892
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15804 13892 15945 13920
rect 15804 13880 15810 13892
rect 15933 13889 15945 13892
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16942 13920 16948 13932
rect 16071 13892 16948 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 12529 13815 12587 13821
rect 13188 13824 13768 13852
rect 11238 13784 11244 13796
rect 10888 13756 11244 13784
rect 7708 13744 7714 13756
rect 11238 13744 11244 13756
rect 11296 13784 11302 13796
rect 12544 13784 12572 13815
rect 13188 13793 13216 13824
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 14458 13852 14464 13864
rect 14384 13824 14464 13852
rect 11296 13756 12572 13784
rect 13173 13787 13231 13793
rect 11296 13744 11302 13756
rect 13173 13753 13185 13787
rect 13219 13753 13231 13787
rect 14182 13784 14188 13796
rect 13173 13747 13231 13753
rect 13280 13756 14188 13784
rect 5258 13676 5264 13728
rect 5316 13676 5322 13728
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 10042 13716 10048 13728
rect 8812 13688 10048 13716
rect 8812 13676 8818 13688
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 13280 13716 13308 13756
rect 14182 13744 14188 13756
rect 14240 13744 14246 13796
rect 14384 13793 14412 13824
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 14918 13812 14924 13864
rect 14976 13812 14982 13864
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15378 13852 15384 13864
rect 15252 13824 15384 13852
rect 15252 13812 15258 13824
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 16114 13812 16120 13864
rect 16172 13812 16178 13864
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 19628 13852 19656 13883
rect 20438 13880 20444 13932
rect 20496 13880 20502 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 21634 13920 21640 13932
rect 20579 13892 21640 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 21836 13920 21864 13951
rect 22756 13944 22784 13960
rect 23753 13957 23765 13960
rect 23799 13957 23811 13991
rect 23753 13951 23811 13957
rect 21836 13892 22324 13920
rect 17828 13824 19656 13852
rect 17828 13812 17834 13824
rect 19978 13812 19984 13864
rect 20036 13852 20042 13864
rect 20625 13855 20683 13861
rect 20036 13824 20116 13852
rect 20036 13812 20042 13824
rect 20088 13793 20116 13824
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 22296 13852 22324 13892
rect 22370 13880 22376 13932
rect 22428 13920 22434 13932
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22428 13892 22569 13920
rect 22428 13880 22434 13892
rect 22557 13889 22569 13892
rect 22603 13920 22615 13923
rect 22664 13920 22784 13944
rect 22603 13916 22784 13920
rect 23768 13920 23796 13951
rect 23842 13948 23848 14000
rect 23900 13948 23906 14000
rect 24578 13948 24584 14000
rect 24636 13988 24642 14000
rect 25041 13991 25099 13997
rect 25041 13988 25053 13991
rect 24636 13960 25053 13988
rect 24636 13948 24642 13960
rect 25041 13957 25053 13960
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 25130 13948 25136 14000
rect 25188 13988 25194 14000
rect 25593 13991 25651 13997
rect 25593 13988 25605 13991
rect 25188 13960 25605 13988
rect 25188 13948 25194 13960
rect 25593 13957 25605 13960
rect 25639 13957 25651 13991
rect 25593 13951 25651 13957
rect 25961 13923 26019 13929
rect 25961 13920 25973 13923
rect 22603 13892 22692 13916
rect 23768 13892 25973 13920
rect 22603 13889 22615 13892
rect 22557 13883 22615 13889
rect 25961 13889 25973 13892
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 22646 13852 22652 13864
rect 20625 13815 20683 13821
rect 20824 13824 22232 13852
rect 22296 13824 22652 13852
rect 14369 13787 14427 13793
rect 14369 13753 14381 13787
rect 14415 13753 14427 13787
rect 14369 13747 14427 13753
rect 20073 13787 20131 13793
rect 20073 13753 20085 13787
rect 20119 13753 20131 13787
rect 20640 13784 20668 13815
rect 20714 13784 20720 13796
rect 20640 13756 20720 13784
rect 20073 13747 20131 13753
rect 20714 13744 20720 13756
rect 20772 13744 20778 13796
rect 10192 13688 13308 13716
rect 10192 13676 10198 13688
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 14642 13716 14648 13728
rect 13412 13688 14648 13716
rect 13412 13676 13418 13688
rect 14642 13676 14648 13688
rect 14700 13676 14706 13728
rect 17392 13719 17450 13725
rect 17392 13685 17404 13719
rect 17438 13716 17450 13719
rect 17494 13716 17500 13728
rect 17438 13688 17500 13716
rect 17438 13685 17450 13688
rect 17392 13679 17450 13685
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20824 13716 20852 13824
rect 22204 13793 22232 13824
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 22830 13812 22836 13864
rect 22888 13852 22894 13864
rect 23750 13852 23756 13864
rect 22888 13824 23756 13852
rect 22888 13812 22894 13824
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 24026 13812 24032 13864
rect 24084 13812 24090 13864
rect 25130 13812 25136 13864
rect 25188 13852 25194 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 25188 13824 25237 13852
rect 25188 13812 25194 13824
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 26145 13855 26203 13861
rect 26145 13852 26157 13855
rect 25271 13824 26157 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 26145 13821 26157 13824
rect 26191 13821 26203 13855
rect 26145 13815 26203 13821
rect 22189 13787 22247 13793
rect 22189 13753 22201 13787
rect 22235 13753 22247 13787
rect 22189 13747 22247 13753
rect 20220 13688 20852 13716
rect 20220 13676 20226 13688
rect 20990 13676 20996 13728
rect 21048 13716 21054 13728
rect 22554 13716 22560 13728
rect 21048 13688 22560 13716
rect 21048 13676 21054 13688
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 24578 13676 24584 13728
rect 24636 13676 24642 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 4430 13521 4436 13524
rect 4420 13515 4436 13521
rect 4420 13481 4432 13515
rect 4420 13475 4436 13481
rect 4430 13472 4436 13475
rect 4488 13472 4494 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 10134 13512 10140 13524
rect 7156 13484 10140 13512
rect 7156 13472 7162 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 11204 13484 11437 13512
rect 11204 13472 11210 13484
rect 11425 13481 11437 13484
rect 11471 13481 11483 13515
rect 12434 13512 12440 13524
rect 11425 13475 11483 13481
rect 11532 13484 12440 13512
rect 5442 13404 5448 13456
rect 5500 13444 5506 13456
rect 5994 13444 6000 13456
rect 5500 13416 6000 13444
rect 5500 13404 5506 13416
rect 5994 13404 6000 13416
rect 6052 13404 6058 13456
rect 8570 13404 8576 13456
rect 8628 13444 8634 13456
rect 11532 13444 11560 13484
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 12860 13484 13737 13512
rect 12860 13472 12866 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 17402 13521 17408 13524
rect 17386 13515 17408 13521
rect 17386 13512 17398 13515
rect 13872 13484 17398 13512
rect 13872 13472 13878 13484
rect 17386 13481 17398 13484
rect 17386 13475 17408 13481
rect 17402 13472 17408 13475
rect 17460 13472 17466 13524
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 17552 13484 18889 13512
rect 17552 13472 17558 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 19518 13512 19524 13524
rect 19208 13484 19524 13512
rect 19208 13472 19214 13484
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 20990 13512 20996 13524
rect 20272 13484 20996 13512
rect 8628 13416 11560 13444
rect 8628 13404 8634 13416
rect 2038 13336 2044 13388
rect 2096 13336 2102 13388
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13376 4215 13379
rect 5166 13376 5172 13388
rect 4203 13348 5172 13376
rect 4203 13345 4215 13348
rect 4157 13339 4215 13345
rect 5166 13336 5172 13348
rect 5224 13376 5230 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 5224 13348 6745 13376
rect 5224 13336 5230 13348
rect 6733 13345 6745 13348
rect 6779 13376 6791 13379
rect 7374 13376 7380 13388
rect 6779 13348 7380 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 8496 13348 10977 13376
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 1946 13308 1952 13320
rect 1811 13280 1952 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 1946 13268 1952 13280
rect 2004 13268 2010 13320
rect 3878 13268 3884 13320
rect 3936 13268 3942 13320
rect 6270 13308 6276 13320
rect 5566 13294 6276 13308
rect 5552 13280 6276 13294
rect 1854 13200 1860 13252
rect 1912 13240 1918 13252
rect 3513 13243 3571 13249
rect 3513 13240 3525 13243
rect 1912 13212 3525 13240
rect 1912 13200 1918 13212
rect 3513 13209 3525 13212
rect 3559 13240 3571 13243
rect 4706 13240 4712 13252
rect 3559 13212 4712 13240
rect 3559 13209 3571 13212
rect 3513 13203 3571 13209
rect 4706 13200 4712 13212
rect 4764 13200 4770 13252
rect 2590 13132 2596 13184
rect 2648 13172 2654 13184
rect 3329 13175 3387 13181
rect 3329 13172 3341 13175
rect 2648 13144 3341 13172
rect 2648 13132 2654 13144
rect 3329 13141 3341 13144
rect 3375 13172 3387 13175
rect 3418 13172 3424 13184
rect 3375 13144 3424 13172
rect 3375 13141 3387 13144
rect 3329 13135 3387 13141
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 4798 13132 4804 13184
rect 4856 13172 4862 13184
rect 5552 13172 5580 13280
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 5810 13200 5816 13252
rect 5868 13240 5874 13252
rect 5994 13240 6000 13252
rect 5868 13212 6000 13240
rect 5868 13200 5874 13212
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 6288 13240 6316 13268
rect 7009 13243 7067 13249
rect 6288 13212 6960 13240
rect 4856 13144 5580 13172
rect 4856 13132 4862 13144
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 6273 13175 6331 13181
rect 6273 13141 6285 13175
rect 6319 13172 6331 13175
rect 6362 13172 6368 13184
rect 6319 13144 6368 13172
rect 6319 13141 6331 13144
rect 6273 13135 6331 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 6546 13172 6552 13184
rect 6503 13144 6552 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 6932 13172 6960 13212
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 7282 13240 7288 13252
rect 7055 13212 7288 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 7466 13240 7472 13252
rect 7392 13212 7472 13240
rect 7392 13172 7420 13212
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 6932 13144 7420 13172
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8496 13181 8524 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11514 13376 11520 13388
rect 11296 13348 11520 13376
rect 11296 13336 11302 13348
rect 11514 13336 11520 13348
rect 11572 13376 11578 13388
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 11572 13348 11621 13376
rect 11572 13336 11578 13348
rect 11609 13345 11621 13348
rect 11655 13345 11667 13379
rect 11609 13339 11667 13345
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 13262 13376 13268 13388
rect 12032 13348 13268 13376
rect 12032 13336 12038 13348
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15194 13376 15200 13388
rect 14599 13348 15200 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15194 13336 15200 13348
rect 15252 13376 15258 13388
rect 16390 13376 16396 13388
rect 15252 13348 16396 13376
rect 15252 13336 15258 13348
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17494 13376 17500 13388
rect 17184 13348 17500 13376
rect 17184 13336 17190 13348
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 20272 13376 20300 13484
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21818 13472 21824 13524
rect 21876 13512 21882 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 21876 13484 22109 13512
rect 21876 13472 21882 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 22370 13472 22376 13524
rect 22428 13512 22434 13524
rect 22465 13515 22523 13521
rect 22465 13512 22477 13515
rect 22428 13484 22477 13512
rect 22428 13472 22434 13484
rect 22465 13481 22477 13484
rect 22511 13481 22523 13515
rect 22465 13475 22523 13481
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23937 13515 23995 13521
rect 23937 13512 23949 13515
rect 23348 13484 23949 13512
rect 23348 13472 23354 13484
rect 23937 13481 23949 13484
rect 23983 13481 23995 13515
rect 23937 13475 23995 13481
rect 21634 13404 21640 13456
rect 21692 13444 21698 13456
rect 22833 13447 22891 13453
rect 22833 13444 22845 13447
rect 21692 13416 22845 13444
rect 21692 13404 21698 13416
rect 22833 13413 22845 13416
rect 22879 13413 22891 13447
rect 23382 13444 23388 13456
rect 22833 13407 22891 13413
rect 23308 13416 23388 13444
rect 17920 13348 20300 13376
rect 20349 13379 20407 13385
rect 17920 13336 17926 13348
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 22186 13376 22192 13388
rect 20395 13348 22192 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 23308 13385 23336 13416
rect 23382 13404 23388 13416
rect 23440 13404 23446 13456
rect 23842 13404 23848 13456
rect 23900 13444 23906 13456
rect 24121 13447 24179 13453
rect 24121 13444 24133 13447
rect 23900 13416 24133 13444
rect 23900 13404 23906 13416
rect 24121 13413 24133 13416
rect 24167 13413 24179 13447
rect 24121 13407 24179 13413
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13345 23351 13379
rect 23293 13339 23351 13345
rect 23474 13336 23480 13388
rect 23532 13336 23538 13388
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 32490 13376 32496 13388
rect 23624 13348 32496 13376
rect 23624 13336 23630 13348
rect 32490 13336 32496 13348
rect 32548 13336 32554 13388
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9140 13240 9168 13271
rect 9398 13268 9404 13320
rect 9456 13268 9462 13320
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13308 10839 13311
rect 11698 13308 11704 13320
rect 10827 13280 11704 13308
rect 10827 13277 10839 13280
rect 10781 13271 10839 13277
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 19150 13308 19156 13320
rect 18538 13280 19156 13308
rect 19150 13268 19156 13280
rect 19208 13268 19214 13320
rect 19337 13311 19395 13317
rect 19337 13277 19349 13311
rect 19383 13308 19395 13311
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 19383 13280 19441 13308
rect 19383 13277 19395 13280
rect 19337 13271 19395 13277
rect 19429 13277 19441 13280
rect 19475 13308 19487 13311
rect 19518 13308 19524 13320
rect 19475 13280 19524 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 19518 13268 19524 13280
rect 19576 13268 19582 13320
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23072 13280 25452 13308
rect 23072 13268 23078 13280
rect 12253 13243 12311 13249
rect 9140 13212 11744 13240
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 7708 13144 8493 13172
rect 7708 13132 7714 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 10410 13132 10416 13184
rect 10468 13132 10474 13184
rect 10870 13132 10876 13184
rect 10928 13132 10934 13184
rect 11716 13172 11744 13212
rect 12253 13209 12265 13243
rect 12299 13240 12311 13243
rect 12342 13240 12348 13252
rect 12299 13212 12348 13240
rect 12299 13209 12311 13212
rect 12253 13203 12311 13209
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 13906 13240 13912 13252
rect 13478 13212 13912 13240
rect 13906 13200 13912 13212
rect 13964 13200 13970 13252
rect 15838 13240 15844 13252
rect 15778 13212 15844 13240
rect 15838 13200 15844 13212
rect 15896 13240 15902 13252
rect 16574 13240 16580 13252
rect 15896 13212 16580 13240
rect 15896 13200 15902 13212
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 18966 13240 18972 13252
rect 18708 13212 18972 13240
rect 13630 13172 13636 13184
rect 11716 13144 13636 13172
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14366 13172 14372 13184
rect 14056 13144 14372 13172
rect 14056 13132 14062 13144
rect 14366 13132 14372 13144
rect 14424 13172 14430 13184
rect 16025 13175 16083 13181
rect 16025 13172 16037 13175
rect 14424 13144 16037 13172
rect 14424 13132 14430 13144
rect 16025 13141 16037 13144
rect 16071 13141 16083 13175
rect 16025 13135 16083 13141
rect 16114 13132 16120 13184
rect 16172 13172 16178 13184
rect 18708 13172 18736 13212
rect 18966 13200 18972 13212
rect 19024 13240 19030 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 19024 13212 20637 13240
rect 19024 13200 19030 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 20625 13203 20683 13209
rect 21174 13200 21180 13252
rect 21232 13200 21238 13252
rect 23201 13243 23259 13249
rect 23201 13209 23213 13243
rect 23247 13240 23259 13243
rect 23247 13212 23336 13240
rect 23247 13209 23259 13212
rect 23201 13203 23259 13209
rect 16172 13144 18736 13172
rect 16172 13132 16178 13144
rect 20346 13132 20352 13184
rect 20404 13172 20410 13184
rect 23106 13172 23112 13184
rect 20404 13144 23112 13172
rect 20404 13132 20410 13144
rect 23106 13132 23112 13144
rect 23164 13132 23170 13184
rect 23308 13172 23336 13212
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 25424 13249 25452 13280
rect 24581 13243 24639 13249
rect 24581 13240 24593 13243
rect 23440 13212 24593 13240
rect 23440 13200 23446 13212
rect 24581 13209 24593 13212
rect 24627 13209 24639 13243
rect 24581 13203 24639 13209
rect 25409 13243 25467 13249
rect 25409 13209 25421 13243
rect 25455 13240 25467 13243
rect 26878 13240 26884 13252
rect 25455 13212 26884 13240
rect 25455 13209 25467 13212
rect 25409 13203 25467 13209
rect 26878 13200 26884 13212
rect 26936 13200 26942 13252
rect 25222 13172 25228 13184
rect 23308 13144 25228 13172
rect 25222 13132 25228 13144
rect 25280 13132 25286 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 3602 12928 3608 12980
rect 3660 12928 3666 12980
rect 5534 12968 5540 12980
rect 4172 12940 5540 12968
rect 3513 12903 3571 12909
rect 3513 12869 3525 12903
rect 3559 12900 3571 12903
rect 4172 12900 4200 12940
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 6638 12968 6644 12980
rect 5776 12940 6644 12968
rect 5776 12928 5782 12940
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 10594 12968 10600 12980
rect 7331 12940 10600 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12529 12971 12587 12977
rect 12529 12968 12541 12971
rect 11848 12940 12541 12968
rect 11848 12928 11854 12940
rect 12529 12937 12541 12940
rect 12575 12937 12587 12971
rect 12529 12931 12587 12937
rect 13446 12928 13452 12980
rect 13504 12968 13510 12980
rect 13630 12968 13636 12980
rect 13504 12940 13636 12968
rect 13504 12928 13510 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 13722 12928 13728 12980
rect 13780 12928 13786 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 14458 12968 14464 12980
rect 14231 12940 14464 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14458 12928 14464 12940
rect 14516 12968 14522 12980
rect 15286 12968 15292 12980
rect 14516 12940 15292 12968
rect 14516 12928 14522 12940
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 16574 12968 16580 12980
rect 16255 12940 16580 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17000 12940 17785 12968
rect 17000 12928 17006 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 20162 12968 20168 12980
rect 18187 12940 20168 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 22189 12971 22247 12977
rect 22189 12968 22201 12971
rect 21232 12940 22201 12968
rect 21232 12928 21238 12940
rect 22189 12937 22201 12940
rect 22235 12937 22247 12971
rect 22189 12931 22247 12937
rect 23106 12928 23112 12980
rect 23164 12968 23170 12980
rect 23474 12968 23480 12980
rect 23164 12940 23480 12968
rect 23164 12928 23170 12940
rect 23474 12928 23480 12940
rect 23532 12968 23538 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23532 12940 24777 12968
rect 23532 12928 23538 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 3559 12872 4200 12900
rect 4249 12903 4307 12909
rect 3559 12869 3571 12872
rect 3513 12863 3571 12869
rect 3620 12844 3648 12872
rect 4249 12869 4261 12903
rect 4295 12900 4307 12903
rect 4338 12900 4344 12912
rect 4295 12872 4344 12900
rect 4295 12869 4307 12872
rect 4249 12863 4307 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 4433 12903 4491 12909
rect 4433 12869 4445 12903
rect 4479 12900 4491 12903
rect 4614 12900 4620 12912
rect 4479 12872 4620 12900
rect 4479 12869 4491 12872
rect 4433 12863 4491 12869
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 4706 12860 4712 12912
rect 4764 12900 4770 12912
rect 4801 12903 4859 12909
rect 4801 12900 4813 12903
rect 4764 12872 4813 12900
rect 4764 12860 4770 12872
rect 4801 12869 4813 12872
rect 4847 12900 4859 12903
rect 5442 12900 5448 12912
rect 4847 12872 5448 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 5629 12903 5687 12909
rect 5629 12869 5641 12903
rect 5675 12900 5687 12903
rect 5810 12900 5816 12912
rect 5675 12872 5816 12900
rect 5675 12869 5687 12872
rect 5629 12863 5687 12869
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 6457 12903 6515 12909
rect 6457 12900 6469 12903
rect 6328 12872 6469 12900
rect 6328 12860 6334 12872
rect 6457 12869 6469 12872
rect 6503 12869 6515 12903
rect 6457 12863 6515 12869
rect 7193 12903 7251 12909
rect 7193 12869 7205 12903
rect 7239 12900 7251 12903
rect 8570 12900 8576 12912
rect 7239 12872 8576 12900
rect 7239 12869 7251 12872
rect 7193 12863 7251 12869
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 2498 12832 2504 12844
rect 1903 12804 2504 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3602 12792 3608 12844
rect 3660 12792 3666 12844
rect 4062 12792 4068 12844
rect 4120 12792 4126 12844
rect 6822 12832 6828 12844
rect 4264 12804 6828 12832
rect 1210 12724 1216 12776
rect 1268 12764 1274 12776
rect 1581 12767 1639 12773
rect 1581 12764 1593 12767
rect 1268 12736 1593 12764
rect 1268 12724 1274 12736
rect 1581 12733 1593 12736
rect 1627 12733 1639 12767
rect 1581 12727 1639 12733
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 3326 12764 3332 12776
rect 2823 12736 3332 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 3326 12724 3332 12736
rect 3384 12764 3390 12776
rect 4080 12764 4108 12792
rect 4264 12776 4292 12804
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 3384 12736 4108 12764
rect 3384 12724 3390 12736
rect 4246 12724 4252 12776
rect 4304 12724 4310 12776
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4856 12736 4905 12764
rect 4856 12724 4862 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 5994 12764 6000 12776
rect 5951 12736 6000 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 5994 12724 6000 12736
rect 6052 12764 6058 12776
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 6052 12736 7389 12764
rect 6052 12724 6058 12736
rect 7377 12733 7389 12736
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 2038 12656 2044 12708
rect 2096 12696 2102 12708
rect 3145 12699 3203 12705
rect 3145 12696 3157 12699
rect 2096 12668 3157 12696
rect 2096 12656 2102 12668
rect 3145 12665 3157 12668
rect 3191 12696 3203 12699
rect 7484 12696 7512 12872
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 8754 12860 8760 12912
rect 8812 12860 8818 12912
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 13170 12900 13176 12912
rect 11931 12872 13176 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 13354 12860 13360 12912
rect 13412 12900 13418 12912
rect 14274 12900 14280 12912
rect 13412 12872 14280 12900
rect 13412 12860 13418 12872
rect 14274 12860 14280 12872
rect 14332 12900 14338 12912
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 14332 12872 15669 12900
rect 14332 12860 14338 12872
rect 15657 12869 15669 12872
rect 15703 12869 15715 12903
rect 18874 12900 18880 12912
rect 15657 12863 15715 12869
rect 16316 12872 18880 12900
rect 10686 12792 10692 12844
rect 10744 12792 10750 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12406 12804 12909 12832
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 9030 12764 9036 12776
rect 8343 12736 9036 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 3191 12668 7512 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 2961 12631 3019 12637
rect 2961 12597 2973 12631
rect 3007 12628 3019 12631
rect 3510 12628 3516 12640
rect 3007 12600 3516 12628
rect 3007 12597 3019 12600
rect 2961 12591 3019 12597
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5626 12628 5632 12640
rect 5307 12600 5632 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 6822 12588 6828 12640
rect 6880 12588 6886 12640
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 8036 12628 8064 12727
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 10008 12736 10057 12764
rect 10008 12724 10014 12736
rect 10045 12733 10057 12736
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 12406 12764 12434 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 13446 12792 13452 12844
rect 13504 12832 13510 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13504 12804 14105 12832
rect 13504 12792 13510 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14826 12832 14832 12844
rect 14093 12795 14151 12801
rect 14292 12804 14832 12832
rect 10192 12736 12434 12764
rect 12989 12767 13047 12773
rect 10192 12724 10198 12736
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 10502 12656 10508 12708
rect 10560 12656 10566 12708
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 11333 12699 11391 12705
rect 11333 12696 11345 12699
rect 10836 12668 11345 12696
rect 10836 12656 10842 12668
rect 11333 12665 11345 12668
rect 11379 12696 11391 12699
rect 12618 12696 12624 12708
rect 11379 12668 12624 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 13004 12696 13032 12727
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14292 12764 14320 12804
rect 14826 12792 14832 12804
rect 14884 12832 14890 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14884 12804 14933 12832
rect 14884 12792 14890 12804
rect 14921 12801 14933 12804
rect 14967 12832 14979 12835
rect 15102 12832 15108 12844
rect 14967 12804 15108 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 15102 12792 15108 12804
rect 15160 12832 15166 12844
rect 16316 12841 16344 12872
rect 18874 12860 18880 12872
rect 18932 12900 18938 12912
rect 18969 12903 19027 12909
rect 18969 12900 18981 12903
rect 18932 12872 18981 12900
rect 18932 12860 18938 12872
rect 18969 12869 18981 12872
rect 19015 12869 19027 12903
rect 18969 12863 19027 12869
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 23566 12900 23572 12912
rect 20680 12872 23572 12900
rect 20680 12860 20686 12872
rect 23566 12860 23572 12872
rect 23624 12860 23630 12912
rect 23934 12860 23940 12912
rect 23992 12860 23998 12912
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 15160 12804 16313 12832
rect 15160 12792 15166 12804
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 17954 12832 17960 12844
rect 17460 12804 17960 12832
rect 17460 12792 17466 12804
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 21177 12835 21235 12841
rect 18279 12804 20208 12832
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 13872 12736 14320 12764
rect 14369 12767 14427 12773
rect 13872 12724 13878 12736
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 15194 12764 15200 12776
rect 14415 12736 15200 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 16850 12724 16856 12776
rect 16908 12724 16914 12776
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12764 18475 12767
rect 18598 12764 18604 12776
rect 18463 12736 18604 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20070 12764 20076 12776
rect 19843 12736 20076 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 17218 12696 17224 12708
rect 13004 12668 17224 12696
rect 17218 12656 17224 12668
rect 17276 12656 17282 12708
rect 17494 12656 17500 12708
rect 17552 12696 17558 12708
rect 19812 12696 19840 12727
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 17552 12668 19840 12696
rect 20180 12696 20208 12804
rect 21177 12801 21189 12835
rect 21223 12832 21235 12835
rect 22094 12832 22100 12844
rect 21223 12804 22100 12832
rect 21223 12801 21235 12804
rect 21177 12795 21235 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 23014 12832 23020 12844
rect 22244 12804 23020 12832
rect 22244 12792 22250 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 23658 12764 23664 12776
rect 23339 12736 23664 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 23934 12724 23940 12776
rect 23992 12764 23998 12776
rect 24486 12764 24492 12776
rect 23992 12736 24492 12764
rect 23992 12724 23998 12736
rect 24486 12724 24492 12736
rect 24544 12764 24550 12776
rect 25041 12767 25099 12773
rect 25041 12764 25053 12767
rect 24544 12736 25053 12764
rect 24544 12724 24550 12736
rect 25041 12733 25053 12736
rect 25087 12733 25099 12767
rect 25041 12727 25099 12733
rect 22462 12696 22468 12708
rect 20180 12668 22468 12696
rect 17552 12656 17558 12668
rect 22462 12656 22468 12668
rect 22520 12656 22526 12708
rect 9306 12628 9312 12640
rect 7432 12600 9312 12628
rect 7432 12588 7438 12600
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 10318 12628 10324 12640
rect 10100 12600 10324 12628
rect 10100 12588 10106 12600
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 11146 12588 11152 12640
rect 11204 12588 11210 12640
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 11480 12600 11621 12628
rect 11480 12588 11486 12600
rect 11609 12597 11621 12600
rect 11655 12628 11667 12631
rect 12250 12628 12256 12640
rect 11655 12600 12256 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 12250 12588 12256 12600
rect 12308 12628 12314 12640
rect 13446 12628 13452 12640
rect 12308 12600 13452 12628
rect 12308 12588 12314 12600
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 14182 12628 14188 12640
rect 14056 12600 14188 12628
rect 14056 12588 14062 12600
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 16850 12628 16856 12640
rect 14700 12600 16856 12628
rect 14700 12588 14706 12600
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 19484 12600 20729 12628
rect 19484 12588 19490 12600
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4338 12424 4344 12436
rect 4019 12396 4344 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 7190 12424 7196 12436
rect 4663 12396 7196 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 3510 12316 3516 12368
rect 3568 12356 3574 12368
rect 3605 12359 3663 12365
rect 3605 12356 3617 12359
rect 3568 12328 3617 12356
rect 3568 12316 3574 12328
rect 3605 12325 3617 12328
rect 3651 12356 3663 12359
rect 3651 12328 4660 12356
rect 3651 12325 3663 12328
rect 3605 12319 3663 12325
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 4246 12288 4252 12300
rect 1903 12260 4252 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1486 12220 1492 12232
rect 992 12192 1492 12220
rect 992 12180 998 12192
rect 1486 12180 1492 12192
rect 1544 12220 1550 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1544 12192 1593 12220
rect 1544 12180 1550 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 4154 12180 4160 12232
rect 4212 12180 4218 12232
rect 4632 12220 4660 12328
rect 4724 12297 4752 12396
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 10870 12424 10876 12436
rect 7883 12396 10876 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11793 12427 11851 12433
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 12526 12424 12532 12436
rect 11839 12396 12532 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 13906 12424 13912 12436
rect 12676 12396 13912 12424
rect 12676 12384 12682 12396
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 14458 12384 14464 12436
rect 14516 12384 14522 12436
rect 15194 12424 15200 12436
rect 14568 12396 15200 12424
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 7340 12328 7696 12356
rect 7340 12316 7346 12328
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 5224 12260 5365 12288
rect 5224 12248 5230 12260
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 7558 12288 7564 12300
rect 7423 12260 7564 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 7668 12288 7696 12328
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 9398 12356 9404 12368
rect 8996 12328 9404 12356
rect 8996 12316 9002 12328
rect 9398 12316 9404 12328
rect 9456 12316 9462 12368
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 12989 12359 13047 12365
rect 11388 12328 12848 12356
rect 11388 12316 11394 12328
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 7668 12260 8401 12288
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9364 12260 9873 12288
rect 9364 12248 9370 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 12066 12288 12072 12300
rect 11287 12260 12072 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 4798 12220 4804 12232
rect 4632 12192 4804 12220
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 9674 12220 9680 12232
rect 8343 12192 9680 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12220 11115 12223
rect 12618 12220 12624 12232
rect 11103 12192 12624 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2832 12124 2973 12152
rect 2832 12112 2838 12124
rect 2961 12121 2973 12124
rect 3007 12121 3019 12155
rect 2961 12115 3019 12121
rect 3145 12155 3203 12161
rect 3145 12121 3157 12155
rect 3191 12152 3203 12155
rect 5074 12152 5080 12164
rect 3191 12124 5080 12152
rect 3191 12121 3203 12124
rect 3145 12115 3203 12121
rect 5074 12112 5080 12124
rect 5132 12112 5138 12164
rect 5629 12155 5687 12161
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 5718 12152 5724 12164
rect 5675 12124 5724 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 6270 12112 6276 12164
rect 6328 12112 6334 12164
rect 9122 12112 9128 12164
rect 9180 12112 9186 12164
rect 9766 12112 9772 12164
rect 9824 12152 9830 12164
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 9824 12124 10977 12152
rect 9824 12112 9830 12124
rect 10965 12121 10977 12124
rect 11011 12121 11023 12155
rect 10965 12115 11023 12121
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 12253 12155 12311 12161
rect 12253 12152 12265 12155
rect 11204 12124 12265 12152
rect 11204 12112 11210 12124
rect 12253 12121 12265 12124
rect 12299 12152 12311 12155
rect 12820 12152 12848 12328
rect 12989 12325 13001 12359
rect 13035 12356 13047 12359
rect 13262 12356 13268 12368
rect 13035 12328 13268 12356
rect 13035 12325 13047 12328
rect 12989 12319 13047 12325
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 14568 12356 14596 12396
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18049 12427 18107 12433
rect 18049 12424 18061 12427
rect 18012 12396 18061 12424
rect 18012 12384 18018 12396
rect 18049 12393 18061 12396
rect 18095 12393 18107 12427
rect 18049 12387 18107 12393
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 18417 12427 18475 12433
rect 18417 12424 18429 12427
rect 18196 12396 18429 12424
rect 18196 12384 18202 12396
rect 18417 12393 18429 12396
rect 18463 12424 18475 12427
rect 18969 12427 19027 12433
rect 18969 12424 18981 12427
rect 18463 12396 18981 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 18969 12393 18981 12396
rect 19015 12424 19027 12427
rect 19150 12424 19156 12436
rect 19015 12396 19156 12424
rect 19015 12393 19027 12396
rect 18969 12387 19027 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21821 12427 21879 12433
rect 21821 12424 21833 12427
rect 20772 12396 21833 12424
rect 20772 12384 20778 12396
rect 21821 12393 21833 12396
rect 21867 12424 21879 12427
rect 21867 12396 22094 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 13648 12328 14596 12356
rect 13648 12297 13676 12328
rect 18874 12316 18880 12368
rect 18932 12316 18938 12368
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 14642 12248 14648 12300
rect 14700 12248 14706 12300
rect 14826 12248 14832 12300
rect 14884 12288 14890 12300
rect 15933 12291 15991 12297
rect 15933 12288 15945 12291
rect 14884 12260 15945 12288
rect 14884 12248 14890 12260
rect 15933 12257 15945 12260
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 16574 12248 16580 12300
rect 16632 12248 16638 12300
rect 17310 12248 17316 12300
rect 17368 12288 17374 12300
rect 19521 12291 19579 12297
rect 19521 12288 19533 12291
rect 17368 12260 19533 12288
rect 17368 12248 17374 12260
rect 19521 12257 19533 12260
rect 19567 12288 19579 12291
rect 19567 12260 19840 12288
rect 19567 12257 19579 12260
rect 19521 12251 19579 12257
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 14660 12220 14688 12248
rect 13403 12192 14688 12220
rect 14737 12223 14795 12229
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14844 12220 14872 12248
rect 14783 12192 14872 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 14976 12192 15577 12220
rect 14976 12180 14982 12192
rect 15565 12189 15577 12192
rect 15611 12220 15623 12223
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 15611 12192 16313 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 18138 12220 18144 12232
rect 17710 12192 18144 12220
rect 16301 12183 16359 12189
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 13449 12155 13507 12161
rect 13449 12152 13461 12155
rect 12299 12124 12434 12152
rect 12820 12124 13461 12152
rect 12299 12121 12311 12124
rect 12253 12115 12311 12121
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 4338 12084 4344 12096
rect 3844 12056 4344 12084
rect 3844 12044 3850 12056
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7616 12056 8217 12084
rect 7616 12044 7622 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 11940 12056 12173 12084
rect 11940 12044 11946 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 12406 12084 12434 12124
rect 13449 12121 13461 12124
rect 13495 12121 13507 12155
rect 19702 12152 19708 12164
rect 13449 12115 13507 12121
rect 17880 12124 19708 12152
rect 13170 12084 13176 12096
rect 12406 12056 13176 12084
rect 12161 12047 12219 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13906 12044 13912 12096
rect 13964 12084 13970 12096
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 13964 12056 14105 12084
rect 13964 12044 13970 12056
rect 14093 12053 14105 12056
rect 14139 12084 14151 12087
rect 14826 12084 14832 12096
rect 14139 12056 14832 12084
rect 14139 12053 14151 12056
rect 14093 12047 14151 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 16206 12044 16212 12096
rect 16264 12084 16270 12096
rect 17880 12084 17908 12124
rect 19702 12112 19708 12124
rect 19760 12112 19766 12164
rect 16264 12056 17908 12084
rect 16264 12044 16270 12056
rect 18414 12044 18420 12096
rect 18472 12084 18478 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 18472 12056 18521 12084
rect 18472 12044 18478 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 18932 12056 19349 12084
rect 18932 12044 18938 12056
rect 19337 12053 19349 12056
rect 19383 12053 19395 12087
rect 19812 12084 19840 12260
rect 20070 12248 20076 12300
rect 20128 12248 20134 12300
rect 22066 12288 22094 12396
rect 24486 12384 24492 12436
rect 24544 12384 24550 12436
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 22066 12260 22569 12288
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22244 12192 22293 12220
rect 22244 12180 22250 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 23934 12220 23940 12232
rect 23690 12192 23940 12220
rect 22281 12183 22339 12189
rect 23934 12180 23940 12192
rect 23992 12180 23998 12232
rect 20346 12112 20352 12164
rect 20404 12112 20410 12164
rect 21082 12112 21088 12164
rect 21140 12112 21146 12164
rect 25038 12152 25044 12164
rect 23860 12124 25044 12152
rect 23860 12084 23888 12124
rect 25038 12112 25044 12124
rect 25096 12112 25102 12164
rect 19812 12056 23888 12084
rect 19337 12047 19395 12053
rect 24026 12044 24032 12096
rect 24084 12044 24090 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 1762 11840 1768 11892
rect 1820 11840 1826 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3510 11880 3516 11892
rect 3467 11852 3516 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4479 11852 5273 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 5626 11840 5632 11892
rect 5684 11840 5690 11892
rect 6454 11840 6460 11892
rect 6512 11840 6518 11892
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 12345 11883 12403 11889
rect 12345 11880 12357 11883
rect 6779 11852 12357 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 12345 11849 12357 11852
rect 12391 11849 12403 11883
rect 14090 11880 14096 11892
rect 12345 11843 12403 11849
rect 13096 11852 14096 11880
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 4154 11812 4160 11824
rect 1719 11784 4160 11812
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 5721 11815 5779 11821
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 6822 11812 6828 11824
rect 5767 11784 6828 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7650 11772 7656 11824
rect 7708 11772 7714 11824
rect 8110 11772 8116 11824
rect 8168 11772 8174 11824
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 9490 11812 9496 11824
rect 9364 11784 9496 11812
rect 9364 11772 9370 11784
rect 9490 11772 9496 11784
rect 9548 11812 9554 11824
rect 9950 11812 9956 11824
rect 9548 11784 9956 11812
rect 9548 11772 9554 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10594 11772 10600 11824
rect 10652 11812 10658 11824
rect 12437 11815 12495 11821
rect 12437 11812 12449 11815
rect 10652 11784 12449 11812
rect 10652 11772 10658 11784
rect 12437 11781 12449 11784
rect 12483 11781 12495 11815
rect 12437 11775 12495 11781
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1946 11744 1952 11756
rect 1535 11716 1952 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2406 11704 2412 11756
rect 2464 11704 2470 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 5258 11744 5264 11756
rect 4571 11716 5264 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9180 11716 9597 11744
rect 9180 11704 9186 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11609 11747 11667 11753
rect 11609 11744 11621 11747
rect 11388 11716 11621 11744
rect 11388 11704 11394 11716
rect 11609 11713 11621 11716
rect 11655 11713 11667 11747
rect 13096 11744 13124 11852
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 14424 11852 17325 11880
rect 14424 11840 14430 11852
rect 17313 11849 17325 11852
rect 17359 11880 17371 11883
rect 18509 11883 18567 11889
rect 17359 11852 18092 11880
rect 17359 11849 17371 11852
rect 17313 11843 17371 11849
rect 13354 11812 13360 11824
rect 13188 11784 13360 11812
rect 13188 11753 13216 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 14826 11812 14832 11824
rect 14674 11784 14832 11812
rect 14826 11772 14832 11784
rect 14884 11812 14890 11824
rect 15289 11815 15347 11821
rect 15289 11812 15301 11815
rect 14884 11784 15301 11812
rect 14884 11772 14890 11784
rect 15289 11781 15301 11784
rect 15335 11812 15347 11815
rect 15838 11812 15844 11824
rect 15335 11784 15844 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 16025 11815 16083 11821
rect 16025 11781 16037 11815
rect 16071 11812 16083 11815
rect 18064 11812 18092 11852
rect 18509 11849 18521 11883
rect 18555 11880 18567 11883
rect 18690 11880 18696 11892
rect 18555 11852 18696 11880
rect 18555 11849 18567 11852
rect 18509 11843 18567 11849
rect 18690 11840 18696 11852
rect 18748 11880 18754 11892
rect 19153 11883 19211 11889
rect 19153 11880 19165 11883
rect 18748 11852 19165 11880
rect 18748 11840 18754 11852
rect 19153 11849 19165 11852
rect 19199 11849 19211 11883
rect 24026 11880 24032 11892
rect 19153 11843 19211 11849
rect 19996 11852 24032 11880
rect 18414 11812 18420 11824
rect 16071 11784 17724 11812
rect 18064 11784 18420 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 11609 11707 11667 11713
rect 12406 11716 13124 11744
rect 13173 11747 13231 11753
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11645 2191 11679
rect 2133 11639 2191 11645
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 5626 11676 5632 11688
rect 4755 11648 5632 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 1946 11568 1952 11620
rect 2004 11608 2010 11620
rect 2148 11608 2176 11639
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5902 11636 5908 11688
rect 5960 11636 5966 11688
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 8680 11648 10333 11676
rect 4890 11608 4896 11620
rect 2004 11580 4896 11608
rect 2004 11568 2010 11580
rect 4890 11568 4896 11580
rect 4948 11568 4954 11620
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5920 11608 5948 11636
rect 5592 11580 5948 11608
rect 5592 11568 5598 11580
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4982 11540 4988 11552
rect 4111 11512 4988 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8680 11540 8708 11648
rect 10321 11645 10333 11648
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11676 11023 11679
rect 12406 11676 12434 11716
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 15930 11704 15936 11756
rect 15988 11704 15994 11756
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 17696 11744 17724 11784
rect 18414 11772 18420 11784
rect 18472 11772 18478 11824
rect 18601 11815 18659 11821
rect 18601 11781 18613 11815
rect 18647 11812 18659 11815
rect 18782 11812 18788 11824
rect 18647 11784 18788 11812
rect 18647 11781 18659 11784
rect 18601 11775 18659 11781
rect 18782 11772 18788 11784
rect 18840 11812 18846 11824
rect 19996 11821 20024 11852
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 19337 11815 19395 11821
rect 19337 11812 19349 11815
rect 18840 11784 19349 11812
rect 18840 11772 18846 11784
rect 19337 11781 19349 11784
rect 19383 11781 19395 11815
rect 19337 11775 19395 11781
rect 19981 11815 20039 11821
rect 19981 11781 19993 11815
rect 20027 11781 20039 11815
rect 19981 11775 20039 11781
rect 22649 11815 22707 11821
rect 22649 11781 22661 11815
rect 22695 11812 22707 11815
rect 22738 11812 22744 11824
rect 22695 11784 22744 11812
rect 22695 11781 22707 11784
rect 22649 11775 22707 11781
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 23934 11812 23940 11824
rect 23874 11784 23940 11812
rect 23934 11772 23940 11784
rect 23992 11812 23998 11824
rect 24397 11815 24455 11821
rect 24397 11812 24409 11815
rect 23992 11784 24409 11812
rect 23992 11772 23998 11784
rect 24397 11781 24409 11784
rect 24443 11781 24455 11815
rect 24397 11775 24455 11781
rect 19426 11744 19432 11756
rect 17696 11716 19432 11744
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 21114 11716 21220 11744
rect 21192 11688 21220 11716
rect 11011 11648 12434 11676
rect 12529 11679 12587 11685
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 14182 11676 14188 11688
rect 13495 11648 14188 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 9030 11568 9036 11620
rect 9088 11608 9094 11620
rect 9125 11611 9183 11617
rect 9125 11608 9137 11611
rect 9088 11580 9137 11608
rect 9088 11568 9094 11580
rect 9125 11577 9137 11580
rect 9171 11577 9183 11611
rect 10336 11608 10364 11639
rect 11514 11608 11520 11620
rect 10336 11580 11520 11608
rect 9125 11571 9183 11577
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 11790 11568 11796 11620
rect 11848 11608 11854 11620
rect 12544 11608 12572 11639
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 17034 11676 17040 11688
rect 16255 11648 17040 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 17034 11636 17040 11648
rect 17092 11636 17098 11688
rect 17586 11636 17592 11688
rect 17644 11636 17650 11688
rect 17770 11636 17776 11688
rect 17828 11676 17834 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 17828 11648 18705 11676
rect 17828 11636 17834 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 19702 11636 19708 11688
rect 19760 11636 19766 11688
rect 21174 11636 21180 11688
rect 21232 11676 21238 11688
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 21232 11648 21925 11676
rect 21232 11636 21238 11648
rect 21913 11645 21925 11648
rect 21959 11645 21971 11679
rect 21913 11639 21971 11645
rect 22186 11636 22192 11688
rect 22244 11676 22250 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 22244 11648 22385 11676
rect 22244 11636 22250 11648
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 22373 11639 22431 11645
rect 11848 11580 12572 11608
rect 11848 11568 11854 11580
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 13170 11608 13176 11620
rect 12676 11580 13176 11608
rect 12676 11568 12682 11580
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 16945 11611 17003 11617
rect 16945 11608 16957 11611
rect 15344 11580 16957 11608
rect 15344 11568 15350 11580
rect 16945 11577 16957 11580
rect 16991 11577 17003 11611
rect 16945 11571 17003 11577
rect 17218 11568 17224 11620
rect 17276 11608 17282 11620
rect 18141 11611 18199 11617
rect 18141 11608 18153 11611
rect 17276 11580 18153 11608
rect 17276 11568 17282 11580
rect 18141 11577 18153 11580
rect 18187 11577 18199 11611
rect 18141 11571 18199 11577
rect 7892 11512 8708 11540
rect 7892 11500 7898 11512
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 10226 11540 10232 11552
rect 8812 11512 10232 11540
rect 8812 11500 8818 11512
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 11204 11512 11989 11540
rect 11204 11500 11210 11512
rect 11977 11509 11989 11512
rect 12023 11509 12035 11543
rect 11977 11503 12035 11509
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 12124 11512 14933 11540
rect 12124 11500 12130 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 19150 11540 19156 11552
rect 15611 11512 19156 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 21450 11500 21456 11552
rect 21508 11500 21514 11552
rect 23382 11500 23388 11552
rect 23440 11540 23446 11552
rect 24121 11543 24179 11549
rect 24121 11540 24133 11543
rect 23440 11512 24133 11540
rect 23440 11500 23446 11512
rect 24121 11509 24133 11512
rect 24167 11540 24179 11543
rect 25130 11540 25136 11552
rect 24167 11512 25136 11540
rect 24167 11509 24179 11512
rect 24121 11503 24179 11509
rect 25130 11500 25136 11512
rect 25188 11500 25194 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 3605 11339 3663 11345
rect 3605 11305 3617 11339
rect 3651 11336 3663 11339
rect 3694 11336 3700 11348
rect 3651 11308 3700 11336
rect 3651 11305 3663 11308
rect 3605 11299 3663 11305
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 5626 11336 5632 11348
rect 4203 11308 5632 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 5776 11308 6561 11336
rect 5776 11296 5782 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 7466 11296 7472 11348
rect 7524 11296 7530 11348
rect 7837 11339 7895 11345
rect 7837 11305 7849 11339
rect 7883 11336 7895 11339
rect 10594 11336 10600 11348
rect 7883 11308 10600 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11606 11296 11612 11348
rect 11664 11336 11670 11348
rect 12250 11336 12256 11348
rect 11664 11308 12256 11336
rect 11664 11296 11670 11308
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 12400 11308 13277 11336
rect 12400 11296 12406 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13354 11296 13360 11348
rect 13412 11296 13418 11348
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13504 11308 13553 11336
rect 13504 11296 13510 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 13541 11299 13599 11305
rect 13817 11339 13875 11345
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 13906 11336 13912 11348
rect 13863 11308 13912 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 16485 11339 16543 11345
rect 16485 11305 16497 11339
rect 16531 11336 16543 11339
rect 16574 11336 16580 11348
rect 16531 11308 16580 11336
rect 16531 11305 16543 11308
rect 16485 11299 16543 11305
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 17402 11296 17408 11348
rect 17460 11336 17466 11348
rect 18598 11336 18604 11348
rect 17460 11308 18604 11336
rect 17460 11296 17466 11308
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 18966 11336 18972 11348
rect 18923 11308 18972 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11336 22707 11339
rect 22830 11336 22836 11348
rect 22695 11308 22836 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23017 11339 23075 11345
rect 23017 11305 23029 11339
rect 23063 11336 23075 11339
rect 23566 11336 23572 11348
rect 23063 11308 23572 11336
rect 23063 11305 23075 11308
rect 23017 11299 23075 11305
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 1627 11240 2774 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 2590 11200 2596 11212
rect 2271 11172 2596 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 1762 11092 1768 11144
rect 1820 11092 1826 11144
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2746 11132 2774 11240
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7156 11240 8432 11268
rect 7156 11228 7162 11240
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5534 11200 5540 11212
rect 5123 11172 5540 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5626 11160 5632 11212
rect 5684 11200 5690 11212
rect 7282 11200 7288 11212
rect 5684 11172 7288 11200
rect 5684 11160 5690 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8404 11209 8432 11240
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 10321 11271 10379 11277
rect 9088 11240 9720 11268
rect 9088 11228 9094 11240
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 7984 11172 8309 11200
rect 7984 11160 7990 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 9582 11160 9588 11212
rect 9640 11160 9646 11212
rect 9692 11209 9720 11240
rect 10321 11237 10333 11271
rect 10367 11268 10379 11271
rect 11330 11268 11336 11280
rect 10367 11240 11336 11268
rect 10367 11237 10379 11240
rect 10321 11231 10379 11237
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 13372 11268 13400 11296
rect 11440 11240 11652 11268
rect 13372 11240 14228 11268
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 2746 11104 4077 11132
rect 2501 11095 2559 11101
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 2516 11064 2544 11095
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 6454 11132 6460 11144
rect 6210 11104 6460 11132
rect 6454 11092 6460 11104
rect 6512 11132 6518 11144
rect 7466 11132 7472 11144
rect 6512 11104 7472 11132
rect 6512 11092 6518 11104
rect 7466 11092 7472 11104
rect 7524 11132 7530 11144
rect 8110 11132 8116 11144
rect 7524 11104 8116 11132
rect 7524 11092 7530 11104
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 9214 11132 9220 11144
rect 8251 11104 9220 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 10410 11132 10416 11144
rect 9539 11104 10416 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 1636 11036 2544 11064
rect 7009 11067 7067 11073
rect 1636 11024 1642 11036
rect 7009 11033 7021 11067
rect 7055 11064 7067 11067
rect 8754 11064 8760 11076
rect 7055 11036 8760 11064
rect 7055 11033 7067 11036
rect 7009 11027 7067 11033
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 9456 11036 10701 11064
rect 9456 11024 9462 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10980 11064 11008 11163
rect 11440 11064 11468 11240
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 11624 11200 11652 11240
rect 13354 11200 13360 11212
rect 11624 11172 13360 11200
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 14200 11209 14228 11240
rect 14185 11203 14243 11209
rect 14185 11169 14197 11203
rect 14231 11200 14243 11203
rect 21542 11200 21548 11212
rect 14231 11172 21548 11200
rect 14231 11169 14243 11172
rect 14185 11163 14243 11169
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 11793 11067 11851 11073
rect 11793 11064 11805 11067
rect 10980 11036 11805 11064
rect 10689 11027 10747 11033
rect 11793 11033 11805 11036
rect 11839 11033 11851 11067
rect 13906 11064 13912 11076
rect 13018 11036 13912 11064
rect 11793 11027 11851 11033
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 14752 11064 14780 11095
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16908 11104 17141 11132
rect 16908 11092 16914 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 18932 11104 19533 11132
rect 18932 11092 18938 11104
rect 19521 11101 19533 11104
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 14918 11064 14924 11076
rect 14608 11036 14924 11064
rect 14608 11024 14614 11036
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 15010 11024 15016 11076
rect 15068 11024 15074 11076
rect 16238 11036 16344 11064
rect 9125 10999 9183 11005
rect 9125 10965 9137 10999
rect 9171 10996 9183 10999
rect 9582 10996 9588 11008
rect 9171 10968 9588 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 10778 10956 10784 11008
rect 10836 10956 10842 11008
rect 15838 10956 15844 11008
rect 15896 10996 15902 11008
rect 16316 10996 16344 11036
rect 16482 11024 16488 11076
rect 16540 11064 16546 11076
rect 17402 11064 17408 11076
rect 16540 11036 17408 11064
rect 16540 11024 16546 11036
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 17862 11064 17868 11076
rect 17512 11036 17868 11064
rect 16761 10999 16819 11005
rect 16761 10996 16773 10999
rect 15896 10968 16773 10996
rect 15896 10956 15902 10968
rect 16761 10965 16773 10968
rect 16807 10996 16819 10999
rect 17512 10996 17540 11036
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 19760 11036 20269 11064
rect 19760 11024 19766 11036
rect 20257 11033 20269 11036
rect 20303 11064 20315 11067
rect 20916 11064 20944 11095
rect 22278 11092 22284 11144
rect 22336 11132 22342 11144
rect 23032 11132 23060 11299
rect 23566 11296 23572 11308
rect 23624 11336 23630 11348
rect 23934 11336 23940 11348
rect 23624 11308 23940 11336
rect 23624 11296 23630 11308
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 31846 11296 31852 11348
rect 31904 11336 31910 11348
rect 32033 11339 32091 11345
rect 32033 11336 32045 11339
rect 31904 11308 32045 11336
rect 31904 11296 31910 11308
rect 32033 11305 32045 11308
rect 32079 11305 32091 11339
rect 32033 11299 32091 11305
rect 26878 11160 26884 11212
rect 26936 11200 26942 11212
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 26936 11172 29745 11200
rect 26936 11160 26942 11172
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 31846 11132 31852 11144
rect 22336 11104 23060 11132
rect 31142 11104 31852 11132
rect 22336 11092 22342 11104
rect 31846 11092 31852 11104
rect 31904 11092 31910 11144
rect 20303 11036 20944 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 27614 11024 27620 11076
rect 27672 11064 27678 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 27672 11036 30021 11064
rect 27672 11024 27678 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 31294 11024 31300 11076
rect 31352 11064 31358 11076
rect 31757 11067 31815 11073
rect 31757 11064 31769 11067
rect 31352 11036 31769 11064
rect 31352 11024 31358 11036
rect 31757 11033 31769 11036
rect 31803 11064 31815 11067
rect 47854 11064 47860 11076
rect 31803 11036 47860 11064
rect 31803 11033 31815 11036
rect 31757 11027 31815 11033
rect 47854 11024 47860 11036
rect 47912 11024 47918 11076
rect 16807 10968 17540 10996
rect 16807 10965 16819 10968
rect 16761 10959 16819 10965
rect 18690 10956 18696 11008
rect 18748 10996 18754 11008
rect 21358 10996 21364 11008
rect 18748 10968 21364 10996
rect 18748 10956 18754 10968
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4488 10764 4813 10792
rect 4488 10752 4494 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 9861 10795 9919 10801
rect 5859 10764 9076 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 1489 10727 1547 10733
rect 1489 10693 1501 10727
rect 1535 10724 1547 10727
rect 2590 10724 2596 10736
rect 1535 10696 2596 10724
rect 1535 10693 1547 10696
rect 1489 10687 1547 10693
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 6730 10724 6736 10736
rect 2746 10696 6736 10724
rect 2746 10656 2774 10696
rect 6730 10684 6736 10696
rect 6788 10684 6794 10736
rect 8294 10684 8300 10736
rect 8352 10684 8358 10736
rect 9048 10724 9076 10764
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 13814 10792 13820 10804
rect 9907 10764 13820 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15286 10792 15292 10804
rect 14875 10764 15292 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 15436 10764 15577 10792
rect 15436 10752 15442 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 15565 10755 15623 10761
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 17092 10764 19257 10792
rect 17092 10752 17098 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 21450 10792 21456 10804
rect 19245 10755 19303 10761
rect 19628 10764 21456 10792
rect 10689 10727 10747 10733
rect 10689 10724 10701 10727
rect 9048 10696 10701 10724
rect 10689 10693 10701 10696
rect 10735 10693 10747 10727
rect 10689 10687 10747 10693
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 11146 10724 11152 10736
rect 10827 10696 11152 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 11146 10684 11152 10696
rect 11204 10724 11210 10736
rect 11974 10724 11980 10736
rect 11204 10696 11980 10724
rect 11204 10684 11210 10696
rect 11974 10684 11980 10696
rect 12032 10684 12038 10736
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12345 10727 12403 10733
rect 12345 10724 12357 10727
rect 12124 10696 12357 10724
rect 12124 10684 12130 10696
rect 12345 10693 12357 10696
rect 12391 10693 12403 10727
rect 13906 10724 13912 10736
rect 13570 10696 13912 10724
rect 12345 10687 12403 10693
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 16758 10684 16764 10736
rect 16816 10724 16822 10736
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 16816 10696 17785 10724
rect 16816 10684 16822 10696
rect 2148 10628 2774 10656
rect 3421 10659 3479 10665
rect 2148 10597 2176 10628
rect 3421 10625 3433 10659
rect 3467 10656 3479 10659
rect 5074 10656 5080 10668
rect 3467 10628 5080 10656
rect 3467 10625 3479 10628
rect 3421 10619 3479 10625
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5350 10616 5356 10668
rect 5408 10616 5414 10668
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 5684 10628 7021 10656
rect 5684 10616 5690 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10962 10656 10968 10668
rect 10376 10628 10968 10656
rect 10376 10616 10382 10628
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1903 10560 2145 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2133 10557 2145 10560
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 6914 10588 6920 10600
rect 3743 10560 6920 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 1026 10480 1032 10532
rect 1084 10520 1090 10532
rect 2424 10520 2452 10551
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7745 10591 7803 10597
rect 7515 10560 7604 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 1084 10492 2452 10520
rect 1084 10480 1090 10492
rect 2590 10480 2596 10532
rect 2648 10520 2654 10532
rect 4617 10523 4675 10529
rect 4617 10520 4629 10523
rect 2648 10492 4629 10520
rect 2648 10480 2654 10492
rect 4617 10489 4629 10492
rect 4663 10489 4675 10523
rect 6549 10523 6607 10529
rect 6549 10520 6561 10523
rect 4617 10483 4675 10489
rect 4724 10492 6561 10520
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 1946 10452 1952 10464
rect 1636 10424 1952 10452
rect 1636 10412 1642 10424
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 4724 10452 4752 10492
rect 6549 10489 6561 10492
rect 6595 10520 6607 10523
rect 7374 10520 7380 10532
rect 6595 10492 7380 10520
rect 6595 10489 6607 10492
rect 6549 10483 6607 10489
rect 7374 10480 7380 10492
rect 7432 10480 7438 10532
rect 3844 10424 4752 10452
rect 3844 10412 3850 10424
rect 5166 10412 5172 10464
rect 5224 10412 5230 10464
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6788 10424 6837 10452
rect 6788 10412 6794 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7466 10452 7472 10464
rect 6972 10424 7472 10452
rect 6972 10412 6978 10424
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 7576 10452 7604 10560
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8110 10588 8116 10600
rect 7791 10560 8116 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 10686 10588 10692 10600
rect 10091 10560 10692 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10888 10597 10916 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 10873 10591 10931 10597
rect 10873 10557 10885 10591
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11296 10560 12081 10588
rect 11296 10548 11302 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 14752 10588 14780 10619
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 15436 10628 15945 10656
rect 15436 10616 15442 10628
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 12069 10551 12127 10557
rect 12176 10560 14780 10588
rect 15013 10591 15071 10597
rect 10226 10480 10232 10532
rect 10284 10520 10290 10532
rect 12176 10520 12204 10560
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15194 10588 15200 10600
rect 15059 10560 15200 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10588 16083 10591
rect 16209 10591 16267 10597
rect 16071 10560 16160 10588
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 10284 10492 12204 10520
rect 10284 10480 10290 10492
rect 7834 10452 7840 10464
rect 7576 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 8260 10424 10333 10452
rect 8260 10412 8266 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11609 10455 11667 10461
rect 11609 10452 11621 10455
rect 11572 10424 11621 10452
rect 11572 10412 11578 10424
rect 11609 10421 11621 10424
rect 11655 10421 11667 10455
rect 11609 10415 11667 10421
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 11848 10424 13829 10452
rect 11848 10412 11854 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14369 10455 14427 10461
rect 14369 10421 14381 10455
rect 14415 10452 14427 10455
rect 16022 10452 16028 10464
rect 14415 10424 16028 10452
rect 14415 10421 14427 10424
rect 14369 10415 14427 10421
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16132 10452 16160 10560
rect 16209 10557 16221 10591
rect 16255 10588 16267 10591
rect 16298 10588 16304 10600
rect 16255 10560 16304 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16632 10560 16865 10588
rect 16632 10548 16638 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 17420 10588 17448 10696
rect 17773 10693 17785 10696
rect 17819 10693 17831 10727
rect 17773 10687 17831 10693
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 17920 10696 18262 10724
rect 17920 10684 17926 10696
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 19628 10588 19656 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21913 10795 21971 10801
rect 21913 10761 21925 10795
rect 21959 10792 21971 10795
rect 22097 10795 22155 10801
rect 22097 10792 22109 10795
rect 21959 10764 22109 10792
rect 21959 10761 21971 10764
rect 21913 10755 21971 10761
rect 22097 10761 22109 10764
rect 22143 10792 22155 10795
rect 22278 10792 22284 10804
rect 22143 10764 22284 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 21542 10724 21548 10736
rect 21206 10696 21548 10724
rect 21542 10684 21548 10696
rect 21600 10724 21606 10736
rect 21928 10724 21956 10755
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 21600 10696 21956 10724
rect 21600 10684 21606 10696
rect 17420 10560 19656 10588
rect 16853 10551 16911 10557
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 22830 10588 22836 10600
rect 20027 10560 22836 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 21358 10480 21364 10532
rect 21416 10520 21422 10532
rect 21453 10523 21511 10529
rect 21453 10520 21465 10523
rect 21416 10492 21465 10520
rect 21416 10480 21422 10492
rect 21453 10489 21465 10492
rect 21499 10489 21511 10523
rect 21453 10483 21511 10489
rect 20530 10452 20536 10464
rect 16132 10424 20536 10452
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 1210 10208 1216 10260
rect 1268 10248 1274 10260
rect 2685 10251 2743 10257
rect 2685 10248 2697 10251
rect 1268 10220 2697 10248
rect 1268 10208 1274 10220
rect 2685 10217 2697 10220
rect 2731 10217 2743 10251
rect 2685 10211 2743 10217
rect 2866 10208 2872 10260
rect 2924 10208 2930 10260
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3602 10248 3608 10260
rect 3283 10220 3608 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 4488 10220 5457 10248
rect 4488 10208 4494 10220
rect 5445 10217 5457 10220
rect 5491 10248 5503 10251
rect 6638 10248 6644 10260
rect 5491 10220 6644 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10778 10248 10784 10260
rect 10091 10220 10784 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 12158 10248 12164 10260
rect 11020 10220 12164 10248
rect 11020 10208 11026 10220
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13964 10220 14105 10248
rect 13964 10208 13970 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 15010 10208 15016 10260
rect 15068 10248 15074 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 15068 10220 16313 10248
rect 15068 10208 15074 10220
rect 16301 10217 16313 10220
rect 16347 10248 16359 10251
rect 17770 10248 17776 10260
rect 16347 10220 17776 10248
rect 16347 10217 16359 10220
rect 16301 10211 16359 10217
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 19794 10248 19800 10260
rect 18932 10220 19800 10248
rect 18932 10208 18938 10220
rect 19794 10208 19800 10220
rect 19852 10208 19858 10260
rect 21542 10208 21548 10260
rect 21600 10208 21606 10260
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1670 10112 1676 10124
rect 1627 10084 1676 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 2884 10112 2912 10208
rect 3418 10140 3424 10192
rect 3476 10180 3482 10192
rect 3881 10183 3939 10189
rect 3881 10180 3893 10183
rect 3476 10152 3893 10180
rect 3476 10140 3482 10152
rect 3881 10149 3893 10152
rect 3927 10149 3939 10183
rect 3881 10143 3939 10149
rect 6365 10183 6423 10189
rect 6365 10149 6377 10183
rect 6411 10180 6423 10183
rect 6454 10180 6460 10192
rect 6411 10152 6460 10180
rect 6411 10149 6423 10152
rect 6365 10143 6423 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 8573 10183 8631 10189
rect 8573 10180 8585 10183
rect 8168 10152 8585 10180
rect 8168 10140 8174 10152
rect 8573 10149 8585 10152
rect 8619 10180 8631 10183
rect 10870 10180 10876 10192
rect 8619 10152 10876 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 3510 10112 3516 10124
rect 1903 10084 3516 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 4246 10072 4252 10124
rect 4304 10072 4310 10124
rect 4522 10072 4528 10124
rect 4580 10072 4586 10124
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 6825 10115 6883 10121
rect 6825 10112 6837 10115
rect 4856 10084 6837 10112
rect 4856 10072 4862 10084
rect 6825 10081 6837 10084
rect 6871 10112 6883 10115
rect 7834 10112 7840 10124
rect 6871 10084 7840 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 8294 10112 8300 10124
rect 8220 10084 8300 10112
rect 1688 9976 1716 10072
rect 2682 10004 2688 10056
rect 2740 10044 2746 10056
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2740 10016 2881 10044
rect 2740 10004 2746 10016
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3418 10044 3424 10056
rect 3191 10016 3424 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 5810 10004 5816 10056
rect 5868 10004 5874 10056
rect 8220 10030 8248 10084
rect 8294 10072 8300 10084
rect 8352 10112 8358 10124
rect 9030 10112 9036 10124
rect 8352 10084 9036 10112
rect 8352 10072 8358 10084
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 11974 10112 11980 10124
rect 10735 10084 11980 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 12636 10084 12848 10112
rect 12636 10056 12664 10084
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 10962 10044 10968 10056
rect 9447 10016 10968 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11238 10004 11244 10056
rect 11296 10004 11302 10056
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 4614 9976 4620 9988
rect 1688 9948 4620 9976
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 7374 9976 7380 9988
rect 7156 9948 7380 9976
rect 7156 9936 7162 9948
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 11517 9979 11575 9985
rect 11517 9945 11529 9979
rect 11563 9976 11575 9979
rect 11790 9976 11796 9988
rect 11563 9948 11796 9976
rect 11563 9945 11575 9948
rect 11517 9939 11575 9945
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 12820 9976 12848 10084
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 14550 10072 14556 10124
rect 14608 10072 14614 10124
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 15194 10112 15200 10124
rect 14875 10084 15200 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15194 10072 15200 10084
rect 15252 10112 15258 10124
rect 16206 10112 16212 10124
rect 15252 10084 16212 10112
rect 15252 10072 15258 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 17144 10084 19441 10112
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17144 10053 17172 10084
rect 19429 10081 19441 10084
rect 19475 10112 19487 10115
rect 19702 10112 19708 10124
rect 19475 10084 19708 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16908 10016 17141 10044
rect 16908 10004 16914 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 21542 10044 21548 10056
rect 20772 10016 21548 10044
rect 20772 10004 20778 10016
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 13906 9976 13912 9988
rect 12742 9948 13912 9976
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 16054 9948 16712 9976
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 3786 9908 3792 9920
rect 2464 9880 3792 9908
rect 2464 9868 2470 9880
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 8444 9880 10425 9908
rect 8444 9868 8450 9880
rect 10413 9877 10425 9880
rect 10459 9877 10471 9911
rect 10413 9871 10471 9877
rect 10505 9911 10563 9917
rect 10505 9877 10517 9911
rect 10551 9908 10563 9911
rect 11422 9908 11428 9920
rect 10551 9880 11428 9908
rect 10551 9877 10563 9880
rect 10505 9871 10563 9877
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 11940 9880 13001 9908
rect 11940 9868 11946 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 16132 9908 16160 9948
rect 16684 9917 16712 9948
rect 17034 9936 17040 9988
rect 17092 9976 17098 9988
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 17092 9948 17417 9976
rect 17092 9936 17098 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 17512 9948 17894 9976
rect 15252 9880 16160 9908
rect 16669 9911 16727 9917
rect 15252 9868 15258 9880
rect 16669 9877 16681 9911
rect 16715 9908 16727 9911
rect 16853 9911 16911 9917
rect 16853 9908 16865 9911
rect 16715 9880 16865 9908
rect 16715 9877 16727 9880
rect 16669 9871 16727 9877
rect 16853 9877 16865 9880
rect 16899 9908 16911 9911
rect 17512 9908 17540 9948
rect 19242 9936 19248 9988
rect 19300 9976 19306 9988
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 19300 9948 19717 9976
rect 19300 9936 19306 9948
rect 19705 9945 19717 9948
rect 19751 9945 19763 9979
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 19705 9939 19763 9945
rect 21008 9948 21649 9976
rect 16899 9880 17540 9908
rect 19720 9908 19748 9939
rect 21008 9908 21036 9948
rect 21637 9945 21649 9948
rect 21683 9976 21695 9979
rect 23382 9976 23388 9988
rect 21683 9948 23388 9976
rect 21683 9945 21695 9948
rect 21637 9939 21695 9945
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 19720 9880 21036 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 21174 9868 21180 9920
rect 21232 9868 21238 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 6454 9664 6460 9716
rect 6512 9664 6518 9716
rect 7650 9664 7656 9716
rect 7708 9704 7714 9716
rect 15470 9704 15476 9716
rect 7708 9676 15476 9704
rect 7708 9664 7714 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 16206 9664 16212 9716
rect 16264 9664 16270 9716
rect 18874 9704 18880 9716
rect 17512 9676 18880 9704
rect 1486 9596 1492 9648
rect 1544 9596 1550 9648
rect 1673 9639 1731 9645
rect 1673 9605 1685 9639
rect 1719 9636 1731 9639
rect 1762 9636 1768 9648
rect 1719 9608 1768 9636
rect 1719 9605 1731 9608
rect 1673 9599 1731 9605
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5767 9608 5825 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 5813 9605 5825 9608
rect 5859 9636 5871 9639
rect 5902 9636 5908 9648
rect 5859 9608 5908 9636
rect 5859 9605 5871 9608
rect 5813 9599 5871 9605
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 8478 9636 8484 9648
rect 7208 9608 8484 9636
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 3786 9528 3792 9580
rect 3844 9528 3850 9580
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 5166 9568 5172 9580
rect 4295 9540 5172 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 5500 9540 7113 9568
rect 5500 9528 5506 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2314 9500 2320 9512
rect 2004 9472 2320 9500
rect 2004 9460 2010 9472
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9469 4583 9503
rect 4525 9463 4583 9469
rect 3602 9392 3608 9444
rect 3660 9392 3666 9444
rect 4540 9432 4568 9463
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 7208 9432 7236 9608
rect 8478 9596 8484 9608
rect 8536 9596 8542 9648
rect 9030 9596 9036 9648
rect 9088 9596 9094 9648
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 10781 9639 10839 9645
rect 10781 9636 10793 9639
rect 10652 9608 10793 9636
rect 10652 9596 10658 9608
rect 10781 9605 10793 9608
rect 10827 9605 10839 9639
rect 10781 9599 10839 9605
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 12618 9596 12624 9648
rect 12676 9596 12682 9648
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 13909 9639 13967 9645
rect 13909 9636 13921 9639
rect 13872 9608 13921 9636
rect 13872 9596 13878 9608
rect 13909 9605 13921 9608
rect 13955 9636 13967 9639
rect 15194 9636 15200 9648
rect 13955 9608 15200 9636
rect 13955 9605 13967 9608
rect 13909 9599 13967 9605
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 16022 9596 16028 9648
rect 16080 9636 16086 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 16080 9608 17141 9636
rect 16080 9596 16086 9608
rect 17129 9605 17141 9608
rect 17175 9636 17187 9639
rect 17512 9636 17540 9676
rect 18874 9664 18880 9676
rect 18932 9664 18938 9716
rect 18506 9636 18512 9648
rect 17175 9608 17540 9636
rect 18354 9608 18512 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 18506 9596 18512 9608
rect 18564 9596 18570 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 24578 9636 24584 9648
rect 19567 9608 24584 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 24578 9596 24584 9608
rect 24636 9596 24642 9648
rect 27798 9596 27804 9648
rect 27856 9636 27862 9648
rect 28629 9639 28687 9645
rect 28629 9636 28641 9639
rect 27856 9608 28641 9636
rect 27856 9596 27862 9608
rect 28629 9605 28641 9608
rect 28675 9636 28687 9639
rect 31294 9636 31300 9648
rect 28675 9608 31300 9636
rect 28675 9605 28687 9608
rect 28629 9599 28687 9605
rect 31294 9596 31300 9608
rect 31352 9596 31358 9648
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9732 9540 10701 9568
rect 9732 9528 9738 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7892 9472 8125 9500
rect 7892 9460 7898 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 10318 9500 10324 9512
rect 8435 9472 10324 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10870 9460 10876 9512
rect 10928 9460 10934 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11296 9472 11713 9500
rect 11296 9460 11302 9472
rect 11701 9469 11713 9472
rect 11747 9500 11759 9503
rect 14458 9500 14464 9512
rect 11747 9472 14464 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14734 9460 14740 9512
rect 14792 9460 14798 9512
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 16758 9500 16764 9512
rect 15344 9472 16764 9500
rect 15344 9460 15350 9472
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 19444 9500 19472 9531
rect 23750 9528 23756 9580
rect 23808 9568 23814 9580
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 23808 9540 27537 9568
rect 23808 9528 23814 9540
rect 27525 9537 27537 9540
rect 27571 9568 27583 9571
rect 27571 9540 28488 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 17276 9472 19472 9500
rect 19705 9503 19763 9509
rect 17276 9460 17282 9472
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 21174 9500 21180 9512
rect 19751 9472 21180 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 23440 9472 27997 9500
rect 23440 9460 23446 9472
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 27985 9463 28043 9469
rect 4540 9404 7236 9432
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 13412 9404 13461 9432
rect 13412 9392 13418 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 13449 9395 13507 9401
rect 13648 9404 14105 9432
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5626 9364 5632 9376
rect 5583 9336 5632 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 8110 9364 8116 9376
rect 7432 9336 8116 9364
rect 7432 9324 7438 9336
rect 8110 9324 8116 9336
rect 8168 9364 8174 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 8168 9336 9873 9364
rect 8168 9324 8174 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9364 10379 9367
rect 11422 9364 11428 9376
rect 10367 9336 11428 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 13538 9364 13544 9376
rect 12492 9336 13544 9364
rect 12492 9324 12498 9336
rect 13538 9324 13544 9336
rect 13596 9364 13602 9376
rect 13648 9364 13676 9404
rect 14093 9401 14105 9404
rect 14139 9401 14151 9435
rect 14093 9395 14151 9401
rect 18506 9392 18512 9444
rect 18564 9432 18570 9444
rect 18564 9404 19012 9432
rect 18564 9392 18570 9404
rect 13596 9336 13676 9364
rect 13596 9324 13602 9336
rect 13998 9324 14004 9376
rect 14056 9364 14062 9376
rect 15746 9364 15752 9376
rect 14056 9336 15752 9364
rect 14056 9324 14062 9336
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 16356 9336 18613 9364
rect 16356 9324 16362 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18984 9364 19012 9404
rect 19058 9392 19064 9444
rect 19116 9392 19122 9444
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 18984 9336 20085 9364
rect 18601 9327 18659 9333
rect 20073 9333 20085 9336
rect 20119 9364 20131 9367
rect 20714 9364 20720 9376
rect 20119 9336 20720 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 27798 9324 27804 9376
rect 27856 9324 27862 9376
rect 28460 9373 28488 9540
rect 28445 9367 28503 9373
rect 28445 9333 28457 9367
rect 28491 9364 28503 9367
rect 31570 9364 31576 9376
rect 28491 9336 31576 9364
rect 28491 9333 28503 9336
rect 28445 9327 28503 9333
rect 31570 9324 31576 9336
rect 31628 9324 31634 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 3421 9163 3479 9169
rect 3421 9129 3433 9163
rect 3467 9160 3479 9163
rect 3786 9160 3792 9172
rect 3467 9132 3792 9160
rect 3467 9129 3479 9132
rect 3421 9123 3479 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 5258 9160 5264 9172
rect 4663 9132 5264 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 3605 9095 3663 9101
rect 3605 9061 3617 9095
rect 3651 9092 3663 9095
rect 4062 9092 4068 9104
rect 3651 9064 4068 9092
rect 3651 9061 3663 9064
rect 3605 9055 3663 9061
rect 4062 9052 4068 9064
rect 4120 9052 4126 9104
rect 1578 8984 1584 9036
rect 1636 8984 1642 9036
rect 1854 8984 1860 9036
rect 1912 8984 1918 9036
rect 4724 9033 4752 9132
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 5534 9120 5540 9172
rect 5592 9120 5598 9172
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 9674 9160 9680 9172
rect 7883 9132 9680 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10134 9120 10140 9172
rect 10192 9120 10198 9172
rect 11563 9163 11621 9169
rect 11563 9129 11575 9163
rect 11609 9160 11621 9163
rect 32398 9160 32404 9172
rect 11609 9132 32404 9160
rect 11609 9129 11621 9132
rect 11563 9123 11621 9129
rect 32398 9120 32404 9132
rect 32456 9120 32462 9172
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 5169 9095 5227 9101
rect 5169 9092 5181 9095
rect 4948 9064 5181 9092
rect 4948 9052 4954 9064
rect 5169 9061 5181 9064
rect 5215 9061 5227 9095
rect 5169 9055 5227 9061
rect 5276 9064 6316 9092
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 1596 8956 1624 8984
rect 1596 8928 2774 8956
rect 2746 8888 2774 8928
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2924 8928 3065 8956
rect 2924 8916 2930 8928
rect 3053 8925 3065 8928
rect 3099 8956 3111 8959
rect 3418 8956 3424 8968
rect 3099 8928 3424 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 5276 8956 5304 9064
rect 6178 8984 6184 9036
rect 6236 8984 6242 9036
rect 6288 9024 6316 9064
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 13630 9092 13636 9104
rect 6880 9064 13636 9092
rect 6880 9052 6886 9064
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 14277 9095 14335 9101
rect 14277 9061 14289 9095
rect 14323 9092 14335 9095
rect 15930 9092 15936 9104
rect 14323 9064 15936 9092
rect 14323 9061 14335 9064
rect 14277 9055 14335 9061
rect 15930 9052 15936 9064
rect 15988 9052 15994 9104
rect 6288 8996 7880 9024
rect 4304 8928 5304 8956
rect 5905 8959 5963 8965
rect 4304 8916 4310 8928
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7742 8956 7748 8968
rect 7423 8928 7748 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 3234 8888 3240 8900
rect 2746 8860 3240 8888
rect 3234 8848 3240 8860
rect 3292 8848 3298 8900
rect 4706 8888 4712 8900
rect 3436 8860 4712 8888
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 3436 8820 3464 8860
rect 4706 8848 4712 8860
rect 4764 8848 4770 8900
rect 5920 8888 5948 8919
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 7852 8956 7880 8996
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8168 8996 8401 9024
rect 8168 8984 8174 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 9024 10839 9027
rect 10827 8996 12434 9024
rect 10827 8993 10839 8996
rect 10781 8987 10839 8993
rect 8662 8956 8668 8968
rect 7852 8928 8668 8956
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 11330 8916 11336 8968
rect 11388 8916 11394 8968
rect 12406 8956 12434 8996
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 13596 8996 14749 9024
rect 13596 8984 13602 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 9024 14979 9027
rect 15286 9024 15292 9036
rect 14967 8996 15292 9024
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 15838 9024 15844 9036
rect 15528 8996 15844 9024
rect 15528 8984 15534 8996
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16850 9024 16856 9036
rect 16071 8996 16856 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 15010 8956 15016 8968
rect 12406 8928 15016 8956
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 9122 8888 9128 8900
rect 5920 8860 9128 8888
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 10505 8891 10563 8897
rect 10505 8857 10517 8891
rect 10551 8888 10563 8891
rect 11882 8888 11888 8900
rect 10551 8860 11888 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 13541 8891 13599 8897
rect 13541 8857 13553 8891
rect 13587 8857 13599 8891
rect 13541 8851 13599 8857
rect 2915 8792 3464 8820
rect 3973 8823 4031 8829
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 7650 8820 7656 8832
rect 4019 8792 7656 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 8202 8780 8208 8832
rect 8260 8780 8266 8832
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 9030 8780 9036 8832
rect 9088 8780 9094 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 9732 8792 10609 8820
rect 9732 8780 9738 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10597 8783 10655 8789
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 11606 8820 11612 8832
rect 11296 8792 11612 8820
rect 11296 8780 11302 8792
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 12492 8792 12633 8820
rect 12492 8780 12498 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 13556 8820 13584 8851
rect 16298 8848 16304 8900
rect 16356 8848 16362 8900
rect 17526 8860 18184 8888
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 13556 8792 14657 8820
rect 12621 8783 12679 8789
rect 14645 8789 14657 8792
rect 14691 8789 14703 8823
rect 14645 8783 14703 8789
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 17586 8820 17592 8832
rect 14792 8792 17592 8820
rect 14792 8780 14798 8792
rect 17586 8780 17592 8792
rect 17644 8820 17650 8832
rect 18156 8829 18184 8860
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17644 8792 17785 8820
rect 17644 8780 17650 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17773 8783 17831 8789
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18506 8820 18512 8832
rect 18187 8792 18512 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18506 8780 18512 8792
rect 18564 8820 18570 8832
rect 18693 8823 18751 8829
rect 18693 8820 18705 8823
rect 18564 8792 18705 8820
rect 18564 8780 18570 8792
rect 18693 8789 18705 8792
rect 18739 8820 18751 8823
rect 18969 8823 19027 8829
rect 18969 8820 18981 8823
rect 18739 8792 18981 8820
rect 18739 8789 18751 8792
rect 18693 8783 18751 8789
rect 18969 8789 18981 8792
rect 19015 8789 19027 8823
rect 18969 8783 19027 8789
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3326 8616 3332 8628
rect 2915 8588 3332 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 3510 8576 3516 8628
rect 3568 8576 3574 8628
rect 3970 8576 3976 8628
rect 4028 8576 4034 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5132 8588 5825 8616
rect 5132 8576 5138 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 6454 8576 6460 8628
rect 6512 8576 6518 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7800 8588 8033 8616
rect 7800 8576 7806 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8168 8588 10180 8616
rect 8168 8576 8174 8588
rect 1118 8508 1124 8560
rect 1176 8548 1182 8560
rect 7377 8551 7435 8557
rect 1176 8520 6040 8548
rect 1176 8508 1182 8520
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1857 8483 1915 8489
rect 1857 8480 1869 8483
rect 1452 8452 1869 8480
rect 1452 8440 1458 8452
rect 1857 8449 1869 8452
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3694 8480 3700 8492
rect 3099 8452 3700 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4246 8480 4252 8492
rect 4203 8452 4252 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 6012 8489 6040 8520
rect 7377 8517 7389 8551
rect 7423 8548 7435 8551
rect 10042 8548 10048 8560
rect 7423 8520 10048 8548
rect 7423 8517 7435 8520
rect 7377 8511 7435 8517
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 10152 8548 10180 8588
rect 11146 8576 11152 8628
rect 11204 8576 11210 8628
rect 11514 8576 11520 8628
rect 11572 8576 11578 8628
rect 12161 8619 12219 8625
rect 12161 8585 12173 8619
rect 12207 8616 12219 8619
rect 13998 8616 14004 8628
rect 12207 8588 14004 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 15378 8616 15384 8628
rect 14323 8588 15384 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8585 15623 8619
rect 15565 8579 15623 8585
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16574 8616 16580 8628
rect 15979 8588 16580 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 11238 8548 11244 8560
rect 10152 8520 11244 8548
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 14734 8548 14740 8560
rect 11532 8520 14740 8548
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7193 8483 7251 8489
rect 6871 8452 7144 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 1302 8372 1308 8424
rect 1360 8412 1366 8424
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 1360 8384 1593 8412
rect 1360 8372 1366 8384
rect 1581 8381 1593 8384
rect 1627 8412 1639 8415
rect 3326 8412 3332 8424
rect 1627 8384 3332 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 4816 8412 4844 8443
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4816 8384 5181 8412
rect 5169 8381 5181 8384
rect 5215 8412 5227 8415
rect 7006 8412 7012 8424
rect 5215 8384 7012 8412
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 4617 8347 4675 8353
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 6914 8344 6920 8356
rect 4663 8316 6920 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7116 8344 7144 8452
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 7558 8480 7564 8492
rect 7239 8452 7564 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 7558 8440 7564 8452
rect 7616 8480 7622 8492
rect 8665 8483 8723 8489
rect 7616 8452 8524 8480
rect 7616 8440 7622 8452
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8110 8412 8116 8424
rect 7791 8384 8116 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8496 8412 8524 8452
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 8754 8480 8760 8492
rect 8711 8452 8760 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 9030 8440 9036 8492
rect 9088 8480 9094 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 9088 8452 9689 8480
rect 9088 8440 9094 8452
rect 9677 8449 9689 8452
rect 9723 8480 9735 8483
rect 10410 8480 10416 8492
rect 9723 8452 10416 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 8496 8384 9996 8412
rect 8389 8375 8447 8381
rect 8404 8344 8432 8375
rect 9858 8344 9864 8356
rect 7116 8316 8340 8344
rect 8404 8316 9864 8344
rect 2222 8236 2228 8288
rect 2280 8276 2286 8288
rect 4430 8276 4436 8288
rect 2280 8248 4436 8276
rect 2280 8236 2286 8248
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7524 8248 7849 8276
rect 7524 8236 7530 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 8312 8276 8340 8316
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 9968 8344 9996 8384
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11532 8412 11560 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12492 8452 12541 8480
rect 12492 8440 12498 8452
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13679 8452 14657 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 15580 8480 15608 8579
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 15838 8508 15844 8560
rect 15896 8548 15902 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 15896 8520 16037 8548
rect 15896 8508 15902 8520
rect 16025 8517 16037 8520
rect 16071 8517 16083 8551
rect 16025 8511 16083 8517
rect 20438 8480 20444 8492
rect 15580 8452 20444 8480
rect 14645 8443 14703 8449
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 10827 8384 11560 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 12618 8372 12624 8424
rect 12676 8372 12682 8424
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8412 12863 8415
rect 12851 8384 14136 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 12526 8344 12532 8356
rect 9968 8316 12532 8344
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 14108 8344 14136 8384
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 14240 8384 14749 8412
rect 14240 8372 14246 8384
rect 14737 8381 14749 8384
rect 14783 8381 14795 8415
rect 14737 8375 14795 8381
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8412 14979 8415
rect 16022 8412 16028 8424
rect 14967 8384 16028 8412
rect 14967 8381 14979 8384
rect 14921 8375 14979 8381
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 20346 8412 20352 8424
rect 16255 8384 20352 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 16482 8344 16488 8356
rect 14108 8316 16488 8344
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 8478 8276 8484 8288
rect 8312 8248 8484 8276
rect 7837 8239 7895 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 10137 8279 10195 8285
rect 10137 8245 10149 8279
rect 10183 8276 10195 8279
rect 10226 8276 10232 8288
rect 10183 8248 10232 8276
rect 10183 8245 10195 8248
rect 10137 8239 10195 8245
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 16390 8276 16396 8288
rect 12860 8248 16396 8276
rect 12860 8236 12866 8248
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1946 8072 1952 8084
rect 1627 8044 1952 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2222 8032 2228 8084
rect 2280 8032 2286 8084
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 3786 8072 3792 8084
rect 2915 8044 3792 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 3878 8032 3884 8084
rect 3936 8032 3942 8084
rect 4246 8032 4252 8084
rect 4304 8032 4310 8084
rect 4614 8032 4620 8084
rect 4672 8032 4678 8084
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 8352 8044 9597 8072
rect 8352 8032 8358 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 12437 8075 12495 8081
rect 12437 8072 12449 8075
rect 9585 8035 9643 8041
rect 11256 8044 12449 8072
rect 2590 7964 2596 8016
rect 2648 8004 2654 8016
rect 3973 8007 4031 8013
rect 3973 8004 3985 8007
rect 2648 7976 3985 8004
rect 2648 7964 2654 7976
rect 3973 7973 3985 7976
rect 4019 7973 4031 8007
rect 3973 7967 4031 7973
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 6788 7976 11192 8004
rect 6788 7964 6794 7976
rect 2222 7896 2228 7948
rect 2280 7936 2286 7948
rect 2280 7908 5580 7936
rect 2280 7896 2286 7908
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 2590 7868 2596 7880
rect 2455 7840 2596 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 1780 7800 1808 7831
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2924 7840 3065 7868
rect 2924 7828 2930 7840
rect 3053 7837 3065 7840
rect 3099 7868 3111 7871
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 3099 7840 4445 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 5552 7868 5580 7908
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7340 7908 7757 7936
rect 7340 7896 7346 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7936 10287 7939
rect 10318 7936 10324 7948
rect 10275 7908 10324 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 8570 7868 8576 7880
rect 5552 7840 8576 7868
rect 4433 7831 4491 7837
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 11054 7868 11060 7880
rect 10091 7840 11060 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11164 7868 11192 7976
rect 11256 7945 11284 8044
rect 12437 8041 12449 8044
rect 12483 8072 12495 8075
rect 12802 8072 12808 8084
rect 12483 8044 12808 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 17218 8072 17224 8084
rect 13035 8044 17224 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 11348 7976 14872 8004
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7905 11299 7939
rect 11241 7899 11299 7905
rect 11348 7868 11376 7976
rect 14844 7945 14872 7976
rect 15194 7964 15200 8016
rect 15252 7964 15258 8016
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13679 7908 14289 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14829 7939 14887 7945
rect 14829 7905 14841 7939
rect 14875 7905 14887 7939
rect 19242 7936 19248 7948
rect 14829 7899 14887 7905
rect 14936 7908 19248 7936
rect 14182 7868 14188 7880
rect 11164 7840 11376 7868
rect 11624 7840 14188 7868
rect 3326 7800 3332 7812
rect 1780 7772 3332 7800
rect 3326 7760 3332 7772
rect 3384 7760 3390 7812
rect 3421 7803 3479 7809
rect 3421 7769 3433 7803
rect 3467 7800 3479 7803
rect 3467 7772 3648 7800
rect 3467 7769 3479 7772
rect 3421 7763 3479 7769
rect 3234 7692 3240 7744
rect 3292 7732 3298 7744
rect 3513 7735 3571 7741
rect 3513 7732 3525 7735
rect 3292 7704 3525 7732
rect 3292 7692 3298 7704
rect 3513 7701 3525 7704
rect 3559 7701 3571 7735
rect 3620 7732 3648 7772
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 9217 7803 9275 7809
rect 9217 7800 9229 7803
rect 6880 7772 9229 7800
rect 6880 7760 6886 7772
rect 9217 7769 9229 7772
rect 9263 7800 9275 7803
rect 9953 7803 10011 7809
rect 9953 7800 9965 7803
rect 9263 7772 9965 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 9953 7769 9965 7772
rect 9999 7800 10011 7803
rect 11624 7800 11652 7840
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14292 7868 14320 7899
rect 14936 7868 14964 7908
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 14292 7840 14964 7868
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15059 7840 15884 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 9999 7772 11652 7800
rect 9999 7769 10011 7772
rect 9953 7763 10011 7769
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 15028 7800 15056 7831
rect 12124 7772 15056 7800
rect 12124 7760 12130 7772
rect 3694 7732 3700 7744
rect 3620 7704 3700 7732
rect 3513 7695 3571 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 11471 7735 11529 7741
rect 11471 7732 11483 7735
rect 5684 7704 11483 7732
rect 5684 7692 5690 7704
rect 11471 7701 11483 7704
rect 11517 7701 11529 7735
rect 11471 7695 11529 7701
rect 13354 7692 13360 7744
rect 13412 7692 13418 7744
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 15856 7741 15884 7840
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 22830 7732 22836 7744
rect 15887 7704 22836 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 22830 7692 22836 7704
rect 22888 7732 22894 7744
rect 23382 7732 23388 7744
rect 22888 7704 23388 7732
rect 22888 7692 22894 7704
rect 23382 7692 23388 7704
rect 23440 7692 23446 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1670 7528 1676 7540
rect 1627 7500 1676 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 4062 7528 4068 7540
rect 1780 7500 4068 7528
rect 1780 7401 1808 7500
rect 4062 7488 4068 7500
rect 4120 7528 4126 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4120 7500 4353 7528
rect 4120 7488 4126 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 11698 7528 11704 7540
rect 9232 7500 11704 7528
rect 1872 7432 3740 7460
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 1302 7284 1308 7336
rect 1360 7324 1366 7336
rect 1872 7324 1900 7432
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3326 7392 3332 7404
rect 3099 7364 3332 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 1360 7296 1900 7324
rect 2424 7324 2452 7355
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 3712 7401 3740 7432
rect 3786 7420 3792 7472
rect 3844 7460 3850 7472
rect 9232 7460 9260 7500
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 11882 7488 11888 7540
rect 11940 7488 11946 7540
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13412 7500 13461 7528
rect 13412 7488 13418 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 27614 7528 27620 7540
rect 23992 7500 27620 7528
rect 23992 7488 23998 7500
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 3844 7432 9260 7460
rect 3844 7420 3850 7432
rect 9582 7420 9588 7472
rect 9640 7460 9646 7472
rect 9640 7432 10916 7460
rect 9640 7420 9646 7432
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3973 7395 4031 7401
rect 3973 7392 3985 7395
rect 3743 7364 3985 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3973 7361 3985 7364
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10888 7392 10916 7432
rect 11422 7420 11428 7472
rect 11480 7460 11486 7472
rect 11480 7432 14320 7460
rect 11480 7420 11486 7432
rect 14292 7401 14320 7432
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 10888 7364 12725 7392
rect 10781 7355 10839 7361
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 2682 7324 2688 7336
rect 2424 7296 2688 7324
rect 1360 7284 1366 7296
rect 2682 7284 2688 7296
rect 2740 7324 2746 7336
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 2740 7296 4169 7324
rect 2740 7284 2746 7296
rect 4157 7293 4169 7296
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 4982 7284 4988 7336
rect 5040 7324 5046 7336
rect 10796 7324 10824 7355
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 23566 7352 23572 7404
rect 23624 7392 23630 7404
rect 24213 7395 24271 7401
rect 24213 7392 24225 7395
rect 23624 7364 24225 7392
rect 23624 7352 23630 7364
rect 24213 7361 24225 7364
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 5040 7296 10824 7324
rect 5040 7284 5046 7296
rect 22462 7284 22468 7336
rect 22520 7284 22526 7336
rect 2222 7216 2228 7268
rect 2280 7216 2286 7268
rect 2869 7259 2927 7265
rect 2869 7225 2881 7259
rect 2915 7256 2927 7259
rect 8386 7256 8392 7268
rect 2915 7228 8392 7256
rect 2915 7225 2927 7228
rect 2869 7219 2927 7225
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 6362 7188 6368 7200
rect 3559 7160 6368 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 12434 7188 12440 7200
rect 10643 7160 12440 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 12529 7191 12587 7197
rect 12529 7157 12541 7191
rect 12575 7188 12587 7191
rect 13998 7188 14004 7200
rect 12575 7160 14004 7188
rect 12575 7157 12587 7160
rect 12529 7151 12587 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 17494 7188 17500 7200
rect 14139 7160 17500 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 3418 6944 3424 6996
rect 3476 6944 3482 6996
rect 23201 6987 23259 6993
rect 23201 6953 23213 6987
rect 23247 6984 23259 6987
rect 23934 6984 23940 6996
rect 23247 6956 23940 6984
rect 23247 6953 23259 6956
rect 23201 6947 23259 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 2869 6919 2927 6925
rect 2869 6885 2881 6919
rect 2915 6916 2927 6919
rect 2915 6888 4292 6916
rect 2915 6885 2927 6888
rect 2869 6879 2927 6885
rect 1302 6808 1308 6860
rect 1360 6848 1366 6860
rect 1360 6820 3096 6848
rect 1360 6808 1366 6820
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2590 6780 2596 6792
rect 2455 6752 2596 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3068 6789 3096 6820
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 3384 6820 4169 6848
rect 3384 6808 3390 6820
rect 4157 6817 4169 6820
rect 4203 6817 4215 6851
rect 4264 6848 4292 6888
rect 23750 6876 23756 6928
rect 23808 6876 23814 6928
rect 9766 6848 9772 6860
rect 4264 6820 9772 6848
rect 4157 6811 4215 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10560 6820 10609 6848
rect 10560 6808 10566 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 20714 6848 20720 6860
rect 19392 6820 20720 6848
rect 19392 6808 19398 6820
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 3053 6783 3111 6789
rect 2832 6752 2912 6780
rect 2832 6740 2838 6752
rect 2884 6712 2912 6752
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3099 6752 3525 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 21726 6740 21732 6792
rect 21784 6780 21790 6792
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 21784 6752 22937 6780
rect 21784 6740 21790 6752
rect 22925 6749 22937 6752
rect 22971 6780 22983 6783
rect 23768 6780 23796 6876
rect 22971 6752 23796 6780
rect 22971 6749 22983 6752
rect 22925 6743 22983 6749
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 1596 6684 2774 6712
rect 2884 6684 3801 6712
rect 1596 6653 1624 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2225 6647 2283 6653
rect 2225 6644 2237 6647
rect 2188 6616 2237 6644
rect 2188 6604 2194 6616
rect 2225 6613 2237 6616
rect 2271 6613 2283 6647
rect 2746 6644 2774 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 7098 6712 7104 6724
rect 3789 6675 3847 6681
rect 3896 6684 7104 6712
rect 3896 6644 3924 6684
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 2746 6616 3924 6644
rect 2225 6607 2283 6613
rect 3970 6604 3976 6656
rect 4028 6604 4034 6656
rect 23382 6604 23388 6656
rect 23440 6604 23446 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 4338 6440 4344 6452
rect 2915 6412 4344 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 22830 6400 22836 6452
rect 22888 6400 22894 6452
rect 1762 6332 1768 6384
rect 1820 6372 1826 6384
rect 3970 6372 3976 6384
rect 1820 6344 3976 6372
rect 1820 6332 1826 6344
rect 3970 6332 3976 6344
rect 4028 6332 4034 6384
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2924 6276 3065 6304
rect 2924 6264 2930 6276
rect 3053 6273 3065 6276
rect 3099 6304 3111 6307
rect 3329 6307 3387 6313
rect 3329 6304 3341 6307
rect 3099 6276 3341 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3329 6273 3341 6276
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 22440 6307 22498 6313
rect 22440 6273 22452 6307
rect 22486 6304 22498 6307
rect 22848 6304 22876 6400
rect 22486 6276 22876 6304
rect 22486 6273 22498 6276
rect 22440 6267 22498 6273
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 1360 6208 1593 6236
rect 1360 6196 1366 6208
rect 1581 6205 1593 6208
rect 1627 6205 1639 6239
rect 1581 6199 1639 6205
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 12250 6236 12256 6248
rect 1903 6208 12256 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 22511 6103 22569 6109
rect 22511 6069 22523 6103
rect 22557 6100 22569 6103
rect 22738 6100 22744 6112
rect 22557 6072 22744 6100
rect 22557 6069 22569 6072
rect 22511 6063 22569 6069
rect 22738 6060 22744 6072
rect 22796 6060 22802 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 1302 5856 1308 5908
rect 1360 5896 1366 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 1360 5868 2697 5896
rect 1360 5856 1366 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 18923 5868 21005 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 20993 5865 21005 5868
rect 21039 5896 21051 5899
rect 22462 5896 22468 5908
rect 21039 5868 22468 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 7558 5788 7564 5840
rect 7616 5828 7622 5840
rect 12618 5828 12624 5840
rect 7616 5800 12624 5828
rect 7616 5788 7622 5800
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 21726 5788 21732 5840
rect 21784 5788 21790 5840
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 5994 5760 6000 5772
rect 1903 5732 6000 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 14056 5732 15577 5760
rect 14056 5720 14062 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 16908 5732 17141 5760
rect 16908 5720 16914 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5692 1639 5695
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 1627 5664 2881 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 12676 5664 15761 5692
rect 12676 5652 12682 5664
rect 15749 5661 15761 5664
rect 15795 5692 15807 5695
rect 15795 5664 17172 5692
rect 15795 5661 15807 5664
rect 15749 5655 15807 5661
rect 16209 5559 16267 5565
rect 16209 5525 16221 5559
rect 16255 5556 16267 5559
rect 17034 5556 17040 5568
rect 16255 5528 17040 5556
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 17144 5556 17172 5664
rect 18506 5652 18512 5704
rect 18564 5692 18570 5704
rect 19337 5695 19395 5701
rect 19337 5692 19349 5695
rect 18564 5664 19349 5692
rect 18564 5652 18570 5664
rect 19337 5661 19349 5664
rect 19383 5661 19395 5695
rect 19337 5655 19395 5661
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20312 5664 20913 5692
rect 20312 5652 20318 5664
rect 20901 5661 20913 5664
rect 20947 5692 20959 5695
rect 21744 5692 21772 5788
rect 22738 5720 22744 5772
rect 22796 5760 22802 5772
rect 24857 5763 24915 5769
rect 24857 5760 24869 5763
rect 22796 5732 24869 5760
rect 22796 5720 22802 5732
rect 24857 5729 24869 5732
rect 24903 5729 24915 5763
rect 24857 5723 24915 5729
rect 26973 5763 27031 5769
rect 26973 5729 26985 5763
rect 27019 5760 27031 5763
rect 28718 5760 28724 5772
rect 27019 5732 28724 5760
rect 27019 5729 27031 5732
rect 26973 5723 27031 5729
rect 28718 5720 28724 5732
rect 28776 5720 28782 5772
rect 28813 5763 28871 5769
rect 28813 5729 28825 5763
rect 28859 5760 28871 5763
rect 28902 5760 28908 5772
rect 28859 5732 28908 5760
rect 28859 5729 28871 5732
rect 28813 5723 28871 5729
rect 28902 5720 28908 5732
rect 28960 5720 28966 5772
rect 20947 5664 21772 5692
rect 24673 5695 24731 5701
rect 20947 5661 20959 5664
rect 20901 5655 20959 5661
rect 24673 5661 24685 5695
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 17402 5584 17408 5636
rect 17460 5584 17466 5636
rect 22186 5624 22192 5636
rect 18708 5596 22192 5624
rect 18708 5556 18736 5596
rect 22186 5584 22192 5596
rect 22244 5624 22250 5636
rect 23382 5624 23388 5636
rect 22244 5596 23388 5624
rect 22244 5584 22250 5596
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 24688 5624 24716 5655
rect 25498 5624 25504 5636
rect 24688 5596 25504 5624
rect 25498 5584 25504 5596
rect 25556 5584 25562 5636
rect 26513 5627 26571 5633
rect 26513 5593 26525 5627
rect 26559 5593 26571 5627
rect 26513 5587 26571 5593
rect 17144 5528 18736 5556
rect 21358 5516 21364 5568
rect 21416 5516 21422 5568
rect 26528 5556 26556 5587
rect 27154 5584 27160 5636
rect 27212 5584 27218 5636
rect 27614 5556 27620 5568
rect 26528 5528 27620 5556
rect 27614 5516 27620 5528
rect 27672 5516 27678 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 22879 5355 22937 5361
rect 22879 5321 22891 5355
rect 22925 5352 22937 5355
rect 27154 5352 27160 5364
rect 22925 5324 27160 5352
rect 22925 5321 22937 5324
rect 22879 5315 22937 5321
rect 27154 5312 27160 5324
rect 27212 5312 27218 5364
rect 28350 5244 28356 5296
rect 28408 5284 28414 5296
rect 28408 5256 30052 5284
rect 28408 5244 28414 5256
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1360 5188 1593 5216
rect 1360 5176 1366 5188
rect 1581 5185 1593 5188
rect 1627 5216 1639 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 1627 5188 2697 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 12492 5188 15669 5216
rect 12492 5176 12498 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 21358 5216 21364 5228
rect 17604 5188 21364 5216
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 9398 5148 9404 5160
rect 1903 5120 9404 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15528 5120 15853 5148
rect 15528 5108 15534 5120
rect 15841 5117 15853 5120
rect 15887 5148 15899 5151
rect 17604 5148 17632 5188
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 22186 5225 22192 5228
rect 22164 5219 22192 5225
rect 22164 5185 22176 5219
rect 22164 5179 22192 5185
rect 22186 5176 22192 5179
rect 22244 5176 22250 5228
rect 22776 5219 22834 5225
rect 22776 5216 22788 5219
rect 22388 5188 22788 5216
rect 15887 5120 17632 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 17678 5108 17684 5160
rect 17736 5108 17742 5160
rect 21376 5148 21404 5176
rect 22388 5148 22416 5188
rect 22776 5185 22788 5188
rect 22822 5185 22834 5219
rect 22776 5179 22834 5185
rect 21376 5120 22416 5148
rect 28629 5151 28687 5157
rect 28629 5117 28641 5151
rect 28675 5117 28687 5151
rect 28629 5111 28687 5117
rect 28644 5080 28672 5111
rect 28810 5108 28816 5160
rect 28868 5108 28874 5160
rect 30024 5157 30052 5256
rect 30009 5151 30067 5157
rect 30009 5117 30021 5151
rect 30055 5148 30067 5151
rect 41414 5148 41420 5160
rect 30055 5120 41420 5148
rect 30055 5117 30067 5120
rect 30009 5111 30067 5117
rect 41414 5108 41420 5120
rect 41472 5108 41478 5160
rect 33502 5080 33508 5092
rect 28644 5052 33508 5080
rect 33502 5040 33508 5052
rect 33560 5040 33566 5092
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 17862 5012 17868 5024
rect 16347 4984 17868 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 20530 5012 20536 5024
rect 18187 4984 20536 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 22235 5015 22293 5021
rect 22235 4981 22247 5015
rect 22281 5012 22293 5015
rect 25958 5012 25964 5024
rect 22281 4984 25964 5012
rect 22281 4981 22293 4984
rect 22235 4975 22293 4981
rect 25958 4972 25964 4984
rect 26016 4972 26022 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 17460 4780 19533 4808
rect 17460 4768 17466 4780
rect 19521 4777 19533 4780
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 20254 4768 20260 4820
rect 20312 4768 20318 4820
rect 24719 4811 24777 4817
rect 24719 4777 24731 4811
rect 24765 4808 24777 4811
rect 28810 4808 28816 4820
rect 24765 4780 28816 4808
rect 24765 4777 24777 4780
rect 24719 4771 24777 4777
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 1581 4675 1639 4681
rect 1581 4672 1593 4675
rect 1360 4644 1593 4672
rect 1360 4632 1366 4644
rect 1581 4641 1593 4644
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 9950 4672 9956 4684
rect 1903 4644 9956 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 1596 4604 1624 4635
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 25777 4675 25835 4681
rect 25777 4641 25789 4675
rect 25823 4672 25835 4675
rect 27798 4672 27804 4684
rect 25823 4644 27804 4672
rect 25823 4641 25835 4644
rect 25777 4635 25835 4641
rect 27798 4632 27804 4644
rect 27856 4632 27862 4684
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 1596 4576 2881 4604
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20254 4604 20260 4616
rect 19475 4576 20260 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 22066 4576 24628 4604
rect 2774 4428 2780 4480
rect 2832 4428 2838 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 19889 4471 19947 4477
rect 19889 4468 19901 4471
rect 17736 4440 19901 4468
rect 17736 4428 17742 4440
rect 19889 4437 19901 4440
rect 19935 4468 19947 4471
rect 22066 4468 22094 4576
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 27246 4564 27252 4616
rect 27304 4604 27310 4616
rect 27617 4607 27675 4613
rect 27617 4604 27629 4607
rect 27304 4576 27629 4604
rect 27304 4564 27310 4576
rect 27617 4573 27629 4576
rect 27663 4573 27675 4607
rect 27617 4567 27675 4573
rect 25958 4496 25964 4548
rect 26016 4496 26022 4548
rect 19935 4440 22094 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 2271 4236 2774 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 2746 4196 2774 4236
rect 1688 4168 1900 4196
rect 2746 4168 3464 4196
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 1688 4128 1716 4168
rect 1268 4100 1716 4128
rect 1268 4088 1274 4100
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 1872 4128 1900 4168
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 1872 4100 2421 4128
rect 2409 4097 2421 4100
rect 2455 4128 2467 4131
rect 2774 4128 2780 4140
rect 2455 4100 2780 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3099 4100 3341 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3436 4128 3464 4168
rect 6822 4128 6828 4140
rect 3436 4100 6828 4128
rect 3329 4091 3387 4097
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 3068 4060 3096 4091
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 1360 4032 3096 4060
rect 1360 4020 1366 4032
rect 3513 3995 3571 4001
rect 3513 3992 3525 3995
rect 2746 3964 3525 3992
rect 1578 3884 1584 3936
rect 1636 3884 1642 3936
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 2746 3924 2774 3964
rect 3513 3961 3525 3964
rect 3559 3961 3571 3995
rect 3513 3955 3571 3961
rect 1820 3896 2774 3924
rect 2869 3927 2927 3933
rect 1820 3884 1826 3896
rect 2869 3893 2881 3927
rect 2915 3924 2927 3927
rect 10594 3924 10600 3936
rect 2915 3896 10600 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 15010 3884 15016 3936
rect 15068 3884 15074 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 1578 3680 1584 3732
rect 1636 3720 1642 3732
rect 9674 3720 9680 3732
rect 1636 3692 9680 3720
rect 1636 3680 1642 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 12066 3680 12072 3732
rect 12124 3680 12130 3732
rect 3513 3655 3571 3661
rect 3513 3652 3525 3655
rect 1596 3624 3525 3652
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1596 3525 1624 3624
rect 3513 3621 3525 3624
rect 3559 3621 3571 3655
rect 3513 3615 3571 3621
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 44082 3652 44088 3664
rect 28960 3624 44088 3652
rect 28960 3612 28966 3624
rect 44082 3612 44088 3624
rect 44140 3612 44146 3664
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 2038 3584 2044 3596
rect 1903 3556 2044 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 27246 3544 27252 3596
rect 27304 3584 27310 3596
rect 46750 3584 46756 3596
rect 27304 3556 46756 3584
rect 27304 3544 27310 3556
rect 46750 3544 46756 3556
rect 46808 3544 46814 3596
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2924 3488 3065 3516
rect 2924 3476 2930 3488
rect 3053 3485 3065 3488
rect 3099 3516 3111 3519
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3099 3488 3341 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 11256 3488 12434 3516
rect 11256 3448 11284 3488
rect 2884 3420 11284 3448
rect 11517 3451 11575 3457
rect 2884 3389 2912 3420
rect 11517 3417 11529 3451
rect 11563 3448 11575 3451
rect 12066 3448 12072 3460
rect 11563 3420 12072 3448
rect 11563 3417 11575 3420
rect 11517 3411 11575 3417
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12406 3448 12434 3488
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 49418 3516 49424 3528
rect 27672 3488 49424 3516
rect 27672 3476 27678 3488
rect 49418 3476 49424 3488
rect 49476 3476 49482 3528
rect 13446 3448 13452 3460
rect 12406 3420 13452 3448
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 20714 3408 20720 3460
rect 20772 3448 20778 3460
rect 38746 3448 38752 3460
rect 20772 3420 38752 3448
rect 20772 3408 20778 3420
rect 38746 3408 38752 3420
rect 38804 3408 38810 3460
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3349 2927 3383
rect 2869 3343 2927 3349
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3476 3352 3801 3380
rect 3476 3340 3482 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 3789 3343 3847 3349
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 9824 3148 14013 3176
rect 9824 3136 9830 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 14001 3139 14059 3145
rect 10410 3108 10416 3120
rect 10258 3080 10416 3108
rect 10410 3068 10416 3080
rect 10468 3108 10474 3120
rect 10781 3111 10839 3117
rect 10781 3108 10793 3111
rect 10468 3080 10793 3108
rect 10468 3068 10474 3080
rect 10781 3077 10793 3080
rect 10827 3077 10839 3111
rect 10781 3071 10839 3077
rect 12618 3068 12624 3120
rect 12676 3068 12682 3120
rect 13909 3111 13967 3117
rect 13909 3077 13921 3111
rect 13955 3108 13967 3111
rect 15470 3108 15476 3120
rect 13955 3080 15476 3108
rect 13955 3077 13967 3080
rect 13909 3071 13967 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15565 3111 15623 3117
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 17678 3108 17684 3120
rect 15611 3080 17684 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 1452 3012 2881 3040
rect 1452 3000 1458 3012
rect 2869 3009 2881 3012
rect 2915 3040 2927 3043
rect 3326 3040 3332 3052
rect 2915 3012 3332 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3559 3012 4169 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1360 2944 1593 2972
rect 1360 2932 1366 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2406 2972 2412 2984
rect 1903 2944 2412 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 1596 2904 1624 2935
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 6564 2972 6592 3003
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7892 3012 8769 3040
rect 7892 3000 7898 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17920 3012 18337 3040
rect 17920 3000 17926 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20530 3000 20536 3052
rect 20588 3000 20594 3052
rect 3988 2944 6592 2972
rect 7193 2975 7251 2981
rect 3786 2904 3792 2916
rect 1596 2876 3792 2904
rect 3786 2864 3792 2876
rect 3844 2864 3850 2916
rect 3988 2913 4016 2944
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 7239 2944 9045 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 17402 2972 17408 2984
rect 10551 2944 17408 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 3973 2907 4031 2913
rect 3973 2873 3985 2907
rect 4019 2873 4031 2907
rect 3973 2867 4031 2873
rect 10060 2876 10916 2904
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 10060 2836 10088 2876
rect 8352 2808 10088 2836
rect 10888 2836 10916 2876
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 12492 2876 15761 2904
rect 12492 2864 12498 2876
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 12713 2839 12771 2845
rect 12713 2836 12725 2839
rect 10888 2808 12725 2836
rect 8352 2796 8358 2808
rect 12713 2805 12725 2808
rect 12759 2805 12771 2839
rect 12713 2799 12771 2805
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17494 2836 17500 2848
rect 16899 2808 17500 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 20070 2836 20076 2848
rect 18187 2808 20076 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20349 2839 20407 2845
rect 20349 2805 20361 2839
rect 20395 2836 20407 2839
rect 22002 2836 22008 2848
rect 20395 2808 22008 2836
rect 20395 2805 20407 2808
rect 20349 2799 20407 2805
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 3326 2592 3332 2644
rect 3384 2592 3390 2644
rect 3786 2592 3792 2644
rect 3844 2592 3850 2644
rect 7558 2632 7564 2644
rect 4908 2604 7564 2632
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 4908 2564 4936 2604
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 25498 2592 25504 2644
rect 25556 2592 25562 2644
rect 27798 2592 27804 2644
rect 27856 2632 27862 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 27856 2604 28181 2632
rect 27856 2592 27862 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 28718 2592 28724 2644
rect 28776 2632 28782 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 28776 2604 30849 2632
rect 28776 2592 28782 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 33502 2592 33508 2644
rect 33560 2592 33566 2644
rect 11606 2564 11612 2576
rect 2915 2536 4936 2564
rect 5552 2536 11612 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1268 2468 1593 2496
rect 1268 2456 1274 2468
rect 1581 2465 1593 2468
rect 1627 2496 1639 2499
rect 3418 2496 3424 2508
rect 1627 2468 3424 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4120 2468 4629 2496
rect 4120 2456 4126 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 5552 2428 5580 2536
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6788 2468 7297 2496
rect 6788 2456 6794 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9456 2468 9965 2496
rect 9456 2456 9462 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12124 2468 12633 2496
rect 12124 2456 12130 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 14792 2468 15301 2496
rect 14792 2456 14798 2468
rect 15289 2465 15301 2468
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17957 2499 18015 2505
rect 17957 2496 17969 2499
rect 17460 2468 17969 2496
rect 17460 2456 17466 2468
rect 17957 2465 17969 2468
rect 18003 2465 18015 2499
rect 17957 2459 18015 2465
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22796 2468 23121 2496
rect 22796 2456 22802 2468
rect 23109 2465 23121 2468
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 31570 2456 31576 2508
rect 31628 2496 31634 2508
rect 36357 2499 36415 2505
rect 36357 2496 36369 2499
rect 31628 2468 36369 2496
rect 31628 2456 31634 2468
rect 36357 2465 36369 2468
rect 36403 2465 36415 2499
rect 36357 2459 36415 2465
rect 4387 2400 5580 2428
rect 7009 2431 7067 2437
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8294 2428 8300 2440
rect 7055 2400 8300 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 3068 2360 3096 2391
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12434 2428 12440 2440
rect 12391 2400 12440 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 15010 2388 15016 2440
rect 15068 2388 15074 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22060 2400 22661 2428
rect 22060 2388 22066 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25464 2400 25697 2428
rect 25464 2388 25470 2400
rect 25685 2397 25697 2400
rect 25731 2428 25743 2431
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25731 2400 25973 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33468 2400 33701 2428
rect 33468 2388 33474 2400
rect 33689 2397 33701 2400
rect 33735 2428 33747 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33735 2400 33977 2428
rect 33735 2397 33747 2400
rect 33689 2391 33747 2397
rect 33965 2397 33977 2400
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36136 2400 37289 2428
rect 36136 2388 36142 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 3513 2363 3571 2369
rect 3513 2360 3525 2363
rect 1360 2332 3525 2360
rect 1360 2320 1366 2332
rect 3513 2329 3525 2332
rect 3559 2329 3571 2363
rect 3513 2323 3571 2329
rect 1811 2295 1869 2301
rect 1811 2261 1823 2295
rect 1857 2292 1869 2295
rect 6546 2292 6552 2304
rect 1857 2264 6552 2292
rect 1857 2261 1869 2264
rect 1811 2255 1869 2261
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 8300 26324 8352 26376
rect 23388 26324 23440 26376
rect 12072 25712 12124 25764
rect 33968 25712 34020 25764
rect 10600 25644 10652 25696
rect 26884 25644 26936 25696
rect 13728 25576 13780 25628
rect 34888 25576 34940 25628
rect 10048 25508 10100 25560
rect 33600 25508 33652 25560
rect 10784 25440 10836 25492
rect 34980 25440 35032 25492
rect 14648 25372 14700 25424
rect 31116 25372 31168 25424
rect 12256 25304 12308 25356
rect 32312 25304 32364 25356
rect 13912 25236 13964 25288
rect 32496 25236 32548 25288
rect 4068 25168 4120 25220
rect 9128 25168 9180 25220
rect 10416 25168 10468 25220
rect 30196 25168 30248 25220
rect 16672 25100 16724 25152
rect 28540 25100 28592 25152
rect 15660 25032 15712 25084
rect 30380 25032 30432 25084
rect 15936 24964 15988 25016
rect 32864 24964 32916 25016
rect 15200 24896 15252 24948
rect 14740 24828 14792 24880
rect 21548 24828 21600 24880
rect 21916 24896 21968 24948
rect 39304 24896 39356 24948
rect 33508 24828 33560 24880
rect 6552 24760 6604 24812
rect 13544 24760 13596 24812
rect 14280 24760 14332 24812
rect 26148 24760 26200 24812
rect 26240 24760 26292 24812
rect 29184 24760 29236 24812
rect 3792 24692 3844 24744
rect 12624 24692 12676 24744
rect 13728 24692 13780 24744
rect 19064 24692 19116 24744
rect 26424 24692 26476 24744
rect 27252 24692 27304 24744
rect 4068 24624 4120 24676
rect 7288 24624 7340 24676
rect 12348 24624 12400 24676
rect 25780 24624 25832 24676
rect 26056 24624 26108 24676
rect 30472 24624 30524 24676
rect 31300 24692 31352 24744
rect 36636 24692 36688 24744
rect 31668 24624 31720 24676
rect 11704 24556 11756 24608
rect 21732 24556 21784 24608
rect 21916 24556 21968 24608
rect 30012 24556 30064 24608
rect 30380 24556 30432 24608
rect 34152 24556 34204 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 2780 24352 2832 24404
rect 4896 24352 4948 24404
rect 6552 24395 6604 24404
rect 6552 24361 6561 24395
rect 6561 24361 6595 24395
rect 6595 24361 6604 24395
rect 6552 24352 6604 24361
rect 11060 24352 11112 24404
rect 11704 24395 11756 24404
rect 11704 24361 11713 24395
rect 11713 24361 11747 24395
rect 11747 24361 11756 24395
rect 11704 24352 11756 24361
rect 14280 24395 14332 24404
rect 14280 24361 14289 24395
rect 14289 24361 14323 24395
rect 14323 24361 14332 24395
rect 14280 24352 14332 24361
rect 11980 24284 12032 24336
rect 3516 24216 3568 24268
rect 2412 24148 2464 24200
rect 3424 24148 3476 24200
rect 4252 24148 4304 24200
rect 1768 24080 1820 24132
rect 3700 24012 3752 24064
rect 6828 24216 6880 24268
rect 9220 24216 9272 24268
rect 14464 24284 14516 24336
rect 8392 24148 8444 24200
rect 8300 24080 8352 24132
rect 9220 24012 9272 24064
rect 10600 24148 10652 24200
rect 12624 24148 12676 24200
rect 18972 24352 19024 24404
rect 18420 24284 18472 24336
rect 25136 24352 25188 24404
rect 25780 24395 25832 24404
rect 25780 24361 25789 24395
rect 25789 24361 25823 24395
rect 25823 24361 25832 24395
rect 25780 24352 25832 24361
rect 27160 24395 27212 24404
rect 27160 24361 27169 24395
rect 27169 24361 27203 24395
rect 27203 24361 27212 24395
rect 27160 24352 27212 24361
rect 29092 24352 29144 24404
rect 18696 24216 18748 24268
rect 18972 24259 19024 24268
rect 18972 24225 18981 24259
rect 18981 24225 19015 24259
rect 19015 24225 19024 24259
rect 18972 24216 19024 24225
rect 19248 24216 19300 24268
rect 19892 24216 19944 24268
rect 20812 24216 20864 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 22100 24216 22152 24268
rect 27620 24284 27672 24336
rect 25228 24216 25280 24268
rect 26424 24216 26476 24268
rect 31576 24352 31628 24404
rect 31668 24352 31720 24404
rect 34152 24395 34204 24404
rect 34152 24361 34161 24395
rect 34161 24361 34195 24395
rect 34195 24361 34204 24395
rect 34152 24352 34204 24361
rect 13820 24080 13872 24132
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 15384 24148 15436 24200
rect 19984 24148 20036 24200
rect 15844 24080 15896 24132
rect 17132 24123 17184 24132
rect 17132 24089 17141 24123
rect 17141 24089 17175 24123
rect 17175 24089 17184 24123
rect 17132 24080 17184 24089
rect 17592 24080 17644 24132
rect 19340 24080 19392 24132
rect 21732 24148 21784 24200
rect 23940 24148 23992 24200
rect 24952 24148 25004 24200
rect 26056 24148 26108 24200
rect 26148 24148 26200 24200
rect 29276 24216 29328 24268
rect 30012 24259 30064 24268
rect 30012 24225 30021 24259
rect 30021 24225 30055 24259
rect 30055 24225 30064 24259
rect 30012 24216 30064 24225
rect 30656 24284 30708 24336
rect 33876 24284 33928 24336
rect 34060 24284 34112 24336
rect 39304 24395 39356 24404
rect 39304 24361 39313 24395
rect 39313 24361 39347 24395
rect 39347 24361 39356 24395
rect 39304 24352 39356 24361
rect 44732 24395 44784 24404
rect 44732 24361 44741 24395
rect 44741 24361 44775 24395
rect 44775 24361 44784 24395
rect 44732 24352 44784 24361
rect 35900 24327 35952 24336
rect 35900 24293 35909 24327
rect 35909 24293 35943 24327
rect 35943 24293 35952 24327
rect 35900 24284 35952 24293
rect 36912 24284 36964 24336
rect 39580 24216 39632 24268
rect 40132 24216 40184 24268
rect 16764 24012 16816 24064
rect 17408 24012 17460 24064
rect 20444 24012 20496 24064
rect 27712 24080 27764 24132
rect 24032 24012 24084 24064
rect 24952 24055 25004 24064
rect 24952 24021 24961 24055
rect 24961 24021 24995 24055
rect 24995 24021 25004 24055
rect 24952 24012 25004 24021
rect 26056 24012 26108 24064
rect 26976 24012 27028 24064
rect 29184 24191 29236 24200
rect 29184 24157 29193 24191
rect 29193 24157 29227 24191
rect 29227 24157 29236 24191
rect 29184 24148 29236 24157
rect 29920 24148 29972 24200
rect 30564 24148 30616 24200
rect 31852 24148 31904 24200
rect 32680 24148 32732 24200
rect 33324 24191 33376 24200
rect 33324 24157 33333 24191
rect 33333 24157 33367 24191
rect 33367 24157 33376 24191
rect 33324 24148 33376 24157
rect 34060 24191 34112 24200
rect 34060 24157 34069 24191
rect 34069 24157 34103 24191
rect 34103 24157 34112 24191
rect 34060 24148 34112 24157
rect 34520 24148 34572 24200
rect 35624 24148 35676 24200
rect 35900 24148 35952 24200
rect 36820 24148 36872 24200
rect 37280 24148 37332 24200
rect 38476 24191 38528 24200
rect 38476 24157 38485 24191
rect 38485 24157 38519 24191
rect 38519 24157 38528 24191
rect 38476 24148 38528 24157
rect 38660 24191 38712 24200
rect 38660 24157 38669 24191
rect 38669 24157 38703 24191
rect 38703 24157 38712 24191
rect 38660 24148 38712 24157
rect 39212 24191 39264 24200
rect 39212 24157 39221 24191
rect 39221 24157 39255 24191
rect 39255 24157 39264 24191
rect 39212 24148 39264 24157
rect 41512 24148 41564 24200
rect 43260 24148 43312 24200
rect 44732 24148 44784 24200
rect 45560 24148 45612 24200
rect 46020 24148 46072 24200
rect 47308 24148 47360 24200
rect 48596 24191 48648 24200
rect 48596 24157 48605 24191
rect 48605 24157 48639 24191
rect 48639 24157 48648 24191
rect 48596 24148 48648 24157
rect 28356 24055 28408 24064
rect 28356 24021 28365 24055
rect 28365 24021 28399 24055
rect 28399 24021 28408 24055
rect 28356 24012 28408 24021
rect 29092 24012 29144 24064
rect 31576 24080 31628 24132
rect 31668 24080 31720 24132
rect 35164 24080 35216 24132
rect 36268 24080 36320 24132
rect 36636 24080 36688 24132
rect 31852 24055 31904 24064
rect 31852 24021 31861 24055
rect 31861 24021 31895 24055
rect 31895 24021 31904 24055
rect 31852 24012 31904 24021
rect 33416 24055 33468 24064
rect 33416 24021 33425 24055
rect 33425 24021 33459 24055
rect 33459 24021 33468 24055
rect 33416 24012 33468 24021
rect 35072 24055 35124 24064
rect 35072 24021 35081 24055
rect 35081 24021 35115 24055
rect 35115 24021 35124 24055
rect 35072 24012 35124 24021
rect 35256 24012 35308 24064
rect 36452 24012 36504 24064
rect 42064 24055 42116 24064
rect 42064 24021 42073 24055
rect 42073 24021 42107 24055
rect 42107 24021 42116 24055
rect 42064 24012 42116 24021
rect 42616 24055 42668 24064
rect 42616 24021 42625 24055
rect 42625 24021 42659 24055
rect 42659 24021 42668 24055
rect 42616 24012 42668 24021
rect 45376 24055 45428 24064
rect 45376 24021 45385 24055
rect 45385 24021 45419 24055
rect 45419 24021 45428 24055
rect 45376 24012 45428 24021
rect 46848 24055 46900 24064
rect 46848 24021 46857 24055
rect 46857 24021 46891 24055
rect 46891 24021 46900 24055
rect 46848 24012 46900 24021
rect 47032 24012 47084 24064
rect 48688 24012 48740 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 3424 23808 3476 23860
rect 6000 23808 6052 23860
rect 6644 23808 6696 23860
rect 12256 23851 12308 23860
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 12348 23851 12400 23860
rect 12348 23817 12357 23851
rect 12357 23817 12391 23851
rect 12391 23817 12400 23851
rect 12348 23808 12400 23817
rect 12440 23808 12492 23860
rect 21916 23808 21968 23860
rect 4068 23740 4120 23792
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 3516 23672 3568 23724
rect 4068 23604 4120 23656
rect 8576 23740 8628 23792
rect 9956 23740 10008 23792
rect 12532 23740 12584 23792
rect 15752 23740 15804 23792
rect 18328 23740 18380 23792
rect 19064 23740 19116 23792
rect 19248 23740 19300 23792
rect 21180 23783 21232 23792
rect 21180 23749 21189 23783
rect 21189 23749 21223 23783
rect 21223 23749 21232 23783
rect 21180 23740 21232 23749
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 6552 23672 6604 23724
rect 7748 23672 7800 23724
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 11152 23672 11204 23724
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 16580 23672 16632 23724
rect 16948 23715 17000 23724
rect 16948 23681 16957 23715
rect 16957 23681 16991 23715
rect 16991 23681 17000 23715
rect 16948 23672 17000 23681
rect 17132 23672 17184 23724
rect 18420 23672 18472 23724
rect 18696 23715 18748 23724
rect 18696 23681 18705 23715
rect 18705 23681 18739 23715
rect 18739 23681 18748 23715
rect 18696 23672 18748 23681
rect 20720 23672 20772 23724
rect 21824 23672 21876 23724
rect 23848 23808 23900 23860
rect 24952 23808 25004 23860
rect 25780 23808 25832 23860
rect 30196 23851 30248 23860
rect 30196 23817 30205 23851
rect 30205 23817 30239 23851
rect 30239 23817 30248 23851
rect 30196 23808 30248 23817
rect 31024 23808 31076 23860
rect 38476 23851 38528 23860
rect 38476 23817 38485 23851
rect 38485 23817 38519 23851
rect 38519 23817 38528 23851
rect 38476 23808 38528 23817
rect 39212 23808 39264 23860
rect 39580 23808 39632 23860
rect 40316 23851 40368 23860
rect 40316 23817 40325 23851
rect 40325 23817 40359 23851
rect 40359 23817 40368 23851
rect 40316 23808 40368 23817
rect 41512 23808 41564 23860
rect 43260 23851 43312 23860
rect 43260 23817 43269 23851
rect 43269 23817 43303 23851
rect 43303 23817 43312 23851
rect 43260 23808 43312 23817
rect 45560 23808 45612 23860
rect 47308 23808 47360 23860
rect 47860 23851 47912 23860
rect 47860 23817 47869 23851
rect 47869 23817 47903 23851
rect 47903 23817 47912 23851
rect 47860 23808 47912 23817
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 1216 23536 1268 23588
rect 1768 23468 1820 23520
rect 7380 23647 7432 23656
rect 7380 23613 7389 23647
rect 7389 23613 7423 23647
rect 7423 23613 7432 23647
rect 7380 23604 7432 23613
rect 7472 23604 7524 23656
rect 11336 23536 11388 23588
rect 17408 23604 17460 23656
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 16764 23536 16816 23588
rect 17592 23536 17644 23588
rect 22376 23604 22428 23656
rect 25412 23740 25464 23792
rect 26424 23740 26476 23792
rect 30104 23783 30156 23792
rect 30104 23749 30113 23783
rect 30113 23749 30147 23783
rect 30147 23749 30156 23783
rect 30104 23740 30156 23749
rect 32312 23783 32364 23792
rect 32312 23749 32321 23783
rect 32321 23749 32355 23783
rect 32355 23749 32364 23783
rect 32312 23740 32364 23749
rect 32864 23740 32916 23792
rect 33600 23740 33652 23792
rect 34888 23783 34940 23792
rect 34888 23749 34897 23783
rect 34897 23749 34931 23783
rect 34931 23749 34940 23783
rect 34888 23740 34940 23749
rect 34980 23740 35032 23792
rect 36544 23740 36596 23792
rect 28540 23672 28592 23724
rect 3884 23468 3936 23520
rect 4988 23468 5040 23520
rect 6552 23511 6604 23520
rect 6552 23477 6561 23511
rect 6561 23477 6595 23511
rect 6595 23477 6604 23511
rect 6552 23468 6604 23477
rect 11428 23468 11480 23520
rect 12256 23468 12308 23520
rect 12808 23468 12860 23520
rect 18696 23468 18748 23520
rect 20076 23468 20128 23520
rect 20628 23468 20680 23520
rect 22100 23468 22152 23520
rect 22836 23468 22888 23520
rect 23756 23511 23808 23520
rect 23756 23477 23765 23511
rect 23765 23477 23799 23511
rect 23799 23477 23808 23511
rect 23756 23468 23808 23477
rect 26148 23604 26200 23656
rect 27160 23647 27212 23656
rect 27160 23613 27169 23647
rect 27169 23613 27203 23647
rect 27203 23613 27212 23647
rect 27160 23604 27212 23613
rect 27528 23604 27580 23656
rect 30380 23672 30432 23724
rect 31392 23672 31444 23724
rect 32128 23604 32180 23656
rect 34704 23715 34756 23724
rect 34704 23681 34713 23715
rect 34713 23681 34747 23715
rect 34747 23681 34756 23715
rect 34704 23672 34756 23681
rect 36268 23715 36320 23724
rect 36268 23681 36277 23715
rect 36277 23681 36311 23715
rect 36311 23681 36320 23715
rect 36268 23672 36320 23681
rect 36360 23672 36412 23724
rect 37648 23672 37700 23724
rect 40960 23672 41012 23724
rect 42064 23672 42116 23724
rect 43720 23715 43772 23724
rect 43720 23681 43729 23715
rect 43729 23681 43763 23715
rect 43763 23681 43772 23715
rect 43720 23672 43772 23681
rect 44180 23672 44232 23724
rect 46664 23672 46716 23724
rect 48320 23715 48372 23724
rect 48320 23681 48329 23715
rect 48329 23681 48363 23715
rect 48363 23681 48372 23715
rect 48320 23672 48372 23681
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 26792 23468 26844 23520
rect 30656 23536 30708 23588
rect 30748 23536 30800 23588
rect 31668 23536 31720 23588
rect 31760 23579 31812 23588
rect 31760 23545 31769 23579
rect 31769 23545 31803 23579
rect 31803 23545 31812 23579
rect 31760 23536 31812 23545
rect 32588 23536 32640 23588
rect 28724 23468 28776 23520
rect 30564 23511 30616 23520
rect 30564 23477 30573 23511
rect 30573 23477 30607 23511
rect 30607 23477 30616 23511
rect 30564 23468 30616 23477
rect 31116 23468 31168 23520
rect 33876 23468 33928 23520
rect 37188 23536 37240 23588
rect 36728 23511 36780 23520
rect 36728 23477 36737 23511
rect 36737 23477 36771 23511
rect 36771 23477 36780 23511
rect 36728 23468 36780 23477
rect 37740 23511 37792 23520
rect 37740 23477 37749 23511
rect 37749 23477 37783 23511
rect 37783 23477 37792 23511
rect 37740 23468 37792 23477
rect 40776 23536 40828 23588
rect 41420 23468 41472 23520
rect 44640 23511 44692 23520
rect 44640 23477 44649 23511
rect 44649 23477 44683 23511
rect 44683 23477 44692 23511
rect 44640 23468 44692 23477
rect 46940 23511 46992 23520
rect 46940 23477 46949 23511
rect 46949 23477 46983 23511
rect 46983 23477 46992 23511
rect 46940 23468 46992 23477
rect 48504 23511 48556 23520
rect 48504 23477 48513 23511
rect 48513 23477 48547 23511
rect 48547 23477 48556 23511
rect 48504 23468 48556 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 3700 23264 3752 23316
rect 3884 23264 3936 23316
rect 3976 23307 4028 23316
rect 3976 23273 3985 23307
rect 3985 23273 4019 23307
rect 4019 23273 4028 23307
rect 3976 23264 4028 23273
rect 3424 23196 3476 23248
rect 17960 23264 18012 23316
rect 24124 23264 24176 23316
rect 24400 23264 24452 23316
rect 26608 23264 26660 23316
rect 3792 23128 3844 23180
rect 6644 23196 6696 23248
rect 12808 23196 12860 23248
rect 19064 23196 19116 23248
rect 19432 23239 19484 23248
rect 19432 23205 19441 23239
rect 19441 23205 19475 23239
rect 19475 23205 19484 23239
rect 19432 23196 19484 23205
rect 19616 23196 19668 23248
rect 23756 23196 23808 23248
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 4712 23171 4764 23180
rect 4712 23137 4721 23171
rect 4721 23137 4755 23171
rect 4755 23137 4764 23171
rect 4712 23128 4764 23137
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 9036 23128 9088 23180
rect 4252 22992 4304 23044
rect 5172 22992 5224 23044
rect 5356 23103 5408 23112
rect 5356 23069 5365 23103
rect 5365 23069 5399 23103
rect 5399 23069 5408 23103
rect 5356 23060 5408 23069
rect 7196 23103 7248 23112
rect 7196 23069 7205 23103
rect 7205 23069 7239 23103
rect 7239 23069 7248 23103
rect 7196 23060 7248 23069
rect 8852 23060 8904 23112
rect 11428 23128 11480 23180
rect 12440 23128 12492 23180
rect 12532 23128 12584 23180
rect 17776 23128 17828 23180
rect 17868 23128 17920 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 26148 23196 26200 23248
rect 27068 23264 27120 23316
rect 27344 23264 27396 23316
rect 28724 23264 28776 23316
rect 29000 23307 29052 23316
rect 29000 23273 29009 23307
rect 29009 23273 29043 23307
rect 29043 23273 29052 23307
rect 29000 23264 29052 23273
rect 30564 23264 30616 23316
rect 31852 23307 31904 23316
rect 31852 23273 31861 23307
rect 31861 23273 31895 23307
rect 31895 23273 31904 23307
rect 31852 23264 31904 23273
rect 32312 23264 32364 23316
rect 32496 23307 32548 23316
rect 32496 23273 32505 23307
rect 32505 23273 32539 23307
rect 32539 23273 32548 23307
rect 32496 23264 32548 23273
rect 33508 23264 33560 23316
rect 33968 23307 34020 23316
rect 33968 23273 33977 23307
rect 33977 23273 34011 23307
rect 34011 23273 34020 23307
rect 33968 23264 34020 23273
rect 34428 23307 34480 23316
rect 34428 23273 34437 23307
rect 34437 23273 34471 23307
rect 34471 23273 34480 23307
rect 34428 23264 34480 23273
rect 16672 23060 16724 23112
rect 16856 23060 16908 23112
rect 7564 22992 7616 23044
rect 8484 22992 8536 23044
rect 4160 22967 4212 22976
rect 4160 22933 4169 22967
rect 4169 22933 4203 22967
rect 4203 22933 4212 22967
rect 4160 22924 4212 22933
rect 7472 22924 7524 22976
rect 9036 22967 9088 22976
rect 9036 22933 9045 22967
rect 9045 22933 9079 22967
rect 9079 22933 9088 22967
rect 9036 22924 9088 22933
rect 9588 23035 9640 23044
rect 9588 23001 9597 23035
rect 9597 23001 9631 23035
rect 9631 23001 9640 23035
rect 9588 22992 9640 23001
rect 12256 22992 12308 23044
rect 14372 23035 14424 23044
rect 14372 23001 14381 23035
rect 14381 23001 14415 23035
rect 14415 23001 14424 23035
rect 14372 22992 14424 23001
rect 11336 22924 11388 22976
rect 12532 22924 12584 22976
rect 12716 22924 12768 22976
rect 13544 22924 13596 22976
rect 17408 23035 17460 23044
rect 17408 23001 17417 23035
rect 17417 23001 17451 23035
rect 17451 23001 17460 23035
rect 17408 22992 17460 23001
rect 17500 22992 17552 23044
rect 17684 22924 17736 22976
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 35072 23196 35124 23248
rect 27160 23128 27212 23180
rect 27620 23128 27672 23180
rect 30748 23128 30800 23180
rect 36820 23307 36872 23316
rect 36820 23273 36829 23307
rect 36829 23273 36863 23307
rect 36863 23273 36872 23307
rect 36820 23264 36872 23273
rect 37280 23307 37332 23316
rect 37280 23273 37289 23307
rect 37289 23273 37323 23307
rect 37323 23273 37332 23307
rect 37280 23264 37332 23273
rect 43720 23264 43772 23316
rect 35624 23196 35676 23248
rect 28540 23060 28592 23112
rect 20352 23035 20404 23044
rect 20352 23001 20361 23035
rect 20361 23001 20395 23035
rect 20395 23001 20404 23035
rect 20352 22992 20404 23001
rect 22100 22992 22152 23044
rect 23848 22992 23900 23044
rect 24492 22992 24544 23044
rect 20536 22924 20588 22976
rect 21824 22967 21876 22976
rect 21824 22933 21833 22967
rect 21833 22933 21867 22967
rect 21867 22933 21876 22967
rect 21824 22924 21876 22933
rect 23204 22924 23256 22976
rect 24124 22924 24176 22976
rect 24952 22967 25004 22976
rect 24952 22933 24961 22967
rect 24961 22933 24995 22967
rect 24995 22933 25004 22967
rect 24952 22924 25004 22933
rect 25412 22924 25464 22976
rect 26056 22924 26108 22976
rect 26516 22924 26568 22976
rect 26792 22967 26844 22976
rect 26792 22933 26801 22967
rect 26801 22933 26835 22967
rect 26835 22933 26844 22967
rect 26792 22924 26844 22933
rect 28356 22924 28408 22976
rect 31852 23060 31904 23112
rect 28816 22992 28868 23044
rect 32036 23060 32088 23112
rect 34980 23060 35032 23112
rect 35716 23103 35768 23112
rect 35716 23069 35725 23103
rect 35725 23069 35759 23103
rect 35759 23069 35768 23103
rect 35716 23060 35768 23069
rect 28908 22924 28960 22976
rect 29184 22924 29236 22976
rect 32864 22992 32916 23044
rect 33324 22992 33376 23044
rect 31484 22967 31536 22976
rect 31484 22933 31493 22967
rect 31493 22933 31527 22967
rect 31527 22933 31536 22967
rect 31484 22924 31536 22933
rect 31944 22967 31996 22976
rect 31944 22933 31953 22967
rect 31953 22933 31987 22967
rect 31987 22933 31996 22967
rect 31944 22924 31996 22933
rect 32496 22924 32548 22976
rect 36268 22992 36320 23044
rect 42616 23060 42668 23112
rect 48688 23060 48740 23112
rect 49056 23103 49108 23112
rect 49056 23069 49065 23103
rect 49065 23069 49099 23103
rect 49099 23069 49108 23103
rect 49056 23060 49108 23069
rect 34888 22967 34940 22976
rect 34888 22933 34897 22967
rect 34897 22933 34931 22967
rect 34931 22933 34940 22967
rect 34888 22924 34940 22933
rect 35072 22924 35124 22976
rect 36176 22967 36228 22976
rect 36176 22933 36185 22967
rect 36185 22933 36219 22967
rect 36219 22933 36228 22967
rect 36176 22924 36228 22933
rect 39948 22924 40000 22976
rect 44548 22967 44600 22976
rect 44548 22933 44557 22967
rect 44557 22933 44591 22967
rect 44591 22933 44600 22967
rect 44548 22924 44600 22933
rect 47216 22924 47268 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 1032 22720 1084 22772
rect 5356 22720 5408 22772
rect 7564 22720 7616 22772
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 11888 22720 11940 22772
rect 12532 22720 12584 22772
rect 12624 22652 12676 22704
rect 12716 22695 12768 22704
rect 12716 22661 12725 22695
rect 12725 22661 12759 22695
rect 12759 22661 12768 22695
rect 12716 22652 12768 22661
rect 12808 22652 12860 22704
rect 18512 22720 18564 22772
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 16672 22652 16724 22704
rect 17684 22652 17736 22704
rect 3424 22584 3476 22636
rect 3792 22627 3844 22636
rect 3792 22593 3801 22627
rect 3801 22593 3835 22627
rect 3835 22593 3844 22627
rect 3792 22584 3844 22593
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 6644 22584 6696 22636
rect 7840 22584 7892 22636
rect 2872 22516 2924 22568
rect 2596 22380 2648 22432
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 7656 22516 7708 22568
rect 4620 22448 4672 22500
rect 7104 22448 7156 22500
rect 8208 22584 8260 22636
rect 10048 22584 10100 22636
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 9864 22516 9916 22568
rect 11704 22516 11756 22568
rect 12348 22584 12400 22636
rect 16764 22584 16816 22636
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 19432 22584 19484 22636
rect 20076 22652 20128 22704
rect 20352 22720 20404 22772
rect 25136 22720 25188 22772
rect 25780 22763 25832 22772
rect 25780 22729 25789 22763
rect 25789 22729 25823 22763
rect 25823 22729 25832 22763
rect 25780 22720 25832 22729
rect 23664 22652 23716 22704
rect 24676 22652 24728 22704
rect 28448 22720 28500 22772
rect 30380 22720 30432 22772
rect 30472 22720 30524 22772
rect 31668 22720 31720 22772
rect 34704 22720 34756 22772
rect 35072 22763 35124 22772
rect 35072 22729 35081 22763
rect 35081 22729 35115 22763
rect 35115 22729 35124 22763
rect 35072 22720 35124 22729
rect 27528 22695 27580 22704
rect 27528 22661 27537 22695
rect 27537 22661 27571 22695
rect 27571 22661 27580 22695
rect 27528 22652 27580 22661
rect 27620 22652 27672 22704
rect 22284 22584 22336 22636
rect 22836 22584 22888 22636
rect 24492 22584 24544 22636
rect 26792 22584 26844 22636
rect 27436 22584 27488 22636
rect 28908 22652 28960 22704
rect 29920 22652 29972 22704
rect 30932 22627 30984 22636
rect 30932 22593 30941 22627
rect 30941 22593 30975 22627
rect 30975 22593 30984 22627
rect 30932 22584 30984 22593
rect 31024 22627 31076 22636
rect 31024 22593 31033 22627
rect 31033 22593 31067 22627
rect 31067 22593 31076 22627
rect 31024 22584 31076 22593
rect 31760 22652 31812 22704
rect 44548 22720 44600 22772
rect 48596 22763 48648 22772
rect 48596 22729 48605 22763
rect 48605 22729 48639 22763
rect 48639 22729 48648 22763
rect 48596 22720 48648 22729
rect 31668 22584 31720 22636
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 32496 22584 32548 22636
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 16856 22559 16908 22568
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 16212 22448 16264 22500
rect 20628 22516 20680 22568
rect 18420 22448 18472 22500
rect 21548 22448 21600 22500
rect 22284 22448 22336 22500
rect 23112 22448 23164 22500
rect 23480 22516 23532 22568
rect 5264 22380 5316 22432
rect 6460 22423 6512 22432
rect 6460 22389 6469 22423
rect 6469 22389 6503 22423
rect 6503 22389 6512 22423
rect 6460 22380 6512 22389
rect 6736 22423 6788 22432
rect 6736 22389 6745 22423
rect 6745 22389 6779 22423
rect 6779 22389 6788 22423
rect 6736 22380 6788 22389
rect 6828 22380 6880 22432
rect 13452 22380 13504 22432
rect 17500 22380 17552 22432
rect 17684 22380 17736 22432
rect 18512 22380 18564 22432
rect 19156 22380 19208 22432
rect 19800 22380 19852 22432
rect 20168 22380 20220 22432
rect 22100 22380 22152 22432
rect 23848 22380 23900 22432
rect 23940 22380 23992 22432
rect 25688 22448 25740 22500
rect 25872 22559 25924 22568
rect 25872 22525 25881 22559
rect 25881 22525 25915 22559
rect 25915 22525 25924 22559
rect 25872 22516 25924 22525
rect 26424 22559 26476 22568
rect 26424 22525 26433 22559
rect 26433 22525 26467 22559
rect 26467 22525 26476 22559
rect 26424 22516 26476 22525
rect 26976 22516 27028 22568
rect 27252 22516 27304 22568
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 26516 22423 26568 22432
rect 26516 22389 26525 22423
rect 26525 22389 26559 22423
rect 26559 22389 26568 22423
rect 26516 22380 26568 22389
rect 27344 22448 27396 22500
rect 28724 22516 28776 22568
rect 31208 22516 31260 22568
rect 33600 22627 33652 22636
rect 33600 22593 33609 22627
rect 33609 22593 33643 22627
rect 33643 22593 33652 22627
rect 33600 22584 33652 22593
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 34980 22627 35032 22636
rect 34980 22593 34989 22627
rect 34989 22593 35023 22627
rect 35023 22593 35032 22627
rect 34980 22584 35032 22593
rect 39948 22695 40000 22704
rect 39948 22661 39957 22695
rect 39957 22661 39991 22695
rect 39991 22661 40000 22695
rect 39948 22652 40000 22661
rect 49240 22584 49292 22636
rect 28264 22380 28316 22432
rect 31484 22448 31536 22500
rect 30104 22423 30156 22432
rect 30104 22389 30113 22423
rect 30113 22389 30147 22423
rect 30147 22389 30156 22423
rect 30104 22380 30156 22389
rect 30932 22380 30984 22432
rect 32496 22423 32548 22432
rect 32496 22389 32505 22423
rect 32505 22389 32539 22423
rect 32539 22389 32548 22423
rect 32496 22380 32548 22389
rect 34428 22516 34480 22568
rect 34612 22516 34664 22568
rect 33416 22448 33468 22500
rect 35716 22380 35768 22432
rect 48320 22380 48372 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 6460 22176 6512 22228
rect 14188 22176 14240 22228
rect 3700 22108 3752 22160
rect 1308 22040 1360 22092
rect 3240 22040 3292 22092
rect 4252 22040 4304 22092
rect 4804 22108 4856 22160
rect 16120 22176 16172 22228
rect 16396 22176 16448 22228
rect 15108 22108 15160 22160
rect 6828 22040 6880 22092
rect 7012 22040 7064 22092
rect 2504 21904 2556 21956
rect 6552 21972 6604 22024
rect 7564 21972 7616 22024
rect 9864 22040 9916 22092
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 9772 22015 9824 22024
rect 9772 21981 9781 22015
rect 9781 21981 9815 22015
rect 9815 21981 9824 22015
rect 9772 21972 9824 21981
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 12624 22040 12676 22092
rect 10048 21972 10100 22024
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 10784 21972 10836 22024
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 13544 22040 13596 22092
rect 18512 22108 18564 22160
rect 20260 22176 20312 22228
rect 21272 22176 21324 22228
rect 23296 22176 23348 22228
rect 5816 21879 5868 21888
rect 5816 21845 5825 21879
rect 5825 21845 5859 21879
rect 5859 21845 5868 21879
rect 5816 21836 5868 21845
rect 6092 21879 6144 21888
rect 6092 21845 6101 21879
rect 6101 21845 6135 21879
rect 6135 21845 6144 21879
rect 6092 21836 6144 21845
rect 6920 21836 6972 21888
rect 8208 21836 8260 21888
rect 8668 21836 8720 21888
rect 9036 21836 9088 21888
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 13912 21904 13964 21956
rect 14648 21904 14700 21956
rect 19432 22040 19484 22092
rect 22008 22108 22060 22160
rect 23756 22108 23808 22160
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 18880 21972 18932 22024
rect 19616 21972 19668 22024
rect 21548 22040 21600 22092
rect 24400 22108 24452 22160
rect 26240 22176 26292 22228
rect 27344 22176 27396 22228
rect 28356 22176 28408 22228
rect 31852 22176 31904 22228
rect 32220 22176 32272 22228
rect 32864 22176 32916 22228
rect 29000 22108 29052 22160
rect 29184 22151 29236 22160
rect 29184 22117 29193 22151
rect 29193 22117 29227 22151
rect 29227 22117 29236 22151
rect 29184 22108 29236 22117
rect 30288 22108 30340 22160
rect 20260 21972 20312 22024
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 22192 21972 22244 22024
rect 23572 21972 23624 22024
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 24676 21972 24728 22024
rect 26700 22040 26752 22092
rect 26792 22040 26844 22092
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 27068 21972 27120 22024
rect 27344 21972 27396 22024
rect 28264 21972 28316 22024
rect 29828 22040 29880 22092
rect 30380 22040 30432 22092
rect 31484 22108 31536 22160
rect 31116 22040 31168 22092
rect 32680 22040 32732 22092
rect 17132 21904 17184 21956
rect 17408 21947 17460 21956
rect 17408 21913 17417 21947
rect 17417 21913 17451 21947
rect 17451 21913 17460 21947
rect 17408 21904 17460 21913
rect 17684 21904 17736 21956
rect 17868 21904 17920 21956
rect 11520 21836 11572 21888
rect 14096 21836 14148 21888
rect 14924 21879 14976 21888
rect 14924 21845 14933 21879
rect 14933 21845 14967 21879
rect 14967 21845 14976 21879
rect 19800 21904 19852 21956
rect 26332 21904 26384 21956
rect 29920 21904 29972 21956
rect 14924 21836 14976 21845
rect 18972 21836 19024 21888
rect 19064 21836 19116 21888
rect 22008 21836 22060 21888
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 23296 21879 23348 21888
rect 23296 21845 23305 21879
rect 23305 21845 23339 21879
rect 23339 21845 23348 21879
rect 23296 21836 23348 21845
rect 24308 21836 24360 21888
rect 25964 21836 26016 21888
rect 28448 21836 28500 21888
rect 29000 21836 29052 21888
rect 30472 22015 30524 22024
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 31208 21904 31260 21956
rect 32772 21972 32824 22024
rect 32864 22015 32916 22024
rect 32864 21981 32873 22015
rect 32873 21981 32907 22015
rect 32907 21981 32916 22015
rect 32864 21972 32916 21981
rect 33324 21972 33376 22024
rect 49056 22015 49108 22024
rect 49056 21981 49065 22015
rect 49065 21981 49099 22015
rect 49099 21981 49108 22015
rect 49056 21972 49108 21981
rect 35256 21904 35308 21956
rect 31668 21836 31720 21888
rect 32404 21836 32456 21888
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 5724 21632 5776 21684
rect 5816 21632 5868 21684
rect 3976 21564 4028 21616
rect 6184 21564 6236 21616
rect 6276 21564 6328 21616
rect 7380 21564 7432 21616
rect 8668 21564 8720 21616
rect 2228 21496 2280 21548
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 7012 21539 7064 21548
rect 7012 21505 7021 21539
rect 7021 21505 7055 21539
rect 7055 21505 7064 21539
rect 7012 21496 7064 21505
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 2780 21428 2832 21437
rect 3332 21428 3384 21480
rect 3424 21360 3476 21412
rect 5264 21428 5316 21480
rect 5356 21428 5408 21480
rect 5816 21471 5868 21480
rect 5816 21437 5825 21471
rect 5825 21437 5859 21471
rect 5859 21437 5868 21471
rect 5816 21428 5868 21437
rect 2136 21292 2188 21344
rect 6828 21360 6880 21412
rect 8944 21496 8996 21548
rect 9680 21632 9732 21684
rect 10968 21675 11020 21684
rect 10968 21641 10977 21675
rect 10977 21641 11011 21675
rect 11011 21641 11020 21675
rect 10968 21632 11020 21641
rect 16304 21632 16356 21684
rect 16672 21632 16724 21684
rect 18972 21632 19024 21684
rect 19616 21632 19668 21684
rect 22836 21632 22888 21684
rect 9588 21564 9640 21616
rect 9404 21428 9456 21480
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 15292 21564 15344 21616
rect 15936 21607 15988 21616
rect 15936 21573 15945 21607
rect 15945 21573 15979 21607
rect 15979 21573 15988 21607
rect 15936 21564 15988 21573
rect 16580 21564 16632 21616
rect 16764 21564 16816 21616
rect 17500 21564 17552 21616
rect 19064 21564 19116 21616
rect 20260 21564 20312 21616
rect 20996 21564 21048 21616
rect 12440 21428 12492 21480
rect 12716 21360 12768 21412
rect 5540 21292 5592 21344
rect 6184 21292 6236 21344
rect 9680 21335 9732 21344
rect 9680 21301 9689 21335
rect 9689 21301 9723 21335
rect 9723 21301 9732 21335
rect 9680 21292 9732 21301
rect 11060 21292 11112 21344
rect 11520 21292 11572 21344
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 14096 21428 14148 21480
rect 24492 21632 24544 21684
rect 23940 21564 23992 21616
rect 25044 21632 25096 21684
rect 27528 21632 27580 21684
rect 30564 21632 30616 21684
rect 36728 21632 36780 21684
rect 25688 21564 25740 21616
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 25964 21539 26016 21548
rect 25964 21505 25973 21539
rect 25973 21505 26007 21539
rect 26007 21505 26016 21539
rect 25964 21496 26016 21505
rect 29000 21564 29052 21616
rect 31576 21564 31628 21616
rect 29828 21496 29880 21548
rect 31944 21539 31996 21548
rect 31944 21505 31953 21539
rect 31953 21505 31987 21539
rect 31987 21505 31996 21539
rect 31944 21496 31996 21505
rect 32312 21496 32364 21548
rect 47860 21496 47912 21548
rect 16212 21471 16264 21480
rect 16212 21437 16221 21471
rect 16221 21437 16255 21471
rect 16255 21437 16264 21471
rect 16212 21428 16264 21437
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 14372 21360 14424 21412
rect 13728 21292 13780 21344
rect 14556 21292 14608 21344
rect 15568 21403 15620 21412
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 18696 21292 18748 21344
rect 18972 21471 19024 21480
rect 18972 21437 18981 21471
rect 18981 21437 19015 21471
rect 19015 21437 19024 21471
rect 18972 21428 19024 21437
rect 19064 21428 19116 21480
rect 21916 21428 21968 21480
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 24676 21428 24728 21480
rect 26240 21471 26292 21480
rect 26240 21437 26249 21471
rect 26249 21437 26283 21471
rect 26283 21437 26292 21471
rect 26240 21428 26292 21437
rect 26700 21428 26752 21480
rect 20168 21360 20220 21412
rect 22376 21360 22428 21412
rect 24768 21360 24820 21412
rect 27804 21471 27856 21480
rect 27804 21437 27813 21471
rect 27813 21437 27847 21471
rect 27847 21437 27856 21471
rect 27804 21428 27856 21437
rect 28356 21428 28408 21480
rect 28724 21471 28776 21480
rect 28724 21437 28733 21471
rect 28733 21437 28767 21471
rect 28767 21437 28776 21471
rect 28724 21428 28776 21437
rect 30104 21428 30156 21480
rect 19432 21292 19484 21344
rect 19708 21292 19760 21344
rect 20996 21335 21048 21344
rect 20996 21301 21005 21335
rect 21005 21301 21039 21335
rect 21039 21301 21048 21335
rect 20996 21292 21048 21301
rect 21916 21292 21968 21344
rect 24124 21292 24176 21344
rect 25228 21292 25280 21344
rect 30288 21360 30340 21412
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 31392 21360 31444 21412
rect 34520 21360 34572 21412
rect 37740 21360 37792 21412
rect 28448 21292 28500 21344
rect 30196 21335 30248 21344
rect 30196 21301 30205 21335
rect 30205 21301 30239 21335
rect 30239 21301 30248 21335
rect 30196 21292 30248 21301
rect 30656 21335 30708 21344
rect 30656 21301 30665 21335
rect 30665 21301 30699 21335
rect 30699 21301 30708 21335
rect 30656 21292 30708 21301
rect 31852 21292 31904 21344
rect 32496 21335 32548 21344
rect 32496 21301 32505 21335
rect 32505 21301 32539 21335
rect 32539 21301 32548 21335
rect 32496 21292 32548 21301
rect 32772 21292 32824 21344
rect 47860 21292 47912 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 6920 21088 6972 21140
rect 12164 21088 12216 21140
rect 12348 21088 12400 21140
rect 14924 21088 14976 21140
rect 15108 21088 15160 21140
rect 7012 21020 7064 21072
rect 4252 20995 4304 21004
rect 4252 20961 4261 20995
rect 4261 20961 4295 20995
rect 4295 20961 4304 20995
rect 4252 20952 4304 20961
rect 11796 21020 11848 21072
rect 12256 21020 12308 21072
rect 14188 21020 14240 21072
rect 14372 21020 14424 21072
rect 17316 21020 17368 21072
rect 8484 20995 8536 21004
rect 8484 20961 8493 20995
rect 8493 20961 8527 20995
rect 8527 20961 8536 20995
rect 8484 20952 8536 20961
rect 8576 20952 8628 21004
rect 11244 20952 11296 21004
rect 1860 20884 1912 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 7656 20884 7708 20936
rect 12072 20952 12124 21004
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 15016 20952 15068 21004
rect 2872 20816 2924 20868
rect 3792 20816 3844 20868
rect 5632 20816 5684 20868
rect 6184 20816 6236 20868
rect 8208 20859 8260 20868
rect 8208 20825 8217 20859
rect 8217 20825 8251 20859
rect 8251 20825 8260 20859
rect 8208 20816 8260 20825
rect 8576 20816 8628 20868
rect 9588 20816 9640 20868
rect 11336 20859 11388 20868
rect 11336 20825 11345 20859
rect 11345 20825 11379 20859
rect 11379 20825 11388 20859
rect 11336 20816 11388 20825
rect 15292 20952 15344 21004
rect 16396 20995 16448 21004
rect 16396 20961 16405 20995
rect 16405 20961 16439 20995
rect 16439 20961 16448 20995
rect 16396 20952 16448 20961
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 18696 20995 18748 21004
rect 18696 20961 18705 20995
rect 18705 20961 18739 20995
rect 18739 20961 18748 20995
rect 18696 20952 18748 20961
rect 22284 21020 22336 21072
rect 22468 21088 22520 21140
rect 25320 21088 25372 21140
rect 26332 21088 26384 21140
rect 24768 21020 24820 21072
rect 27528 21020 27580 21072
rect 28816 21020 28868 21072
rect 31944 21088 31996 21140
rect 32588 21088 32640 21140
rect 29184 21020 29236 21072
rect 32772 21020 32824 21072
rect 19708 20995 19760 21004
rect 19708 20961 19717 20995
rect 19717 20961 19751 20995
rect 19751 20961 19760 20995
rect 19708 20952 19760 20961
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 23848 20995 23900 21004
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 25320 20995 25372 21004
rect 25320 20961 25329 20995
rect 25329 20961 25363 20995
rect 25363 20961 25372 20995
rect 25320 20952 25372 20961
rect 27804 20952 27856 21004
rect 28540 20995 28592 21004
rect 28540 20961 28549 20995
rect 28549 20961 28583 20995
rect 28583 20961 28592 20995
rect 28540 20952 28592 20961
rect 30012 20995 30064 21004
rect 30012 20961 30021 20995
rect 30021 20961 30055 20995
rect 30055 20961 30064 20995
rect 30012 20952 30064 20961
rect 30564 20952 30616 21004
rect 31208 20952 31260 21004
rect 31668 20952 31720 21004
rect 36452 20952 36504 21004
rect 15200 20816 15252 20868
rect 5816 20748 5868 20800
rect 6368 20748 6420 20800
rect 7012 20748 7064 20800
rect 7564 20791 7616 20800
rect 7564 20757 7573 20791
rect 7573 20757 7607 20791
rect 7607 20757 7616 20791
rect 7564 20748 7616 20757
rect 9404 20748 9456 20800
rect 11428 20791 11480 20800
rect 11428 20757 11437 20791
rect 11437 20757 11471 20791
rect 11471 20757 11480 20791
rect 11428 20748 11480 20757
rect 11612 20748 11664 20800
rect 11888 20748 11940 20800
rect 13544 20748 13596 20800
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 14372 20748 14424 20800
rect 19064 20884 19116 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 24216 20884 24268 20936
rect 25780 20884 25832 20936
rect 26056 20927 26108 20936
rect 26056 20893 26065 20927
rect 26065 20893 26099 20927
rect 26099 20893 26108 20927
rect 26056 20884 26108 20893
rect 28448 20884 28500 20936
rect 28908 20884 28960 20936
rect 29552 20884 29604 20936
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 32680 20927 32732 20936
rect 32680 20893 32689 20927
rect 32689 20893 32723 20927
rect 32723 20893 32732 20927
rect 32680 20884 32732 20893
rect 19708 20816 19760 20868
rect 20996 20816 21048 20868
rect 16764 20748 16816 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 17500 20748 17552 20800
rect 17684 20748 17736 20800
rect 18880 20748 18932 20800
rect 21180 20791 21232 20800
rect 21180 20757 21189 20791
rect 21189 20757 21223 20791
rect 21223 20757 21232 20791
rect 21180 20748 21232 20757
rect 21824 20816 21876 20868
rect 21916 20748 21968 20800
rect 23572 20816 23624 20868
rect 26240 20816 26292 20868
rect 27344 20816 27396 20868
rect 22468 20791 22520 20800
rect 22468 20757 22477 20791
rect 22477 20757 22511 20791
rect 22511 20757 22520 20791
rect 22468 20748 22520 20757
rect 22560 20791 22612 20800
rect 22560 20757 22569 20791
rect 22569 20757 22603 20791
rect 22603 20757 22612 20791
rect 22560 20748 22612 20757
rect 22652 20748 22704 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 23940 20748 23992 20800
rect 30656 20816 30708 20868
rect 31852 20859 31904 20868
rect 31852 20825 31861 20859
rect 31861 20825 31895 20859
rect 31895 20825 31904 20859
rect 31852 20816 31904 20825
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 31944 20791 31996 20800
rect 31944 20757 31953 20791
rect 31953 20757 31987 20791
rect 31987 20757 31996 20791
rect 31944 20748 31996 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 3884 20476 3936 20528
rect 4344 20476 4396 20528
rect 6828 20544 6880 20596
rect 6920 20476 6972 20528
rect 9220 20476 9272 20528
rect 9404 20476 9456 20528
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 3976 20408 4028 20460
rect 3332 20340 3384 20392
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 6092 20408 6144 20460
rect 8668 20408 8720 20460
rect 11980 20408 12032 20460
rect 6828 20340 6880 20392
rect 7288 20383 7340 20392
rect 7288 20349 7297 20383
rect 7297 20349 7331 20383
rect 7331 20349 7340 20383
rect 7288 20340 7340 20349
rect 8852 20340 8904 20392
rect 9404 20383 9456 20392
rect 9404 20349 9413 20383
rect 9413 20349 9447 20383
rect 9447 20349 9456 20383
rect 9404 20340 9456 20349
rect 10968 20340 11020 20392
rect 5908 20272 5960 20324
rect 10692 20272 10744 20324
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 16948 20544 17000 20596
rect 17776 20544 17828 20596
rect 18512 20587 18564 20596
rect 18512 20553 18521 20587
rect 18521 20553 18555 20587
rect 18555 20553 18564 20587
rect 18512 20544 18564 20553
rect 18880 20587 18932 20596
rect 18880 20553 18889 20587
rect 18889 20553 18923 20587
rect 18923 20553 18932 20587
rect 18880 20544 18932 20553
rect 19432 20544 19484 20596
rect 15292 20476 15344 20528
rect 17224 20476 17276 20528
rect 13544 20408 13596 20460
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 15384 20408 15436 20460
rect 7656 20204 7708 20256
rect 8484 20204 8536 20256
rect 9036 20204 9088 20256
rect 10048 20204 10100 20256
rect 10876 20204 10928 20256
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 11612 20204 11664 20256
rect 13636 20204 13688 20256
rect 14556 20340 14608 20392
rect 15016 20340 15068 20392
rect 15200 20340 15252 20392
rect 21916 20476 21968 20528
rect 22468 20544 22520 20596
rect 23756 20544 23808 20596
rect 22100 20408 22152 20460
rect 23388 20408 23440 20460
rect 24216 20408 24268 20460
rect 25688 20408 25740 20460
rect 26056 20544 26108 20596
rect 26608 20544 26660 20596
rect 27528 20544 27580 20596
rect 29000 20544 29052 20596
rect 30840 20544 30892 20596
rect 27712 20476 27764 20528
rect 31760 20587 31812 20596
rect 31760 20553 31769 20587
rect 31769 20553 31803 20587
rect 31803 20553 31812 20587
rect 31760 20544 31812 20553
rect 27252 20408 27304 20460
rect 27620 20408 27672 20460
rect 28356 20451 28408 20460
rect 28356 20417 28365 20451
rect 28365 20417 28399 20451
rect 28399 20417 28408 20451
rect 28356 20408 28408 20417
rect 29736 20408 29788 20460
rect 36912 20408 36964 20460
rect 18788 20340 18840 20392
rect 18880 20340 18932 20392
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 16120 20272 16172 20324
rect 17408 20272 17460 20324
rect 20628 20340 20680 20392
rect 24676 20340 24728 20392
rect 25964 20340 26016 20392
rect 16580 20204 16632 20256
rect 17132 20204 17184 20256
rect 18880 20204 18932 20256
rect 22560 20272 22612 20324
rect 21824 20204 21876 20256
rect 22192 20204 22244 20256
rect 30196 20340 30248 20392
rect 30288 20340 30340 20392
rect 29644 20272 29696 20324
rect 25688 20204 25740 20256
rect 27252 20204 27304 20256
rect 28816 20204 28868 20256
rect 30196 20204 30248 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 5448 20000 5500 20052
rect 6276 19975 6328 19984
rect 6276 19941 6285 19975
rect 6285 19941 6319 19975
rect 6319 19941 6328 19975
rect 6276 19932 6328 19941
rect 8852 20000 8904 20052
rect 9496 20000 9548 20052
rect 10784 20000 10836 20052
rect 11796 20043 11848 20052
rect 11796 20009 11805 20043
rect 11805 20009 11839 20043
rect 11839 20009 11848 20043
rect 11796 20000 11848 20009
rect 12072 20000 12124 20052
rect 17132 20000 17184 20052
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 19340 20000 19392 20052
rect 19524 20000 19576 20052
rect 9036 19864 9088 19916
rect 13544 19932 13596 19984
rect 13728 19932 13780 19984
rect 14096 19932 14148 19984
rect 14556 19932 14608 19984
rect 10876 19907 10928 19916
rect 10876 19873 10885 19907
rect 10885 19873 10919 19907
rect 10919 19873 10928 19907
rect 10876 19864 10928 19873
rect 13360 19864 13412 19916
rect 15476 19864 15528 19916
rect 17500 19864 17552 19916
rect 17684 19907 17736 19916
rect 17684 19873 17693 19907
rect 17693 19873 17727 19907
rect 17727 19873 17736 19907
rect 17684 19864 17736 19873
rect 4436 19796 4488 19848
rect 10784 19796 10836 19848
rect 2872 19728 2924 19780
rect 4528 19728 4580 19780
rect 4804 19771 4856 19780
rect 4804 19737 4813 19771
rect 4813 19737 4847 19771
rect 4847 19737 4856 19771
rect 4804 19728 4856 19737
rect 6276 19728 6328 19780
rect 8668 19728 8720 19780
rect 8300 19660 8352 19712
rect 8852 19660 8904 19712
rect 9496 19728 9548 19780
rect 11060 19728 11112 19780
rect 14464 19796 14516 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 21548 19932 21600 19984
rect 49240 20000 49292 20052
rect 22744 19932 22796 19984
rect 11152 19660 11204 19712
rect 13268 19728 13320 19780
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 13912 19660 13964 19712
rect 14648 19660 14700 19712
rect 15292 19728 15344 19780
rect 18328 19728 18380 19780
rect 16396 19660 16448 19712
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 17684 19660 17736 19712
rect 17868 19660 17920 19712
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 18788 19864 18840 19916
rect 21180 19864 21232 19916
rect 23848 19907 23900 19916
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 19064 19796 19116 19848
rect 19708 19796 19760 19848
rect 21548 19796 21600 19848
rect 22284 19796 22336 19848
rect 23756 19839 23808 19848
rect 23756 19805 23765 19839
rect 23765 19805 23799 19839
rect 23799 19805 23808 19839
rect 23756 19796 23808 19805
rect 27804 19932 27856 19984
rect 26148 19864 26200 19916
rect 28632 19907 28684 19916
rect 28632 19873 28641 19907
rect 28641 19873 28675 19907
rect 28675 19873 28684 19907
rect 28632 19864 28684 19873
rect 29000 19864 29052 19916
rect 31760 19932 31812 19984
rect 46940 19932 46992 19984
rect 32036 19864 32088 19916
rect 18972 19728 19024 19780
rect 19340 19728 19392 19780
rect 19892 19728 19944 19780
rect 21916 19728 21968 19780
rect 22744 19771 22796 19780
rect 22744 19737 22753 19771
rect 22753 19737 22787 19771
rect 22787 19737 22796 19771
rect 22744 19728 22796 19737
rect 25596 19728 25648 19780
rect 25780 19796 25832 19848
rect 27252 19796 27304 19848
rect 27988 19796 28040 19848
rect 28448 19796 28500 19848
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 30380 19796 30432 19848
rect 31668 19796 31720 19848
rect 26424 19728 26476 19780
rect 23296 19703 23348 19712
rect 23296 19669 23305 19703
rect 23305 19669 23339 19703
rect 23339 19669 23348 19703
rect 23296 19660 23348 19669
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 23756 19660 23808 19712
rect 27988 19703 28040 19712
rect 27988 19669 27997 19703
rect 27997 19669 28031 19703
rect 28031 19669 28040 19703
rect 27988 19660 28040 19669
rect 29736 19660 29788 19712
rect 30380 19703 30432 19712
rect 30380 19669 30389 19703
rect 30389 19669 30423 19703
rect 30423 19669 30432 19703
rect 30380 19660 30432 19669
rect 37188 19660 37240 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 5264 19499 5316 19508
rect 5264 19465 5273 19499
rect 5273 19465 5307 19499
rect 5307 19465 5316 19499
rect 5264 19456 5316 19465
rect 6736 19456 6788 19508
rect 7564 19456 7616 19508
rect 10692 19456 10744 19508
rect 11888 19456 11940 19508
rect 14096 19456 14148 19508
rect 4160 19388 4212 19440
rect 2136 19320 2188 19372
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3608 19363 3660 19372
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 8668 19320 8720 19372
rect 9128 19388 9180 19440
rect 10324 19320 10376 19372
rect 4252 19252 4304 19304
rect 6552 19252 6604 19304
rect 4988 19184 5040 19236
rect 5356 19184 5408 19236
rect 5448 19184 5500 19236
rect 10140 19295 10192 19304
rect 10140 19261 10149 19295
rect 10149 19261 10183 19295
rect 10183 19261 10192 19295
rect 10140 19252 10192 19261
rect 6920 19184 6972 19236
rect 10232 19184 10284 19236
rect 11428 19388 11480 19440
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 11060 19252 11112 19304
rect 11612 19320 11664 19372
rect 11980 19388 12032 19440
rect 13268 19388 13320 19440
rect 13820 19388 13872 19440
rect 13912 19431 13964 19440
rect 13912 19397 13921 19431
rect 13921 19397 13955 19431
rect 13955 19397 13964 19431
rect 13912 19388 13964 19397
rect 14648 19456 14700 19508
rect 13452 19320 13504 19372
rect 14464 19388 14516 19440
rect 17960 19456 18012 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 19340 19456 19392 19508
rect 23296 19456 23348 19508
rect 17132 19388 17184 19440
rect 14556 19320 14608 19372
rect 13728 19252 13780 19304
rect 15292 19320 15344 19372
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 4620 19116 4672 19168
rect 6092 19116 6144 19168
rect 6460 19116 6512 19168
rect 8484 19116 8536 19168
rect 9496 19116 9548 19168
rect 10784 19116 10836 19168
rect 13820 19116 13872 19168
rect 14924 19295 14976 19304
rect 14924 19261 14933 19295
rect 14933 19261 14967 19295
rect 14967 19261 14976 19295
rect 14924 19252 14976 19261
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 19432 19388 19484 19440
rect 22652 19388 22704 19440
rect 25688 19456 25740 19508
rect 26240 19456 26292 19508
rect 26792 19456 26844 19508
rect 27252 19499 27304 19508
rect 27252 19465 27261 19499
rect 27261 19465 27295 19499
rect 27295 19465 27304 19499
rect 27252 19456 27304 19465
rect 27712 19499 27764 19508
rect 27712 19465 27721 19499
rect 27721 19465 27755 19499
rect 27755 19465 27764 19499
rect 27712 19456 27764 19465
rect 27804 19456 27856 19508
rect 30380 19456 30432 19508
rect 32128 19456 32180 19508
rect 17684 19320 17736 19372
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 18512 19320 18564 19372
rect 19064 19320 19116 19372
rect 21916 19320 21968 19372
rect 25320 19388 25372 19440
rect 28816 19388 28868 19440
rect 17316 19252 17368 19304
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 17684 19184 17736 19236
rect 14464 19116 14516 19168
rect 16028 19116 16080 19168
rect 17776 19116 17828 19168
rect 18696 19116 18748 19168
rect 20628 19252 20680 19304
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 22836 19320 22888 19372
rect 24492 19320 24544 19372
rect 24860 19252 24912 19304
rect 22008 19227 22060 19236
rect 22008 19193 22017 19227
rect 22017 19193 22051 19227
rect 22051 19193 22060 19227
rect 22008 19184 22060 19193
rect 22100 19184 22152 19236
rect 25044 19320 25096 19372
rect 29644 19320 29696 19372
rect 30656 19363 30708 19372
rect 30656 19329 30665 19363
rect 30665 19329 30699 19363
rect 30699 19329 30708 19363
rect 30656 19320 30708 19329
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 26884 19252 26936 19304
rect 27436 19295 27488 19304
rect 27436 19261 27445 19295
rect 27445 19261 27479 19295
rect 27479 19261 27488 19295
rect 27436 19252 27488 19261
rect 28264 19295 28316 19304
rect 28264 19261 28273 19295
rect 28273 19261 28307 19295
rect 28307 19261 28316 19295
rect 28264 19252 28316 19261
rect 30932 19252 30984 19304
rect 31852 19320 31904 19372
rect 23480 19116 23532 19168
rect 23572 19116 23624 19168
rect 24124 19116 24176 19168
rect 27804 19116 27856 19168
rect 28632 19116 28684 19168
rect 30288 19116 30340 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 1400 18776 1452 18828
rect 15016 18912 15068 18964
rect 8576 18887 8628 18896
rect 8576 18853 8585 18887
rect 8585 18853 8619 18887
rect 8619 18853 8628 18887
rect 8576 18844 8628 18853
rect 8484 18776 8536 18828
rect 4528 18708 4580 18760
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 8208 18708 8260 18760
rect 9128 18776 9180 18828
rect 9864 18844 9916 18896
rect 9956 18819 10008 18828
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 10324 18776 10376 18828
rect 10508 18776 10560 18828
rect 11152 18776 11204 18828
rect 6276 18640 6328 18692
rect 6736 18640 6788 18692
rect 2504 18572 2556 18624
rect 3424 18572 3476 18624
rect 4712 18572 4764 18624
rect 4804 18572 4856 18624
rect 8760 18640 8812 18692
rect 8944 18640 8996 18692
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 11244 18708 11296 18760
rect 13544 18819 13596 18828
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 8576 18572 8628 18624
rect 9128 18572 9180 18624
rect 9220 18572 9272 18624
rect 10048 18640 10100 18692
rect 10232 18640 10284 18692
rect 11704 18640 11756 18692
rect 12808 18683 12860 18692
rect 12808 18649 12817 18683
rect 12817 18649 12851 18683
rect 12851 18649 12860 18683
rect 12808 18640 12860 18649
rect 22008 18912 22060 18964
rect 22560 18912 22612 18964
rect 17224 18844 17276 18896
rect 16212 18776 16264 18828
rect 16764 18776 16816 18828
rect 18328 18844 18380 18896
rect 21088 18844 21140 18896
rect 19708 18776 19760 18828
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 21548 18776 21600 18828
rect 30748 18912 30800 18964
rect 29736 18844 29788 18896
rect 30932 18844 30984 18896
rect 48504 18912 48556 18964
rect 23664 18776 23716 18828
rect 25780 18776 25832 18828
rect 26424 18776 26476 18828
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 16948 18708 17000 18760
rect 18604 18708 18656 18760
rect 15476 18683 15528 18692
rect 15476 18649 15485 18683
rect 15485 18649 15519 18683
rect 15519 18649 15528 18683
rect 15476 18640 15528 18649
rect 15936 18640 15988 18692
rect 11244 18572 11296 18624
rect 11612 18572 11664 18624
rect 12716 18572 12768 18624
rect 15384 18572 15436 18624
rect 16396 18572 16448 18624
rect 19708 18640 19760 18692
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 17040 18572 17092 18624
rect 17132 18572 17184 18624
rect 18696 18572 18748 18624
rect 20260 18572 20312 18624
rect 22100 18572 22152 18624
rect 22928 18640 22980 18692
rect 24124 18708 24176 18760
rect 26792 18708 26844 18760
rect 23848 18640 23900 18692
rect 23020 18572 23072 18624
rect 23388 18615 23440 18624
rect 23388 18581 23397 18615
rect 23397 18581 23431 18615
rect 23431 18581 23440 18615
rect 23388 18572 23440 18581
rect 23664 18572 23716 18624
rect 25964 18640 26016 18692
rect 25136 18572 25188 18624
rect 27712 18708 27764 18760
rect 29828 18708 29880 18760
rect 27068 18640 27120 18692
rect 46848 18776 46900 18828
rect 29736 18615 29788 18624
rect 29736 18581 29745 18615
rect 29745 18581 29779 18615
rect 29779 18581 29788 18615
rect 29736 18572 29788 18581
rect 30104 18615 30156 18624
rect 30104 18581 30113 18615
rect 30113 18581 30147 18615
rect 30147 18581 30156 18615
rect 30104 18572 30156 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 5908 18368 5960 18420
rect 6736 18368 6788 18420
rect 7288 18368 7340 18420
rect 8944 18368 8996 18420
rect 7932 18300 7984 18352
rect 9128 18300 9180 18352
rect 10140 18368 10192 18420
rect 13360 18368 13412 18420
rect 15016 18411 15068 18420
rect 15016 18377 15025 18411
rect 15025 18377 15059 18411
rect 15059 18377 15068 18411
rect 15016 18368 15068 18377
rect 17684 18368 17736 18420
rect 4252 18232 4304 18284
rect 5632 18275 5684 18284
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 6460 18232 6512 18284
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 3700 18164 3752 18216
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 6092 18164 6144 18216
rect 4712 18096 4764 18148
rect 8392 18232 8444 18284
rect 12808 18300 12860 18352
rect 10232 18232 10284 18284
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 7196 18207 7248 18216
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7196 18164 7248 18173
rect 8576 18164 8628 18216
rect 9496 18164 9548 18216
rect 12072 18164 12124 18216
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 14096 18300 14148 18352
rect 14648 18300 14700 18352
rect 21456 18368 21508 18420
rect 15936 18232 15988 18284
rect 16580 18232 16632 18284
rect 15108 18164 15160 18216
rect 16948 18164 17000 18216
rect 3424 18028 3476 18080
rect 3700 18028 3752 18080
rect 5448 18028 5500 18080
rect 9588 18028 9640 18080
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 9864 18028 9916 18080
rect 10416 18028 10468 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 12164 18096 12216 18148
rect 16396 18096 16448 18148
rect 16856 18096 16908 18148
rect 17132 18096 17184 18148
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 17592 18232 17644 18284
rect 20260 18232 20312 18284
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 22652 18368 22704 18420
rect 22928 18368 22980 18420
rect 23480 18368 23532 18420
rect 26792 18411 26844 18420
rect 26792 18377 26801 18411
rect 26801 18377 26835 18411
rect 26835 18377 26844 18411
rect 26792 18368 26844 18377
rect 30104 18368 30156 18420
rect 30748 18411 30800 18420
rect 30748 18377 30757 18411
rect 30757 18377 30791 18411
rect 30791 18377 30800 18411
rect 30748 18368 30800 18377
rect 23020 18300 23072 18352
rect 23848 18300 23900 18352
rect 26056 18343 26108 18352
rect 26056 18309 26065 18343
rect 26065 18309 26099 18343
rect 26099 18309 26108 18343
rect 26056 18300 26108 18309
rect 21088 18232 21140 18241
rect 25044 18232 25096 18284
rect 28264 18300 28316 18352
rect 28632 18300 28684 18352
rect 29644 18300 29696 18352
rect 30656 18343 30708 18352
rect 30656 18309 30665 18343
rect 30665 18309 30699 18343
rect 30699 18309 30708 18343
rect 31300 18343 31352 18352
rect 30656 18300 30708 18309
rect 31300 18309 31309 18343
rect 31309 18309 31343 18343
rect 31343 18309 31352 18343
rect 31300 18300 31352 18309
rect 18144 18164 18196 18216
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 18972 18164 19024 18216
rect 19800 18164 19852 18216
rect 12716 18028 12768 18080
rect 13820 18028 13872 18080
rect 15660 18028 15712 18080
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 16764 18028 16816 18080
rect 18328 18028 18380 18080
rect 19708 18096 19760 18148
rect 21180 18207 21232 18216
rect 21180 18173 21189 18207
rect 21189 18173 21223 18207
rect 21223 18173 21232 18207
rect 21180 18164 21232 18173
rect 20996 18096 21048 18148
rect 26240 18164 26292 18216
rect 27068 18164 27120 18216
rect 30380 18096 30432 18148
rect 34612 18164 34664 18216
rect 41420 18096 41472 18148
rect 24676 18028 24728 18080
rect 27344 18028 27396 18080
rect 29828 18071 29880 18080
rect 29828 18037 29837 18071
rect 29837 18037 29871 18071
rect 29871 18037 29880 18071
rect 29828 18028 29880 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 8392 17824 8444 17876
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 1860 17756 1912 17808
rect 6184 17756 6236 17808
rect 7840 17799 7892 17808
rect 7840 17765 7849 17799
rect 7849 17765 7883 17799
rect 7883 17765 7892 17799
rect 7840 17756 7892 17765
rect 8024 17756 8076 17808
rect 8852 17756 8904 17808
rect 10324 17756 10376 17808
rect 11520 17756 11572 17808
rect 7932 17688 7984 17740
rect 4160 17620 4212 17672
rect 4620 17620 4672 17672
rect 6276 17620 6328 17672
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7656 17620 7708 17672
rect 8392 17620 8444 17672
rect 8576 17620 8628 17672
rect 9404 17688 9456 17740
rect 10048 17688 10100 17740
rect 11428 17688 11480 17740
rect 10876 17620 10928 17672
rect 13452 17824 13504 17876
rect 13728 17867 13780 17876
rect 13728 17833 13737 17867
rect 13737 17833 13771 17867
rect 13771 17833 13780 17867
rect 13728 17824 13780 17833
rect 15844 17824 15896 17876
rect 16212 17824 16264 17876
rect 16396 17824 16448 17876
rect 13268 17756 13320 17808
rect 14924 17756 14976 17808
rect 12624 17688 12676 17740
rect 12808 17688 12860 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 16948 17688 17000 17740
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 15016 17620 15068 17672
rect 940 17552 992 17604
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 2136 17484 2188 17536
rect 4804 17484 4856 17536
rect 7472 17552 7524 17604
rect 8024 17484 8076 17536
rect 9220 17552 9272 17604
rect 9404 17552 9456 17604
rect 12256 17552 12308 17604
rect 12716 17552 12768 17604
rect 13820 17552 13872 17604
rect 14924 17552 14976 17604
rect 15292 17552 15344 17604
rect 12072 17484 12124 17536
rect 15016 17484 15068 17536
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 15200 17484 15252 17536
rect 15936 17484 15988 17536
rect 16304 17484 16356 17536
rect 17776 17688 17828 17740
rect 21088 17756 21140 17808
rect 19432 17731 19484 17740
rect 19432 17697 19441 17731
rect 19441 17697 19475 17731
rect 19475 17697 19484 17731
rect 19432 17688 19484 17697
rect 20996 17688 21048 17740
rect 22284 17756 22336 17808
rect 26240 17756 26292 17808
rect 28448 17756 28500 17808
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 20444 17620 20496 17672
rect 24584 17688 24636 17740
rect 24676 17688 24728 17740
rect 25780 17688 25832 17740
rect 28356 17688 28408 17740
rect 22008 17620 22060 17672
rect 29644 17688 29696 17740
rect 30288 17731 30340 17740
rect 30288 17697 30297 17731
rect 30297 17697 30331 17731
rect 30331 17697 30340 17731
rect 30288 17688 30340 17697
rect 28816 17620 28868 17672
rect 31024 17620 31076 17672
rect 34520 17620 34572 17672
rect 18880 17552 18932 17604
rect 18328 17484 18380 17536
rect 18696 17527 18748 17536
rect 18696 17493 18705 17527
rect 18705 17493 18739 17527
rect 18739 17493 18748 17527
rect 18696 17484 18748 17493
rect 19892 17484 19944 17536
rect 23848 17552 23900 17604
rect 25136 17595 25188 17604
rect 21916 17484 21968 17536
rect 23480 17484 23532 17536
rect 25136 17561 25145 17595
rect 25145 17561 25179 17595
rect 25179 17561 25188 17595
rect 25136 17552 25188 17561
rect 26792 17552 26844 17604
rect 27344 17595 27396 17604
rect 27344 17561 27353 17595
rect 27353 17561 27387 17595
rect 27387 17561 27396 17595
rect 27344 17552 27396 17561
rect 24400 17527 24452 17536
rect 24400 17493 24409 17527
rect 24409 17493 24443 17527
rect 24443 17493 24452 17527
rect 30932 17552 30984 17604
rect 24400 17484 24452 17493
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 28816 17484 28868 17493
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 5080 17212 5132 17264
rect 7748 17280 7800 17332
rect 9128 17280 9180 17332
rect 9496 17280 9548 17332
rect 8392 17255 8444 17264
rect 8392 17221 8401 17255
rect 8401 17221 8435 17255
rect 8435 17221 8444 17255
rect 8392 17212 8444 17221
rect 3792 17144 3844 17196
rect 1124 17076 1176 17128
rect 4436 17076 4488 17128
rect 6092 17144 6144 17196
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 8576 17144 8628 17196
rect 9496 17144 9548 17196
rect 11428 17212 11480 17264
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 12532 17323 12584 17332
rect 12532 17289 12541 17323
rect 12541 17289 12575 17323
rect 12575 17289 12584 17323
rect 12532 17280 12584 17289
rect 14648 17280 14700 17332
rect 14832 17280 14884 17332
rect 17040 17280 17092 17332
rect 17776 17280 17828 17332
rect 17868 17280 17920 17332
rect 13820 17212 13872 17264
rect 14280 17212 14332 17264
rect 18328 17212 18380 17264
rect 20076 17212 20128 17264
rect 2504 17008 2556 17060
rect 5172 16940 5224 16992
rect 5356 16940 5408 16992
rect 5632 17008 5684 17060
rect 5816 17119 5868 17128
rect 5816 17085 5825 17119
rect 5825 17085 5859 17119
rect 5859 17085 5868 17119
rect 5816 17076 5868 17085
rect 7840 17076 7892 17128
rect 8208 17076 8260 17128
rect 8760 17076 8812 17128
rect 9404 17076 9456 17128
rect 9772 17076 9824 17128
rect 10140 17119 10192 17128
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 10692 17076 10744 17128
rect 12532 17144 12584 17196
rect 13912 17144 13964 17196
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 14924 17187 14976 17196
rect 14924 17153 14933 17187
rect 14933 17153 14967 17187
rect 14967 17153 14976 17187
rect 14924 17144 14976 17153
rect 15292 17144 15344 17196
rect 15844 17144 15896 17196
rect 17132 17144 17184 17196
rect 17224 17187 17276 17196
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 20904 17212 20956 17264
rect 23940 17280 23992 17332
rect 24216 17280 24268 17332
rect 22284 17212 22336 17264
rect 23112 17212 23164 17264
rect 28816 17280 28868 17332
rect 29644 17280 29696 17332
rect 30196 17280 30248 17332
rect 30932 17323 30984 17332
rect 30932 17289 30941 17323
rect 30941 17289 30975 17323
rect 30975 17289 30984 17323
rect 30932 17280 30984 17289
rect 26240 17212 26292 17264
rect 26792 17255 26844 17264
rect 26792 17221 26801 17255
rect 26801 17221 26835 17255
rect 26835 17221 26844 17255
rect 26792 17212 26844 17221
rect 13728 17076 13780 17128
rect 14188 17119 14240 17128
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 15476 17076 15528 17128
rect 15936 17076 15988 17128
rect 6460 16983 6512 16992
rect 6460 16949 6469 16983
rect 6469 16949 6503 16983
rect 6503 16949 6512 16983
rect 6460 16940 6512 16949
rect 6644 17008 6696 17060
rect 8576 17008 8628 17060
rect 9404 16940 9456 16992
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 9588 16940 9640 16992
rect 12072 17008 12124 17060
rect 17776 17076 17828 17128
rect 17960 17008 18012 17060
rect 18972 17076 19024 17128
rect 22652 17144 22704 17196
rect 20352 17076 20404 17128
rect 21088 17008 21140 17060
rect 11612 16940 11664 16992
rect 12716 16940 12768 16992
rect 15752 16940 15804 16992
rect 16488 16940 16540 16992
rect 17408 16940 17460 16992
rect 17500 16940 17552 16992
rect 19892 16983 19944 16992
rect 19892 16949 19901 16983
rect 19901 16949 19935 16983
rect 19935 16949 19944 16983
rect 19892 16940 19944 16949
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 21916 17076 21968 17128
rect 21824 17008 21876 17060
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 24400 17144 24452 17196
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 28356 17212 28408 17264
rect 31024 17212 31076 17264
rect 23756 17119 23808 17128
rect 23756 17085 23765 17119
rect 23765 17085 23799 17119
rect 23799 17085 23808 17119
rect 23756 17076 23808 17085
rect 23848 17119 23900 17128
rect 23848 17085 23857 17119
rect 23857 17085 23891 17119
rect 23891 17085 23900 17119
rect 23848 17076 23900 17085
rect 24584 17076 24636 17128
rect 27620 17076 27672 17128
rect 30288 17076 30340 17128
rect 30196 17008 30248 17060
rect 34520 17212 34572 17264
rect 48320 17212 48372 17264
rect 21548 16940 21600 16992
rect 21732 16940 21784 16992
rect 23296 16983 23348 16992
rect 23296 16949 23305 16983
rect 23305 16949 23339 16983
rect 23339 16949 23348 16983
rect 23296 16940 23348 16949
rect 24584 16940 24636 16992
rect 25044 16940 25096 16992
rect 25136 16940 25188 16992
rect 25964 16940 26016 16992
rect 27252 16940 27304 16992
rect 47216 17008 47268 17060
rect 47032 16940 47084 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 5080 16736 5132 16788
rect 5724 16736 5776 16788
rect 2596 16668 2648 16720
rect 6184 16668 6236 16720
rect 9220 16736 9272 16788
rect 10416 16736 10468 16788
rect 11520 16736 11572 16788
rect 11888 16736 11940 16788
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 12624 16736 12676 16788
rect 13728 16736 13780 16788
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 6828 16600 6880 16652
rect 8208 16600 8260 16652
rect 9312 16668 9364 16720
rect 9404 16668 9456 16720
rect 18880 16736 18932 16788
rect 14556 16668 14608 16720
rect 15016 16711 15068 16720
rect 15016 16677 15025 16711
rect 15025 16677 15059 16711
rect 15059 16677 15068 16711
rect 15016 16668 15068 16677
rect 15568 16668 15620 16720
rect 19708 16736 19760 16788
rect 20076 16736 20128 16788
rect 23756 16736 23808 16788
rect 30196 16736 30248 16788
rect 22008 16668 22060 16720
rect 25688 16711 25740 16720
rect 1216 16464 1268 16516
rect 4896 16575 4948 16584
rect 4896 16541 4905 16575
rect 4905 16541 4939 16575
rect 4939 16541 4948 16575
rect 4896 16532 4948 16541
rect 5724 16464 5776 16516
rect 7288 16464 7340 16516
rect 7748 16464 7800 16516
rect 6736 16396 6788 16448
rect 6920 16396 6972 16448
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 8208 16396 8260 16405
rect 9220 16507 9272 16516
rect 9220 16473 9229 16507
rect 9229 16473 9263 16507
rect 9263 16473 9272 16507
rect 9220 16464 9272 16473
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 11612 16600 11664 16652
rect 10968 16532 11020 16584
rect 12532 16600 12584 16652
rect 14280 16600 14332 16652
rect 14464 16600 14516 16652
rect 15752 16600 15804 16652
rect 16304 16600 16356 16652
rect 17224 16600 17276 16652
rect 11796 16464 11848 16516
rect 15292 16532 15344 16584
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 15568 16532 15620 16584
rect 20444 16600 20496 16652
rect 20720 16600 20772 16652
rect 22652 16643 22704 16652
rect 22652 16609 22661 16643
rect 22661 16609 22695 16643
rect 22695 16609 22704 16643
rect 22652 16600 22704 16609
rect 23756 16643 23808 16652
rect 23756 16609 23765 16643
rect 23765 16609 23799 16643
rect 23799 16609 23808 16643
rect 23756 16600 23808 16609
rect 25044 16600 25096 16652
rect 25688 16677 25697 16711
rect 25697 16677 25731 16711
rect 25731 16677 25740 16711
rect 25688 16668 25740 16677
rect 25964 16668 26016 16720
rect 25780 16600 25832 16652
rect 25872 16643 25924 16652
rect 25872 16609 25881 16643
rect 25881 16609 25915 16643
rect 25915 16609 25924 16643
rect 25872 16600 25924 16609
rect 26976 16600 27028 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27252 16643 27304 16652
rect 27252 16609 27261 16643
rect 27261 16609 27295 16643
rect 27295 16609 27304 16643
rect 27252 16600 27304 16609
rect 27804 16600 27856 16652
rect 28264 16643 28316 16652
rect 28264 16609 28273 16643
rect 28273 16609 28307 16643
rect 28307 16609 28316 16643
rect 28264 16600 28316 16609
rect 29000 16600 29052 16652
rect 17776 16532 17828 16584
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 23296 16532 23348 16584
rect 23664 16532 23716 16584
rect 24216 16532 24268 16584
rect 24492 16532 24544 16584
rect 17960 16464 18012 16516
rect 10508 16396 10560 16448
rect 13176 16396 13228 16448
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 14372 16396 14424 16448
rect 15568 16396 15620 16448
rect 16212 16396 16264 16448
rect 16488 16396 16540 16448
rect 16764 16396 16816 16448
rect 19984 16464 20036 16516
rect 21088 16464 21140 16516
rect 18972 16396 19024 16448
rect 23388 16464 23440 16516
rect 25596 16532 25648 16584
rect 21548 16396 21600 16448
rect 22468 16396 22520 16448
rect 23848 16396 23900 16448
rect 24584 16396 24636 16448
rect 25136 16396 25188 16448
rect 25872 16396 25924 16448
rect 27620 16532 27672 16584
rect 28448 16464 28500 16516
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 3884 16192 3936 16244
rect 4896 16192 4948 16244
rect 5632 16192 5684 16244
rect 6000 16192 6052 16244
rect 7380 16192 7432 16244
rect 4344 16167 4396 16176
rect 4344 16133 4353 16167
rect 4353 16133 4387 16167
rect 4387 16133 4396 16167
rect 4344 16124 4396 16133
rect 5448 16124 5500 16176
rect 6644 16124 6696 16176
rect 7104 16124 7156 16176
rect 1860 16056 1912 16108
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 7012 16056 7064 16108
rect 12532 16192 12584 16244
rect 13728 16235 13780 16244
rect 13728 16201 13737 16235
rect 13737 16201 13771 16235
rect 13771 16201 13780 16235
rect 13728 16192 13780 16201
rect 16304 16192 16356 16244
rect 1124 15988 1176 16040
rect 6092 15988 6144 16040
rect 6368 15988 6420 16040
rect 7564 15988 7616 16040
rect 4436 15920 4488 15972
rect 8760 16124 8812 16176
rect 10048 16124 10100 16176
rect 12256 16124 12308 16176
rect 16488 16124 16540 16176
rect 8484 16099 8536 16108
rect 8484 16065 8493 16099
rect 8493 16065 8527 16099
rect 8527 16065 8536 16099
rect 8484 16056 8536 16065
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 10968 16056 11020 16108
rect 8208 15988 8260 16040
rect 9956 15988 10008 16040
rect 10140 15988 10192 16040
rect 10876 15988 10928 16040
rect 11796 16056 11848 16108
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 14924 16056 14976 16108
rect 16396 16056 16448 16108
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 17592 16192 17644 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 18696 16192 18748 16244
rect 21180 16192 21232 16244
rect 21456 16192 21508 16244
rect 16672 16124 16724 16176
rect 17592 16056 17644 16108
rect 11244 15988 11296 16040
rect 11428 15988 11480 16040
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12256 16031 12308 16040
rect 12256 15997 12265 16031
rect 12265 15997 12299 16031
rect 12299 15997 12308 16031
rect 12256 15988 12308 15997
rect 12624 15988 12676 16040
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 5816 15852 5868 15904
rect 10784 15920 10836 15972
rect 10968 15963 11020 15972
rect 10968 15929 10977 15963
rect 10977 15929 11011 15963
rect 11011 15929 11020 15963
rect 10968 15920 11020 15929
rect 8760 15852 8812 15904
rect 9864 15852 9916 15904
rect 11704 15852 11756 15904
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 15568 15988 15620 16040
rect 18880 16124 18932 16176
rect 24952 16192 25004 16244
rect 27620 16192 27672 16244
rect 27804 16192 27856 16244
rect 19156 16056 19208 16108
rect 19432 16056 19484 16108
rect 20076 16056 20128 16108
rect 14004 15852 14056 15904
rect 17500 15920 17552 15972
rect 21640 15988 21692 16040
rect 22376 16056 22428 16108
rect 23664 16099 23716 16108
rect 23664 16065 23673 16099
rect 23673 16065 23707 16099
rect 23707 16065 23716 16099
rect 23664 16056 23716 16065
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 22836 15920 22888 15972
rect 23848 15988 23900 16040
rect 24032 15988 24084 16040
rect 25412 16124 25464 16176
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 26240 16056 26292 16108
rect 27068 16056 27120 16108
rect 27252 15988 27304 16040
rect 20168 15852 20220 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 22192 15852 22244 15904
rect 25228 15852 25280 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 5448 15648 5500 15700
rect 6276 15648 6328 15700
rect 7196 15648 7248 15700
rect 8208 15648 8260 15700
rect 3792 15580 3844 15632
rect 1308 15512 1360 15564
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 3424 15444 3476 15496
rect 4068 15444 4120 15496
rect 5540 15512 5592 15564
rect 5816 15512 5868 15564
rect 8668 15648 8720 15700
rect 10048 15648 10100 15700
rect 10416 15648 10468 15700
rect 13360 15648 13412 15700
rect 14556 15648 14608 15700
rect 14740 15648 14792 15700
rect 15936 15648 15988 15700
rect 17776 15648 17828 15700
rect 8576 15580 8628 15632
rect 9128 15580 9180 15632
rect 9220 15580 9272 15632
rect 8484 15512 8536 15564
rect 9404 15512 9456 15564
rect 10416 15512 10468 15564
rect 10784 15512 10836 15564
rect 12072 15623 12124 15632
rect 12072 15589 12081 15623
rect 12081 15589 12115 15623
rect 12115 15589 12124 15623
rect 12072 15580 12124 15589
rect 13636 15580 13688 15632
rect 19892 15623 19944 15632
rect 19892 15589 19901 15623
rect 19901 15589 19935 15623
rect 19935 15589 19944 15623
rect 19892 15580 19944 15589
rect 21640 15648 21692 15700
rect 24584 15648 24636 15700
rect 29736 15648 29788 15700
rect 12808 15512 12860 15564
rect 14372 15512 14424 15564
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 6092 15308 6144 15360
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 6644 15444 6696 15496
rect 7380 15444 7432 15496
rect 8116 15444 8168 15496
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 15476 15444 15528 15496
rect 8484 15376 8536 15428
rect 9220 15419 9272 15428
rect 9220 15385 9229 15419
rect 9229 15385 9263 15419
rect 9263 15385 9272 15419
rect 9220 15376 9272 15385
rect 11336 15419 11388 15428
rect 11336 15385 11345 15419
rect 11345 15385 11379 15419
rect 11379 15385 11388 15419
rect 11336 15376 11388 15385
rect 16028 15376 16080 15428
rect 20076 15512 20128 15564
rect 21088 15512 21140 15564
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 22100 15512 22152 15564
rect 22376 15444 22428 15496
rect 26976 15580 27028 15632
rect 34520 15580 34572 15632
rect 25780 15555 25832 15564
rect 25780 15521 25789 15555
rect 25789 15521 25823 15555
rect 25823 15521 25832 15555
rect 25780 15512 25832 15521
rect 23296 15444 23348 15496
rect 25596 15487 25648 15496
rect 25596 15453 25605 15487
rect 25605 15453 25639 15487
rect 25639 15453 25648 15487
rect 25596 15444 25648 15453
rect 17316 15419 17368 15428
rect 7380 15308 7432 15360
rect 7472 15308 7524 15360
rect 8576 15308 8628 15360
rect 9588 15308 9640 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 11428 15308 11480 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 13728 15308 13780 15360
rect 13912 15308 13964 15360
rect 15476 15351 15528 15360
rect 15476 15317 15485 15351
rect 15485 15317 15519 15351
rect 15519 15317 15528 15351
rect 17316 15385 17325 15419
rect 17325 15385 17359 15419
rect 17359 15385 17368 15419
rect 17316 15376 17368 15385
rect 17592 15376 17644 15428
rect 20260 15376 20312 15428
rect 15476 15308 15528 15317
rect 16396 15308 16448 15360
rect 17408 15308 17460 15360
rect 19340 15308 19392 15360
rect 22652 15376 22704 15428
rect 23572 15376 23624 15428
rect 23940 15419 23992 15428
rect 23940 15385 23949 15419
rect 23949 15385 23983 15419
rect 23983 15385 23992 15419
rect 23940 15376 23992 15385
rect 25412 15376 25464 15428
rect 26332 15376 26384 15428
rect 21916 15308 21968 15360
rect 22376 15351 22428 15360
rect 22376 15317 22385 15351
rect 22385 15317 22419 15351
rect 22419 15317 22428 15351
rect 22376 15308 22428 15317
rect 23480 15308 23532 15360
rect 23848 15308 23900 15360
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 40776 15308 40828 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 3516 15147 3568 15156
rect 3516 15113 3525 15147
rect 3525 15113 3559 15147
rect 3559 15113 3568 15147
rect 3516 15104 3568 15113
rect 4804 15104 4856 15156
rect 5908 15104 5960 15156
rect 6184 15104 6236 15156
rect 4712 15036 4764 15088
rect 5448 15036 5500 15088
rect 5724 15036 5776 15088
rect 3700 15011 3752 15020
rect 3700 14977 3709 15011
rect 3709 14977 3743 15011
rect 3743 14977 3752 15011
rect 3700 14968 3752 14977
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 5908 14968 5960 15020
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6644 14968 6696 14977
rect 7932 14968 7984 15020
rect 8576 15011 8628 15020
rect 8576 14977 8585 15011
rect 8585 14977 8619 15011
rect 8619 14977 8628 15011
rect 8576 14968 8628 14977
rect 9312 15104 9364 15156
rect 9496 15104 9548 15156
rect 9312 14968 9364 15020
rect 12440 15104 12492 15156
rect 10600 15036 10652 15088
rect 10968 15036 11020 15088
rect 1124 14900 1176 14952
rect 4804 14900 4856 14952
rect 5724 14900 5776 14952
rect 6092 14900 6144 14952
rect 6460 14900 6512 14952
rect 1860 14764 1912 14816
rect 5816 14764 5868 14816
rect 6092 14764 6144 14816
rect 7564 14832 7616 14884
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 8944 14900 8996 14952
rect 9680 14900 9732 14952
rect 11888 14968 11940 15020
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 14832 15104 14884 15156
rect 14188 15079 14240 15088
rect 10416 14900 10468 14952
rect 10968 14943 11020 14952
rect 10968 14909 10977 14943
rect 10977 14909 11011 14943
rect 11011 14909 11020 14943
rect 10968 14900 11020 14909
rect 14188 15045 14197 15079
rect 14197 15045 14231 15079
rect 14231 15045 14240 15079
rect 14188 15036 14240 15045
rect 14740 15036 14792 15088
rect 16856 15104 16908 15156
rect 16304 15036 16356 15088
rect 16580 15036 16632 15088
rect 16764 15036 16816 15088
rect 18328 15036 18380 15088
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 13820 14968 13872 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 18420 14968 18472 15020
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 22100 15104 22152 15156
rect 23572 15104 23624 15156
rect 23848 15104 23900 15156
rect 24952 15104 25004 15156
rect 27068 15147 27120 15156
rect 27068 15113 27077 15147
rect 27077 15113 27111 15147
rect 27111 15113 27120 15147
rect 27068 15104 27120 15113
rect 21548 15036 21600 15088
rect 21824 15036 21876 15088
rect 18880 14968 18932 14977
rect 19708 14968 19760 15020
rect 20996 14968 21048 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 23940 14968 23992 15020
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 7840 14764 7892 14816
rect 10508 14832 10560 14884
rect 10784 14832 10836 14884
rect 14280 14900 14332 14952
rect 14924 14900 14976 14952
rect 16396 14900 16448 14952
rect 20168 14900 20220 14952
rect 9588 14764 9640 14816
rect 9680 14764 9732 14816
rect 16304 14807 16356 14816
rect 16304 14773 16313 14807
rect 16313 14773 16347 14807
rect 16347 14773 16356 14807
rect 16304 14764 16356 14773
rect 17224 14832 17276 14884
rect 19984 14832 20036 14884
rect 26148 14900 26200 14952
rect 30564 14900 30616 14952
rect 18604 14764 18656 14816
rect 19156 14807 19208 14816
rect 19156 14773 19165 14807
rect 19165 14773 19199 14807
rect 19199 14773 19208 14807
rect 19156 14764 19208 14773
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 20536 14764 20588 14816
rect 21916 14832 21968 14884
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 5908 14560 5960 14612
rect 6092 14560 6144 14612
rect 1308 14424 1360 14476
rect 5448 14492 5500 14544
rect 7472 14492 7524 14544
rect 7656 14492 7708 14544
rect 7932 14492 7984 14544
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 9588 14560 9640 14612
rect 13360 14560 13412 14612
rect 13544 14560 13596 14612
rect 13820 14560 13872 14612
rect 14740 14560 14792 14612
rect 14924 14560 14976 14612
rect 26884 14560 26936 14612
rect 26976 14603 27028 14612
rect 26976 14569 26985 14603
rect 26985 14569 27019 14603
rect 27019 14569 27028 14603
rect 26976 14560 27028 14569
rect 4436 14424 4488 14476
rect 5816 14424 5868 14476
rect 6736 14424 6788 14476
rect 4252 14356 4304 14408
rect 2688 14288 2740 14340
rect 3516 14263 3568 14272
rect 3516 14229 3525 14263
rect 3525 14229 3559 14263
rect 3559 14229 3568 14263
rect 3516 14220 3568 14229
rect 4528 14220 4580 14272
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 5172 14356 5224 14408
rect 10784 14492 10836 14544
rect 21364 14492 21416 14544
rect 21732 14535 21784 14544
rect 21732 14501 21741 14535
rect 21741 14501 21775 14535
rect 21775 14501 21784 14535
rect 21732 14492 21784 14501
rect 23664 14492 23716 14544
rect 25780 14492 25832 14544
rect 9772 14424 9824 14476
rect 10140 14424 10192 14476
rect 10692 14424 10744 14476
rect 12808 14424 12860 14476
rect 15936 14424 15988 14476
rect 16304 14424 16356 14476
rect 17132 14424 17184 14476
rect 17592 14424 17644 14476
rect 19156 14424 19208 14476
rect 19800 14424 19852 14476
rect 5724 14331 5776 14340
rect 5724 14297 5733 14331
rect 5733 14297 5767 14331
rect 5767 14297 5776 14331
rect 5724 14288 5776 14297
rect 6276 14288 6328 14340
rect 7748 14288 7800 14340
rect 7380 14220 7432 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 8944 14220 8996 14272
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 9772 14220 9824 14229
rect 10876 14356 10928 14408
rect 11060 14356 11112 14408
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 14280 14356 14332 14408
rect 16580 14356 16632 14408
rect 10508 14220 10560 14272
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 10784 14220 10836 14272
rect 13912 14220 13964 14272
rect 15016 14220 15068 14272
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 17408 14288 17460 14340
rect 17592 14288 17644 14340
rect 22008 14424 22060 14476
rect 23940 14424 23992 14476
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 26608 14424 26660 14476
rect 19432 14288 19484 14340
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 21364 14220 21416 14272
rect 21916 14288 21968 14340
rect 23848 14288 23900 14340
rect 22652 14220 22704 14272
rect 22744 14220 22796 14272
rect 26976 14356 27028 14408
rect 25136 14288 25188 14340
rect 25872 14288 25924 14340
rect 26332 14288 26384 14340
rect 24584 14263 24636 14272
rect 24584 14229 24593 14263
rect 24593 14229 24627 14263
rect 24627 14229 24636 14263
rect 24584 14220 24636 14229
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 4712 14016 4764 14068
rect 6368 14016 6420 14068
rect 2320 13948 2372 14000
rect 5724 13991 5776 14000
rect 5724 13957 5733 13991
rect 5733 13957 5767 13991
rect 5767 13957 5776 13991
rect 5724 13948 5776 13957
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 9588 14016 9640 14068
rect 8576 13991 8628 14000
rect 8576 13957 8585 13991
rect 8585 13957 8619 13991
rect 8619 13957 8628 13991
rect 8576 13948 8628 13957
rect 11060 14016 11112 14068
rect 12072 14016 12124 14068
rect 14188 14016 14240 14068
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 16764 14016 16816 14068
rect 17316 14016 17368 14068
rect 20628 14016 20680 14068
rect 21088 14016 21140 14068
rect 25780 14016 25832 14068
rect 25872 14059 25924 14068
rect 25872 14025 25881 14059
rect 25881 14025 25915 14059
rect 25915 14025 25924 14059
rect 25872 14016 25924 14025
rect 26884 14016 26936 14068
rect 35072 14016 35124 14068
rect 1860 13880 1912 13932
rect 1308 13812 1360 13864
rect 4252 13880 4304 13932
rect 3424 13744 3476 13796
rect 4804 13812 4856 13864
rect 5264 13880 5316 13932
rect 14004 13948 14056 14000
rect 16580 13948 16632 14000
rect 21364 13948 21416 14000
rect 5724 13812 5776 13864
rect 6092 13812 6144 13864
rect 6644 13812 6696 13864
rect 5908 13744 5960 13796
rect 6460 13744 6512 13796
rect 7472 13855 7524 13864
rect 7472 13821 7481 13855
rect 7481 13821 7515 13855
rect 7515 13821 7524 13855
rect 7472 13812 7524 13821
rect 10876 13880 10928 13932
rect 11336 13880 11388 13932
rect 12072 13880 12124 13932
rect 7656 13744 7708 13796
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 10968 13812 11020 13864
rect 11520 13812 11572 13864
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 12256 13812 12308 13864
rect 15568 13880 15620 13932
rect 15752 13880 15804 13932
rect 16948 13880 17000 13932
rect 11244 13744 11296 13796
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 8760 13676 8812 13728
rect 10048 13676 10100 13728
rect 10140 13676 10192 13728
rect 14188 13744 14240 13796
rect 14464 13812 14516 13864
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 15200 13812 15252 13864
rect 15384 13812 15436 13864
rect 16120 13855 16172 13864
rect 16120 13821 16129 13855
rect 16129 13821 16163 13855
rect 16163 13821 16172 13855
rect 16120 13812 16172 13821
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17776 13812 17828 13864
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 21640 13880 21692 13932
rect 19984 13812 20036 13864
rect 22376 13880 22428 13932
rect 23848 13991 23900 14000
rect 23848 13957 23857 13991
rect 23857 13957 23891 13991
rect 23891 13957 23900 13991
rect 23848 13948 23900 13957
rect 24584 13948 24636 14000
rect 25136 13948 25188 14000
rect 22652 13855 22704 13864
rect 20720 13744 20772 13796
rect 13360 13676 13412 13728
rect 14648 13676 14700 13728
rect 17500 13676 17552 13728
rect 20168 13676 20220 13728
rect 22652 13821 22661 13855
rect 22661 13821 22695 13855
rect 22695 13821 22704 13855
rect 22652 13812 22704 13821
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 23756 13812 23808 13864
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 25136 13812 25188 13864
rect 20996 13676 21048 13728
rect 22560 13676 22612 13728
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 4436 13515 4488 13524
rect 4436 13481 4466 13515
rect 4466 13481 4488 13515
rect 4436 13472 4488 13481
rect 7104 13472 7156 13524
rect 10140 13472 10192 13524
rect 11152 13472 11204 13524
rect 5448 13404 5500 13456
rect 6000 13404 6052 13456
rect 8576 13404 8628 13456
rect 12440 13472 12492 13524
rect 12808 13472 12860 13524
rect 13820 13472 13872 13524
rect 17408 13515 17460 13524
rect 17408 13481 17432 13515
rect 17432 13481 17460 13515
rect 17408 13472 17460 13481
rect 17500 13472 17552 13524
rect 19156 13472 19208 13524
rect 19524 13472 19576 13524
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 5172 13336 5224 13388
rect 7380 13336 7432 13388
rect 1952 13268 2004 13320
rect 3884 13311 3936 13320
rect 3884 13277 3893 13311
rect 3893 13277 3927 13311
rect 3927 13277 3936 13311
rect 3884 13268 3936 13277
rect 1860 13200 1912 13252
rect 4712 13200 4764 13252
rect 2596 13132 2648 13184
rect 3424 13132 3476 13184
rect 4804 13132 4856 13184
rect 6276 13268 6328 13320
rect 5816 13200 5868 13252
rect 6000 13200 6052 13252
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6368 13132 6420 13184
rect 6552 13132 6604 13184
rect 7288 13200 7340 13252
rect 7472 13200 7524 13252
rect 7656 13132 7708 13184
rect 11244 13336 11296 13388
rect 11520 13336 11572 13388
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 13268 13336 13320 13388
rect 15200 13336 15252 13388
rect 16396 13336 16448 13388
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 17132 13379 17184 13388
rect 17132 13345 17141 13379
rect 17141 13345 17175 13379
rect 17175 13345 17184 13379
rect 17132 13336 17184 13345
rect 17500 13336 17552 13388
rect 17868 13336 17920 13388
rect 20996 13472 21048 13524
rect 21824 13472 21876 13524
rect 22376 13472 22428 13524
rect 23296 13472 23348 13524
rect 21640 13404 21692 13456
rect 22192 13336 22244 13388
rect 23388 13404 23440 13456
rect 23848 13404 23900 13456
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23480 13336 23532 13345
rect 23572 13336 23624 13388
rect 32496 13336 32548 13388
rect 9404 13311 9456 13320
rect 9404 13277 9413 13311
rect 9413 13277 9447 13311
rect 9447 13277 9456 13311
rect 9404 13268 9456 13277
rect 11704 13268 11756 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 19156 13268 19208 13320
rect 19524 13268 19576 13320
rect 23020 13268 23072 13320
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 12348 13200 12400 13252
rect 13912 13200 13964 13252
rect 15844 13200 15896 13252
rect 16580 13200 16632 13252
rect 13636 13132 13688 13184
rect 14004 13132 14056 13184
rect 14372 13132 14424 13184
rect 16120 13132 16172 13184
rect 18972 13200 19024 13252
rect 21180 13200 21232 13252
rect 20352 13132 20404 13184
rect 23112 13132 23164 13184
rect 23388 13200 23440 13252
rect 26884 13200 26936 13252
rect 25228 13132 25280 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 5540 12928 5592 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 6644 12928 6696 12980
rect 10600 12928 10652 12980
rect 11796 12928 11848 12980
rect 13452 12928 13504 12980
rect 13636 12928 13688 12980
rect 13728 12971 13780 12980
rect 13728 12937 13737 12971
rect 13737 12937 13771 12971
rect 13771 12937 13780 12971
rect 13728 12928 13780 12937
rect 14464 12928 14516 12980
rect 15292 12928 15344 12980
rect 16580 12928 16632 12980
rect 16948 12928 17000 12980
rect 20168 12928 20220 12980
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 21180 12928 21232 12980
rect 23112 12928 23164 12980
rect 23480 12928 23532 12980
rect 4344 12860 4396 12912
rect 4620 12860 4672 12912
rect 4712 12860 4764 12912
rect 5448 12860 5500 12912
rect 5816 12860 5868 12912
rect 6276 12860 6328 12912
rect 2504 12792 2556 12844
rect 3608 12792 3660 12844
rect 4068 12792 4120 12844
rect 1216 12724 1268 12776
rect 3332 12724 3384 12776
rect 6828 12792 6880 12844
rect 4252 12724 4304 12776
rect 4804 12724 4856 12776
rect 6000 12724 6052 12776
rect 2044 12656 2096 12708
rect 8576 12860 8628 12912
rect 8760 12860 8812 12912
rect 13176 12860 13228 12912
rect 13360 12860 13412 12912
rect 14280 12860 14332 12912
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 3516 12588 3568 12640
rect 5632 12588 5684 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7380 12588 7432 12640
rect 9036 12724 9088 12776
rect 9956 12724 10008 12776
rect 10140 12724 10192 12776
rect 13452 12792 13504 12844
rect 10508 12699 10560 12708
rect 10508 12665 10517 12699
rect 10517 12665 10551 12699
rect 10551 12665 10560 12699
rect 10508 12656 10560 12665
rect 10784 12656 10836 12708
rect 12624 12656 12676 12708
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 13820 12724 13872 12776
rect 14832 12792 14884 12844
rect 15108 12792 15160 12844
rect 18880 12860 18932 12912
rect 20628 12860 20680 12912
rect 23572 12860 23624 12912
rect 23940 12860 23992 12912
rect 17408 12792 17460 12844
rect 17960 12792 18012 12844
rect 15200 12724 15252 12776
rect 16856 12767 16908 12776
rect 16856 12733 16865 12767
rect 16865 12733 16899 12767
rect 16899 12733 16908 12767
rect 16856 12724 16908 12733
rect 18604 12724 18656 12776
rect 17224 12656 17276 12708
rect 17500 12656 17552 12708
rect 20076 12724 20128 12776
rect 22100 12792 22152 12844
rect 22192 12792 22244 12844
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 21456 12724 21508 12776
rect 23664 12724 23716 12776
rect 23940 12724 23992 12776
rect 24492 12724 24544 12776
rect 22468 12656 22520 12708
rect 9312 12588 9364 12640
rect 10048 12588 10100 12640
rect 10324 12588 10376 12640
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 11428 12588 11480 12640
rect 12256 12588 12308 12640
rect 13452 12588 13504 12640
rect 14004 12588 14056 12640
rect 14188 12588 14240 12640
rect 14648 12588 14700 12640
rect 16856 12588 16908 12640
rect 19432 12588 19484 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 4344 12384 4396 12436
rect 3516 12316 3568 12368
rect 4252 12248 4304 12300
rect 940 12180 992 12232
rect 1492 12180 1544 12232
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 7196 12384 7248 12436
rect 10876 12384 10928 12436
rect 12532 12384 12584 12436
rect 12624 12384 12676 12436
rect 13912 12384 13964 12436
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 7288 12316 7340 12368
rect 5172 12248 5224 12300
rect 7564 12248 7616 12300
rect 8944 12316 8996 12368
rect 9404 12316 9456 12368
rect 11336 12316 11388 12368
rect 9312 12248 9364 12300
rect 12072 12248 12124 12300
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 4804 12180 4856 12232
rect 9680 12180 9732 12232
rect 12624 12180 12676 12232
rect 2780 12112 2832 12164
rect 5080 12112 5132 12164
rect 5724 12112 5776 12164
rect 6276 12112 6328 12164
rect 9128 12155 9180 12164
rect 9128 12121 9137 12155
rect 9137 12121 9171 12155
rect 9171 12121 9180 12155
rect 9128 12112 9180 12121
rect 9772 12112 9824 12164
rect 11152 12112 11204 12164
rect 13268 12316 13320 12368
rect 15200 12384 15252 12436
rect 17960 12384 18012 12436
rect 18144 12384 18196 12436
rect 19156 12384 19208 12436
rect 20720 12384 20772 12436
rect 18880 12359 18932 12368
rect 18880 12325 18889 12359
rect 18889 12325 18923 12359
rect 18923 12325 18932 12359
rect 18880 12316 18932 12325
rect 14648 12248 14700 12300
rect 14832 12248 14884 12300
rect 16580 12291 16632 12300
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 17316 12248 17368 12300
rect 14924 12180 14976 12232
rect 18144 12180 18196 12232
rect 3792 12044 3844 12096
rect 4344 12044 4396 12096
rect 7564 12044 7616 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 11888 12044 11940 12096
rect 13176 12044 13228 12096
rect 13912 12044 13964 12096
rect 14832 12044 14884 12096
rect 16212 12044 16264 12096
rect 19708 12112 19760 12164
rect 18420 12044 18472 12096
rect 18880 12044 18932 12096
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 24492 12427 24544 12436
rect 24492 12393 24501 12427
rect 24501 12393 24535 12427
rect 24535 12393 24544 12427
rect 24492 12384 24544 12393
rect 22192 12180 22244 12232
rect 23940 12180 23992 12232
rect 20352 12155 20404 12164
rect 20352 12121 20361 12155
rect 20361 12121 20395 12155
rect 20395 12121 20404 12155
rect 20352 12112 20404 12121
rect 21088 12112 21140 12164
rect 25044 12112 25096 12164
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 1768 11883 1820 11892
rect 1768 11849 1777 11883
rect 1777 11849 1811 11883
rect 1811 11849 1820 11883
rect 1768 11840 1820 11849
rect 3516 11840 3568 11892
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 6460 11883 6512 11892
rect 6460 11849 6469 11883
rect 6469 11849 6503 11883
rect 6503 11849 6512 11883
rect 6460 11840 6512 11849
rect 4160 11772 4212 11824
rect 6828 11772 6880 11824
rect 7656 11815 7708 11824
rect 7656 11781 7665 11815
rect 7665 11781 7699 11815
rect 7699 11781 7708 11815
rect 7656 11772 7708 11781
rect 8116 11772 8168 11824
rect 9312 11772 9364 11824
rect 9496 11772 9548 11824
rect 9956 11772 10008 11824
rect 10600 11772 10652 11824
rect 1952 11704 2004 11756
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 5264 11704 5316 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 9128 11704 9180 11756
rect 11336 11704 11388 11756
rect 14096 11840 14148 11892
rect 14372 11840 14424 11892
rect 13360 11772 13412 11824
rect 14832 11772 14884 11824
rect 15844 11772 15896 11824
rect 18696 11840 18748 11892
rect 1952 11568 2004 11620
rect 5632 11636 5684 11688
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 4896 11568 4948 11620
rect 5540 11568 5592 11620
rect 4988 11500 5040 11552
rect 7840 11500 7892 11552
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 18420 11772 18472 11824
rect 18788 11772 18840 11824
rect 24032 11840 24084 11892
rect 22744 11772 22796 11824
rect 23940 11772 23992 11824
rect 19432 11704 19484 11756
rect 9036 11568 9088 11620
rect 11520 11568 11572 11620
rect 11796 11568 11848 11620
rect 14188 11636 14240 11688
rect 17040 11636 17092 11688
rect 17592 11679 17644 11688
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 17592 11636 17644 11645
rect 17776 11636 17828 11688
rect 19708 11679 19760 11688
rect 19708 11645 19717 11679
rect 19717 11645 19751 11679
rect 19751 11645 19760 11679
rect 19708 11636 19760 11645
rect 21180 11636 21232 11688
rect 22192 11636 22244 11688
rect 12624 11568 12676 11620
rect 13176 11568 13228 11620
rect 15292 11568 15344 11620
rect 17224 11568 17276 11620
rect 8760 11500 8812 11552
rect 10232 11500 10284 11552
rect 11152 11500 11204 11552
rect 12072 11500 12124 11552
rect 19156 11500 19208 11552
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 23388 11500 23440 11552
rect 25136 11500 25188 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 3700 11296 3752 11348
rect 5632 11296 5684 11348
rect 5724 11296 5776 11348
rect 7472 11339 7524 11348
rect 7472 11305 7481 11339
rect 7481 11305 7515 11339
rect 7515 11305 7524 11339
rect 7472 11296 7524 11305
rect 10600 11296 10652 11348
rect 11612 11296 11664 11348
rect 12256 11296 12308 11348
rect 12348 11296 12400 11348
rect 13360 11296 13412 11348
rect 13452 11296 13504 11348
rect 13912 11296 13964 11348
rect 16580 11296 16632 11348
rect 17408 11296 17460 11348
rect 18604 11296 18656 11348
rect 18972 11296 19024 11348
rect 22836 11296 22888 11348
rect 2596 11160 2648 11212
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 7104 11228 7156 11280
rect 5540 11160 5592 11212
rect 5632 11160 5684 11212
rect 7288 11160 7340 11212
rect 7932 11160 7984 11212
rect 9036 11228 9088 11280
rect 9588 11203 9640 11212
rect 9588 11169 9597 11203
rect 9597 11169 9631 11203
rect 9631 11169 9640 11203
rect 9588 11160 9640 11169
rect 11336 11228 11388 11280
rect 1584 11024 1636 11076
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 6460 11092 6512 11144
rect 7472 11092 7524 11144
rect 8116 11092 8168 11144
rect 9220 11092 9272 11144
rect 10416 11092 10468 11144
rect 8760 11024 8812 11076
rect 9404 11024 9456 11076
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 13360 11160 13412 11212
rect 21548 11160 21600 11212
rect 13912 11024 13964 11076
rect 14556 11024 14608 11076
rect 16856 11092 16908 11144
rect 18880 11092 18932 11144
rect 14924 11024 14976 11076
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 9588 10956 9640 11008
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 15844 10956 15896 11008
rect 16488 11024 16540 11076
rect 17408 11067 17460 11076
rect 17408 11033 17417 11067
rect 17417 11033 17451 11067
rect 17451 11033 17460 11067
rect 17408 11024 17460 11033
rect 17868 11024 17920 11076
rect 19708 11024 19760 11076
rect 22284 11092 22336 11144
rect 23572 11296 23624 11348
rect 23940 11296 23992 11348
rect 31852 11296 31904 11348
rect 26884 11160 26936 11212
rect 31852 11092 31904 11144
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 27620 11024 27672 11076
rect 31300 11024 31352 11076
rect 47860 11024 47912 11076
rect 18696 10956 18748 11008
rect 21364 10956 21416 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 4436 10752 4488 10804
rect 2596 10684 2648 10736
rect 6736 10684 6788 10736
rect 8300 10684 8352 10736
rect 13820 10752 13872 10804
rect 15292 10752 15344 10804
rect 15384 10752 15436 10804
rect 17040 10752 17092 10804
rect 11152 10684 11204 10736
rect 11980 10684 12032 10736
rect 12072 10684 12124 10736
rect 13912 10684 13964 10736
rect 16764 10684 16816 10736
rect 5080 10616 5132 10668
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 5632 10616 5684 10668
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 10324 10616 10376 10668
rect 1032 10480 1084 10532
rect 6920 10548 6972 10600
rect 2596 10480 2648 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 1952 10412 2004 10464
rect 3792 10412 3844 10464
rect 7380 10480 7432 10532
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 6736 10412 6788 10464
rect 6920 10412 6972 10464
rect 7472 10412 7524 10464
rect 8116 10548 8168 10600
rect 10692 10548 10744 10600
rect 10968 10616 11020 10668
rect 11244 10548 11296 10600
rect 15384 10616 15436 10668
rect 10232 10480 10284 10532
rect 15200 10548 15252 10600
rect 7840 10412 7892 10464
rect 8208 10412 8260 10464
rect 11520 10412 11572 10464
rect 11796 10412 11848 10464
rect 16028 10412 16080 10464
rect 16304 10548 16356 10600
rect 16580 10548 16632 10600
rect 17868 10684 17920 10736
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 21456 10752 21508 10804
rect 21548 10684 21600 10736
rect 22284 10752 22336 10804
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 22836 10548 22888 10600
rect 21364 10480 21416 10532
rect 20536 10412 20588 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 1216 10208 1268 10260
rect 2872 10208 2924 10260
rect 3608 10208 3660 10260
rect 4436 10208 4488 10260
rect 6644 10208 6696 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 10784 10208 10836 10260
rect 10968 10208 11020 10260
rect 12164 10208 12216 10260
rect 13912 10208 13964 10260
rect 15016 10208 15068 10260
rect 17776 10208 17828 10260
rect 18880 10251 18932 10260
rect 18880 10217 18889 10251
rect 18889 10217 18923 10251
rect 18923 10217 18932 10251
rect 18880 10208 18932 10217
rect 19800 10208 19852 10260
rect 21548 10251 21600 10260
rect 21548 10217 21557 10251
rect 21557 10217 21591 10251
rect 21591 10217 21600 10251
rect 21548 10208 21600 10217
rect 1676 10072 1728 10124
rect 3424 10140 3476 10192
rect 6460 10183 6512 10192
rect 6460 10149 6469 10183
rect 6469 10149 6503 10183
rect 6503 10149 6512 10183
rect 6460 10140 6512 10149
rect 8116 10140 8168 10192
rect 10876 10140 10928 10192
rect 3516 10072 3568 10124
rect 4252 10115 4304 10124
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 4804 10072 4856 10124
rect 7840 10072 7892 10124
rect 2688 10004 2740 10056
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 8300 10072 8352 10124
rect 9036 10072 9088 10124
rect 11980 10072 12032 10124
rect 10968 10004 11020 10056
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 12624 10004 12676 10056
rect 4620 9936 4672 9988
rect 7104 9979 7156 9988
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 7380 9936 7432 9988
rect 11796 9936 11848 9988
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 15200 10072 15252 10124
rect 16212 10072 16264 10124
rect 16856 10004 16908 10056
rect 19708 10072 19760 10124
rect 20720 10004 20772 10056
rect 21548 10004 21600 10056
rect 13912 9936 13964 9988
rect 2412 9868 2464 9920
rect 3792 9868 3844 9920
rect 8392 9868 8444 9920
rect 11428 9868 11480 9920
rect 11888 9868 11940 9920
rect 15200 9868 15252 9920
rect 17040 9936 17092 9988
rect 19248 9936 19300 9988
rect 23388 9936 23440 9988
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 6460 9707 6512 9716
rect 6460 9673 6469 9707
rect 6469 9673 6503 9707
rect 6503 9673 6512 9707
rect 6460 9664 6512 9673
rect 7656 9664 7708 9716
rect 15476 9664 15528 9716
rect 16212 9707 16264 9716
rect 16212 9673 16221 9707
rect 16221 9673 16255 9707
rect 16255 9673 16264 9707
rect 16212 9664 16264 9673
rect 1492 9639 1544 9648
rect 1492 9605 1501 9639
rect 1501 9605 1535 9639
rect 1535 9605 1544 9639
rect 1492 9596 1544 9605
rect 1768 9596 1820 9648
rect 3240 9639 3292 9648
rect 3240 9605 3249 9639
rect 3249 9605 3283 9639
rect 3283 9605 3292 9639
rect 3240 9596 3292 9605
rect 5908 9596 5960 9648
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 5172 9528 5224 9580
rect 5448 9528 5500 9580
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2320 9460 2372 9512
rect 3608 9435 3660 9444
rect 3608 9401 3617 9435
rect 3617 9401 3651 9435
rect 3651 9401 3660 9435
rect 3608 9392 3660 9401
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 8484 9596 8536 9648
rect 9036 9596 9088 9648
rect 10600 9596 10652 9648
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 12624 9596 12676 9648
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 15200 9596 15252 9648
rect 16028 9596 16080 9648
rect 18880 9664 18932 9716
rect 18512 9596 18564 9648
rect 24584 9596 24636 9648
rect 27804 9596 27856 9648
rect 31300 9596 31352 9648
rect 9680 9528 9732 9580
rect 7840 9460 7892 9512
rect 10324 9460 10376 9512
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 11244 9460 11296 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 15292 9460 15344 9512
rect 16764 9460 16816 9512
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17224 9460 17276 9512
rect 23756 9528 23808 9580
rect 21180 9460 21232 9512
rect 23388 9460 23440 9512
rect 13360 9392 13412 9444
rect 5632 9324 5684 9376
rect 7380 9324 7432 9376
rect 8116 9324 8168 9376
rect 11428 9324 11480 9376
rect 12440 9324 12492 9376
rect 13544 9324 13596 9376
rect 18512 9392 18564 9444
rect 14004 9324 14056 9376
rect 15752 9324 15804 9376
rect 16304 9324 16356 9376
rect 19064 9435 19116 9444
rect 19064 9401 19073 9435
rect 19073 9401 19107 9435
rect 19107 9401 19116 9435
rect 19064 9392 19116 9401
rect 20720 9324 20772 9376
rect 27804 9367 27856 9376
rect 27804 9333 27813 9367
rect 27813 9333 27847 9367
rect 27847 9333 27856 9367
rect 27804 9324 27856 9333
rect 31576 9324 31628 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 3792 9120 3844 9172
rect 4068 9052 4120 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 5264 9120 5316 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 9680 9120 9732 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 32404 9120 32456 9172
rect 4896 9052 4948 9104
rect 2872 8916 2924 8968
rect 3424 8916 3476 8968
rect 4252 8916 4304 8968
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 6828 9052 6880 9104
rect 13636 9052 13688 9104
rect 15936 9052 15988 9104
rect 3240 8848 3292 8900
rect 4712 8848 4764 8900
rect 7748 8916 7800 8968
rect 8116 8984 8168 9036
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 8668 8916 8720 8968
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 13544 8984 13596 9036
rect 15292 8984 15344 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 15844 8984 15896 9036
rect 16856 8984 16908 9036
rect 15016 8916 15068 8968
rect 9128 8848 9180 8900
rect 11888 8848 11940 8900
rect 7656 8780 7708 8832
rect 8208 8823 8260 8832
rect 8208 8789 8217 8823
rect 8217 8789 8251 8823
rect 8251 8789 8260 8823
rect 8208 8780 8260 8789
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 9680 8780 9732 8832
rect 11244 8780 11296 8832
rect 11612 8780 11664 8832
rect 12440 8780 12492 8832
rect 16304 8891 16356 8900
rect 16304 8857 16313 8891
rect 16313 8857 16347 8891
rect 16347 8857 16356 8891
rect 16304 8848 16356 8857
rect 14740 8780 14792 8832
rect 17592 8780 17644 8832
rect 18512 8780 18564 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 3332 8576 3384 8628
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 5080 8576 5132 8628
rect 6460 8619 6512 8628
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 6460 8576 6512 8585
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 7748 8576 7800 8628
rect 8116 8576 8168 8628
rect 1124 8508 1176 8560
rect 1400 8440 1452 8492
rect 3700 8440 3752 8492
rect 4252 8440 4304 8492
rect 10048 8508 10100 8560
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 14004 8576 14056 8628
rect 15384 8576 15436 8628
rect 11244 8508 11296 8560
rect 1308 8372 1360 8424
rect 3332 8372 3384 8424
rect 7012 8372 7064 8424
rect 6920 8304 6972 8356
rect 7564 8440 7616 8492
rect 8116 8372 8168 8424
rect 8760 8440 8812 8492
rect 9036 8440 9088 8492
rect 10416 8440 10468 8492
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 9864 8347 9916 8356
rect 2228 8236 2280 8288
rect 4436 8236 4488 8288
rect 7472 8236 7524 8288
rect 9864 8313 9873 8347
rect 9873 8313 9907 8347
rect 9907 8313 9916 8347
rect 9864 8304 9916 8313
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 14740 8508 14792 8560
rect 12440 8440 12492 8492
rect 16580 8576 16632 8628
rect 15844 8508 15896 8560
rect 20444 8440 20496 8492
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 12532 8304 12584 8356
rect 14188 8372 14240 8424
rect 16028 8372 16080 8424
rect 20352 8372 20404 8424
rect 16488 8304 16540 8356
rect 8484 8236 8536 8288
rect 10232 8236 10284 8288
rect 12808 8236 12860 8288
rect 16396 8236 16448 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 1952 8032 2004 8084
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 3792 8032 3844 8084
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 8300 8032 8352 8084
rect 2596 7964 2648 8016
rect 6736 7964 6788 8016
rect 2228 7896 2280 7948
rect 2596 7828 2648 7880
rect 2872 7828 2924 7880
rect 7288 7896 7340 7948
rect 10324 7896 10376 7948
rect 8576 7828 8628 7880
rect 11060 7828 11112 7880
rect 12808 8032 12860 8084
rect 17224 8032 17276 8084
rect 15200 8007 15252 8016
rect 15200 7973 15209 8007
rect 15209 7973 15243 8007
rect 15243 7973 15252 8007
rect 15200 7964 15252 7973
rect 14188 7871 14240 7880
rect 3332 7760 3384 7812
rect 3240 7692 3292 7744
rect 6828 7760 6880 7812
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 19248 7896 19300 7948
rect 12072 7760 12124 7812
rect 3700 7692 3752 7744
rect 5632 7692 5684 7744
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 22836 7692 22888 7744
rect 23388 7692 23440 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 1676 7488 1728 7540
rect 4068 7488 4120 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 1308 7284 1360 7336
rect 3332 7352 3384 7404
rect 3792 7420 3844 7472
rect 11704 7488 11756 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 13360 7488 13412 7540
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 27620 7488 27672 7540
rect 9588 7420 9640 7472
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 11428 7420 11480 7472
rect 2688 7284 2740 7336
rect 4988 7284 5040 7336
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 23572 7352 23624 7404
rect 22468 7327 22520 7336
rect 22468 7293 22477 7327
rect 22477 7293 22511 7327
rect 22511 7293 22520 7327
rect 22468 7284 22520 7293
rect 2228 7259 2280 7268
rect 2228 7225 2237 7259
rect 2237 7225 2271 7259
rect 2271 7225 2280 7259
rect 2228 7216 2280 7225
rect 8392 7216 8444 7268
rect 6368 7148 6420 7200
rect 12440 7148 12492 7200
rect 14004 7148 14056 7200
rect 17500 7148 17552 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 3424 6987 3476 6996
rect 3424 6953 3433 6987
rect 3433 6953 3467 6987
rect 3467 6953 3476 6987
rect 3424 6944 3476 6953
rect 23940 6944 23992 6996
rect 1308 6808 1360 6860
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2596 6740 2648 6792
rect 2780 6740 2832 6792
rect 3332 6808 3384 6860
rect 23756 6919 23808 6928
rect 23756 6885 23765 6919
rect 23765 6885 23799 6919
rect 23799 6885 23808 6919
rect 23756 6876 23808 6885
rect 9772 6808 9824 6860
rect 10508 6808 10560 6860
rect 19340 6808 19392 6860
rect 20720 6808 20772 6860
rect 21732 6740 21784 6792
rect 2136 6604 2188 6656
rect 7104 6672 7156 6724
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 23388 6647 23440 6656
rect 23388 6613 23397 6647
rect 23397 6613 23431 6647
rect 23431 6613 23440 6647
rect 23388 6604 23440 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 4344 6400 4396 6452
rect 22836 6443 22888 6452
rect 22836 6409 22845 6443
rect 22845 6409 22879 6443
rect 22879 6409 22888 6443
rect 22836 6400 22888 6409
rect 1768 6332 1820 6384
rect 3976 6332 4028 6384
rect 2872 6264 2924 6316
rect 1308 6196 1360 6248
rect 12256 6196 12308 6248
rect 22744 6060 22796 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 1308 5856 1360 5908
rect 22468 5856 22520 5908
rect 7564 5788 7616 5840
rect 12624 5788 12676 5840
rect 21732 5831 21784 5840
rect 21732 5797 21741 5831
rect 21741 5797 21775 5831
rect 21775 5797 21784 5831
rect 21732 5788 21784 5797
rect 6000 5720 6052 5772
rect 14004 5720 14056 5772
rect 16856 5720 16908 5772
rect 1308 5652 1360 5704
rect 12624 5652 12676 5704
rect 17040 5516 17092 5568
rect 18512 5652 18564 5704
rect 20260 5652 20312 5704
rect 22744 5720 22796 5772
rect 28724 5720 28776 5772
rect 28908 5720 28960 5772
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 22192 5584 22244 5636
rect 23388 5584 23440 5636
rect 25504 5584 25556 5636
rect 21364 5559 21416 5568
rect 21364 5525 21373 5559
rect 21373 5525 21407 5559
rect 21407 5525 21416 5559
rect 21364 5516 21416 5525
rect 27160 5627 27212 5636
rect 27160 5593 27169 5627
rect 27169 5593 27203 5627
rect 27203 5593 27212 5627
rect 27160 5584 27212 5593
rect 27620 5516 27672 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 27160 5312 27212 5364
rect 28356 5244 28408 5296
rect 1308 5176 1360 5228
rect 12440 5176 12492 5228
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 9404 5108 9456 5160
rect 15476 5108 15528 5160
rect 21364 5176 21416 5228
rect 22192 5219 22244 5228
rect 22192 5185 22210 5219
rect 22210 5185 22244 5219
rect 22192 5176 22244 5185
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 28816 5151 28868 5160
rect 28816 5117 28825 5151
rect 28825 5117 28859 5151
rect 28859 5117 28868 5151
rect 28816 5108 28868 5117
rect 41420 5108 41472 5160
rect 33508 5040 33560 5092
rect 17868 4972 17920 5024
rect 20536 4972 20588 5024
rect 25964 4972 26016 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 17408 4768 17460 4820
rect 20260 4811 20312 4820
rect 20260 4777 20269 4811
rect 20269 4777 20303 4811
rect 20303 4777 20312 4811
rect 20260 4768 20312 4777
rect 28816 4768 28868 4820
rect 1308 4632 1360 4684
rect 9956 4632 10008 4684
rect 27804 4632 27856 4684
rect 20260 4564 20312 4616
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 17684 4428 17736 4480
rect 27252 4564 27304 4616
rect 25964 4539 26016 4548
rect 25964 4505 25973 4539
rect 25973 4505 26007 4539
rect 26007 4505 26016 4539
rect 25964 4496 26016 4505
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1216 4088 1268 4140
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 2780 4088 2832 4140
rect 1308 4020 1360 4072
rect 6828 4088 6880 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 1768 3884 1820 3936
rect 10600 3884 10652 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 1584 3680 1636 3732
rect 9680 3680 9732 3732
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 1308 3476 1360 3528
rect 28908 3612 28960 3664
rect 44088 3612 44140 3664
rect 2044 3544 2096 3596
rect 27252 3544 27304 3596
rect 46756 3544 46808 3596
rect 2872 3476 2924 3528
rect 12072 3408 12124 3460
rect 27620 3476 27672 3528
rect 49424 3476 49476 3528
rect 13452 3408 13504 3460
rect 20720 3408 20772 3460
rect 38752 3408 38804 3460
rect 3424 3340 3476 3392
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 9772 3136 9824 3188
rect 10416 3068 10468 3120
rect 12624 3111 12676 3120
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 15476 3068 15528 3120
rect 17684 3068 17736 3120
rect 1400 3000 1452 3052
rect 3332 3000 3384 3052
rect 1308 2932 1360 2984
rect 2412 2932 2464 2984
rect 7840 3000 7892 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17868 3000 17920 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 3792 2864 3844 2916
rect 17408 2932 17460 2984
rect 8300 2796 8352 2848
rect 12440 2864 12492 2916
rect 17500 2796 17552 2848
rect 20076 2796 20128 2848
rect 22008 2796 22060 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 7564 2592 7616 2644
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 27804 2592 27856 2644
rect 28724 2592 28776 2644
rect 33508 2635 33560 2644
rect 33508 2601 33517 2635
rect 33517 2601 33551 2635
rect 33551 2601 33560 2635
rect 33508 2592 33560 2601
rect 1216 2456 1268 2508
rect 3424 2456 3476 2508
rect 4068 2456 4120 2508
rect 11612 2524 11664 2576
rect 6736 2456 6788 2508
rect 9404 2456 9456 2508
rect 12072 2456 12124 2508
rect 14740 2456 14792 2508
rect 17408 2456 17460 2508
rect 20168 2456 20220 2508
rect 22744 2456 22796 2508
rect 31576 2456 31628 2508
rect 1308 2320 1360 2372
rect 8300 2388 8352 2440
rect 9772 2388 9824 2440
rect 12440 2388 12492 2440
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 22008 2388 22060 2440
rect 25412 2388 25464 2440
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 30748 2388 30800 2440
rect 33416 2388 33468 2440
rect 36084 2431 36136 2440
rect 36084 2397 36093 2431
rect 36093 2397 36127 2431
rect 36127 2397 36136 2431
rect 36084 2388 36136 2397
rect 6552 2252 6604 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 2226 26200 2282 27000
rect 2870 26330 2926 27000
rect 2870 26302 3372 26330
rect 2870 26200 2926 26302
rect 1768 24132 1820 24138
rect 1768 24074 1820 24080
rect 1780 23610 1808 24074
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 1216 23588 1268 23594
rect 1216 23530 1268 23536
rect 1688 23582 1808 23610
rect 1032 22772 1084 22778
rect 1032 22714 1084 22720
rect 940 17604 992 17610
rect 940 17546 992 17552
rect 952 17105 980 17546
rect 938 17096 994 17105
rect 938 17031 994 17040
rect 940 12232 992 12238
rect 938 12200 940 12209
rect 992 12200 994 12209
rect 938 12135 994 12144
rect 1044 10538 1072 22714
rect 1124 17128 1176 17134
rect 1124 17070 1176 17076
rect 1136 16697 1164 17070
rect 1122 16688 1178 16697
rect 1228 16674 1256 23530
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1504 19417 1532 23151
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17921 1440 18770
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 1490 16688 1546 16697
rect 1228 16646 1348 16674
rect 1122 16623 1178 16632
rect 1216 16516 1268 16522
rect 1216 16458 1268 16464
rect 1228 16289 1256 16458
rect 1214 16280 1270 16289
rect 1214 16215 1270 16224
rect 1124 16040 1176 16046
rect 1124 15982 1176 15988
rect 1136 15881 1164 15982
rect 1122 15872 1178 15881
rect 1122 15807 1178 15816
rect 1320 15688 1348 16646
rect 1490 16623 1546 16632
rect 1504 16574 1532 16623
rect 1504 16546 1624 16574
rect 1228 15660 1348 15688
rect 1122 15056 1178 15065
rect 1122 14991 1178 15000
rect 1136 14958 1164 14991
rect 1124 14952 1176 14958
rect 1124 14894 1176 14900
rect 1228 14770 1256 15660
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1136 14742 1256 14770
rect 1032 10532 1084 10538
rect 1032 10474 1084 10480
rect 1136 8566 1164 14742
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1214 13424 1270 13433
rect 1214 13359 1270 13368
rect 1228 12782 1256 13359
rect 1216 12776 1268 12782
rect 1216 12718 1268 12724
rect 1228 10266 1256 12718
rect 1596 12434 1624 16546
rect 1412 12406 1624 12434
rect 1306 10976 1362 10985
rect 1306 10911 1362 10920
rect 1216 10260 1268 10266
rect 1216 10202 1268 10208
rect 1124 8560 1176 8566
rect 1124 8502 1176 8508
rect 1320 8430 1348 10911
rect 1412 8498 1440 12406
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1504 9654 1532 12174
rect 1688 12152 1716 23582
rect 1768 23520 1820 23526
rect 2148 23497 2176 23666
rect 1768 23462 1820 23468
rect 2134 23488 2190 23497
rect 1780 20466 1808 23462
rect 2134 23423 2190 23432
rect 2240 22234 2268 26200
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2778 24440 2834 24449
rect 2950 24443 3258 24452
rect 2778 24375 2780 24384
rect 2832 24375 2834 24384
rect 2780 24346 2832 24352
rect 2412 24200 2464 24206
rect 2412 24142 2464 24148
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2136 21344 2188 21350
rect 2136 21286 2188 21292
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1766 19816 1822 19825
rect 1766 19751 1822 19760
rect 1596 12124 1716 12152
rect 1596 11082 1624 12124
rect 1780 12050 1808 19751
rect 1872 17814 1900 20878
rect 2148 19378 2176 21286
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 2056 17513 2084 18158
rect 2136 17536 2188 17542
rect 2042 17504 2098 17513
rect 2136 17478 2188 17484
rect 2042 17439 2098 17448
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1872 14822 1900 16050
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1858 13968 1914 13977
rect 1858 13903 1860 13912
rect 1912 13903 1914 13912
rect 1860 13874 1912 13880
rect 2042 13832 2098 13841
rect 2042 13767 2098 13776
rect 1950 13424 2006 13433
rect 2056 13394 2084 13767
rect 1950 13359 2006 13368
rect 2044 13388 2096 13394
rect 1964 13326 1992 13359
rect 2044 13330 2096 13336
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1688 12022 1808 12050
rect 1688 11778 1716 12022
rect 1766 11928 1822 11937
rect 1766 11863 1768 11872
rect 1820 11863 1822 11872
rect 1768 11834 1820 11840
rect 1688 11750 1808 11778
rect 1674 11656 1730 11665
rect 1674 11591 1730 11600
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10010 1624 10406
rect 1688 10130 1716 11591
rect 1780 11150 1808 11750
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1596 9982 1716 10010
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1596 9042 1624 9687
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1308 8424 1360 8430
rect 1308 8366 1360 8372
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1320 7342 1348 7647
rect 1688 7546 1716 9982
rect 1780 9654 1808 11086
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1872 9042 1900 13194
rect 1964 11762 1992 13262
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 1964 10470 1992 11562
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1308 7336 1360 7342
rect 1308 7278 1360 7284
rect 1308 6860 1360 6866
rect 1308 6802 1360 6808
rect 1320 6497 1348 6802
rect 1780 6798 1808 8871
rect 1964 8090 1992 9454
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1306 6488 1362 6497
rect 1306 6423 1362 6432
rect 1780 6390 1808 6734
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1320 6089 1348 6190
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1320 5914 1348 6015
rect 1308 5908 1360 5914
rect 1308 5850 1360 5856
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 1360 5672 1362 5681
rect 1306 5607 1362 5616
rect 1306 5264 1362 5273
rect 1306 5199 1308 5208
rect 1360 5199 1362 5208
rect 1308 5170 1360 5176
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 1320 4690 1348 4791
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1766 4448 1822 4457
rect 1766 4383 1822 4392
rect 1780 4146 1808 4383
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1228 3641 1256 4082
rect 1308 4072 1360 4078
rect 1306 4040 1308 4049
rect 1360 4040 1362 4049
rect 1306 3975 1362 3984
rect 1780 3942 1808 4082
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1596 3738 1624 3878
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1214 3632 1270 3641
rect 2056 3602 2084 12650
rect 2148 6662 2176 17478
rect 2240 9586 2268 21490
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2332 9518 2360 13942
rect 2424 11762 2452 24142
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2504 21956 2556 21962
rect 2504 21898 2556 21904
rect 2516 18714 2544 21898
rect 2608 18986 2636 22374
rect 2792 22250 2820 22986
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2780 21480 2832 21486
rect 2884 21457 2912 22510
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 3252 21593 3280 22034
rect 3238 21584 3294 21593
rect 3238 21519 3294 21528
rect 3344 21486 3372 26302
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 3528 24274 3556 26200
rect 3606 25664 3662 25673
rect 3606 25599 3662 25608
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3436 23866 3464 24142
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 3436 22642 3464 23190
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 3332 21480 3384 21486
rect 2780 21422 2832 21428
rect 2870 21448 2926 21457
rect 2792 19961 2820 21422
rect 3332 21422 3384 21428
rect 2870 21383 2926 21392
rect 3424 21412 3476 21418
rect 3424 21354 3476 21360
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2778 19952 2834 19961
rect 2884 19938 2912 20810
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2884 19910 3004 19938
rect 2778 19887 2834 19896
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2778 19680 2834 19689
rect 2778 19615 2834 19624
rect 2792 19496 2820 19615
rect 2700 19468 2820 19496
rect 2700 19145 2728 19468
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2686 19136 2742 19145
rect 2686 19071 2742 19080
rect 2608 18958 2728 18986
rect 2516 18686 2636 18714
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2516 17066 2544 18566
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2516 12850 2544 17002
rect 2608 16726 2636 18686
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2700 14346 2728 18958
rect 2792 18329 2820 19314
rect 2884 18737 2912 19722
rect 2976 19553 3004 19910
rect 3344 19689 3372 20334
rect 3330 19680 3386 19689
rect 3330 19615 3386 19624
rect 2962 19544 3018 19553
rect 3436 19530 3464 21354
rect 2962 19479 3018 19488
rect 3344 19502 3464 19530
rect 3344 19145 3372 19502
rect 3330 19136 3386 19145
rect 2950 19068 3258 19077
rect 3330 19071 3386 19080
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2870 18728 2926 18737
rect 2870 18663 2926 18672
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 3344 18193 3372 19071
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 2778 18184 2834 18193
rect 2778 18119 2834 18128
rect 3330 18184 3386 18193
rect 3330 18119 3386 18128
rect 2792 16810 2820 18119
rect 3436 18086 3464 18566
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3422 17912 3478 17921
rect 3422 17847 3424 17856
rect 3476 17847 3478 17856
rect 3424 17818 3476 17824
rect 3528 17218 3556 23666
rect 3620 23202 3648 25599
rect 4066 25256 4122 25265
rect 4066 25191 4068 25200
rect 4120 25191 4122 25200
rect 4068 25162 4120 25168
rect 4066 24848 4122 24857
rect 4066 24783 4122 24792
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3712 23322 3740 24006
rect 3700 23316 3752 23322
rect 3700 23258 3752 23264
rect 3620 23174 3740 23202
rect 3804 23186 3832 24686
rect 4080 24682 4108 24783
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 3882 24032 3938 24041
rect 3882 23967 3938 23976
rect 3896 23526 3924 23967
rect 4068 23792 4120 23798
rect 4172 23780 4200 26200
rect 4802 24848 4858 24857
rect 4802 24783 4858 24792
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4120 23752 4200 23780
rect 4068 23734 4120 23740
rect 4068 23656 4120 23662
rect 4066 23624 4068 23633
rect 4120 23624 4122 23633
rect 4066 23559 4122 23568
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3988 23322 4200 23338
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 3976 23316 4200 23322
rect 4028 23310 4200 23316
rect 3976 23258 4028 23264
rect 3606 22808 3662 22817
rect 3606 22743 3662 22752
rect 3620 21729 3648 22743
rect 3712 22250 3740 23174
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3792 22636 3844 22642
rect 3792 22578 3844 22584
rect 3804 22409 3832 22578
rect 3790 22400 3846 22409
rect 3790 22335 3846 22344
rect 3896 22250 3924 23258
rect 4172 23066 4200 23310
rect 4264 23225 4292 24142
rect 4816 23730 4844 24783
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4250 23216 4306 23225
rect 4250 23151 4306 23160
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4172 23050 4292 23066
rect 4172 23044 4304 23050
rect 4172 23038 4252 23044
rect 4252 22986 4304 22992
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4172 22681 4200 22918
rect 4158 22672 4214 22681
rect 4158 22607 4214 22616
rect 4066 22536 4122 22545
rect 4122 22494 4200 22522
rect 4066 22471 4122 22480
rect 3712 22222 3832 22250
rect 3896 22222 4016 22250
rect 3700 22160 3752 22166
rect 3700 22102 3752 22108
rect 3606 21720 3662 21729
rect 3606 21655 3662 21664
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3344 17190 3556 17218
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2792 16782 2912 16810
rect 2778 16552 2834 16561
rect 2778 16487 2834 16496
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2608 12730 2636 13126
rect 2516 12702 2636 12730
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2516 10724 2544 12702
rect 2792 12170 2820 16487
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 11121 2636 11154
rect 2594 11112 2650 11121
rect 2792 11064 2820 12106
rect 2594 11047 2650 11056
rect 2700 11036 2820 11064
rect 2596 10736 2648 10742
rect 2516 10696 2596 10724
rect 2596 10678 2648 10684
rect 2608 10538 2636 10678
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2700 10062 2728 11036
rect 2778 10568 2834 10577
rect 2778 10503 2834 10512
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2240 8090 2268 8230
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2240 7274 2268 7890
rect 2228 7268 2280 7274
rect 2228 7210 2280 7216
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1214 3567 1270 3576
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1320 3233 1348 3470
rect 1306 3224 1362 3233
rect 1306 3159 1362 3168
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1320 2825 1348 2926
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1228 2417 1256 2450
rect 1214 2408 1270 2417
rect 1214 2343 1270 2352
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 2009 1348 2314
rect 1306 2000 1362 2009
rect 1306 1935 1362 1944
rect 1412 800 1440 2994
rect 2424 2990 2452 9862
rect 2792 9466 2820 10503
rect 2884 10266 2912 16782
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 3344 13705 3372 17190
rect 3422 16688 3478 16697
rect 3422 16623 3424 16632
rect 3476 16623 3478 16632
rect 3424 16594 3476 16600
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3436 14074 3464 15438
rect 3528 15162 3556 16050
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3330 13696 3386 13705
rect 2950 13628 3258 13637
rect 3330 13631 3386 13640
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3436 13190 3464 13738
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2608 9438 2820 9466
rect 2608 8022 2636 9438
rect 2778 9344 2834 9353
rect 2778 9279 2834 9288
rect 2792 8242 2820 9279
rect 2884 8974 2912 10095
rect 3240 9648 3292 9654
rect 3238 9616 3240 9625
rect 3292 9616 3294 9625
rect 3238 9551 3294 9560
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 2870 8528 2926 8537
rect 3252 8514 3280 8842
rect 3344 8634 3372 12718
rect 3528 12646 3556 14214
rect 3620 12986 3648 19314
rect 3712 18222 3740 22102
rect 3804 22094 3832 22222
rect 3804 22066 3924 22094
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3712 16833 3740 18022
rect 3804 17320 3832 20810
rect 3896 20534 3924 22066
rect 3988 21622 4016 22222
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3988 20777 4016 20878
rect 3974 20768 4030 20777
rect 3974 20703 4030 20712
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3804 17292 3924 17320
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3698 16824 3754 16833
rect 3698 16759 3754 16768
rect 3712 15026 3740 16759
rect 3804 16289 3832 17138
rect 3790 16280 3846 16289
rect 3896 16250 3924 17292
rect 3790 16215 3846 16224
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3528 12374 3556 12582
rect 3516 12368 3568 12374
rect 3436 12328 3516 12356
rect 3436 11354 3464 12328
rect 3516 12310 3568 12316
rect 3514 12200 3570 12209
rect 3514 12135 3570 12144
rect 3528 11898 3556 12135
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3514 11656 3570 11665
rect 3514 11591 3570 11600
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 10282 3556 11591
rect 3436 10254 3556 10282
rect 3620 10266 3648 12786
rect 3712 11354 3740 14962
rect 3804 12102 3832 15574
rect 3884 13320 3936 13326
rect 3882 13288 3884 13297
rect 3936 13288 3938 13297
rect 3882 13223 3938 13232
rect 3882 13016 3938 13025
rect 3882 12951 3938 12960
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3790 11520 3846 11529
rect 3790 11455 3846 11464
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3698 11248 3754 11257
rect 3698 11183 3754 11192
rect 3608 10260 3660 10266
rect 3436 10198 3464 10254
rect 3608 10202 3660 10208
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3424 10056 3476 10062
rect 3422 10024 3424 10033
rect 3476 10024 3478 10033
rect 3422 9959 3478 9968
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 8634 3464 8910
rect 3528 8634 3556 10066
rect 3606 9480 3662 9489
rect 3606 9415 3608 9424
rect 3660 9415 3662 9424
rect 3608 9386 3660 9392
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3252 8486 3464 8514
rect 3712 8498 3740 11183
rect 3804 11121 3832 11455
rect 3790 11112 3846 11121
rect 3790 11047 3846 11056
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 9926 3832 10406
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3804 9489 3832 9522
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3804 9178 3832 9415
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 2870 8463 2926 8472
rect 2700 8214 2820 8242
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2608 7886 2636 7958
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2700 7342 2728 8214
rect 2778 8120 2834 8129
rect 2778 8055 2834 8064
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2792 7154 2820 8055
rect 2884 7886 2912 8463
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 3344 8072 3372 8366
rect 3252 8044 3372 8072
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 3252 7750 3280 8044
rect 3330 7848 3386 7857
rect 3330 7783 3332 7792
rect 3384 7783 3386 7792
rect 3332 7754 3384 7760
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 2870 7304 2926 7313
rect 2870 7239 2926 7248
rect 2700 7126 2820 7154
rect 2596 6792 2648 6798
rect 2700 6746 2728 7126
rect 2780 6792 2832 6798
rect 2648 6740 2780 6746
rect 2596 6734 2832 6740
rect 2608 6718 2820 6734
rect 2884 6322 2912 7239
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3344 6905 3372 7346
rect 3436 7002 3464 8486
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3712 7750 3740 8434
rect 3896 8090 3924 12951
rect 3988 8634 4016 20402
rect 4172 19446 4200 22494
rect 4620 22500 4672 22506
rect 4620 22442 4672 22448
rect 4252 22092 4304 22098
rect 4252 22034 4304 22040
rect 4264 22001 4292 22034
rect 4250 21992 4306 22001
rect 4250 21927 4306 21936
rect 4250 21040 4306 21049
rect 4250 20975 4252 20984
rect 4304 20975 4306 20984
rect 4252 20946 4304 20952
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4264 18290 4292 19246
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4068 15496 4120 15502
rect 4066 15464 4068 15473
rect 4120 15464 4122 15473
rect 4066 15399 4122 15408
rect 4172 15026 4200 17614
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4264 17513 4292 17546
rect 4250 17504 4306 17513
rect 4250 17439 4306 17448
rect 4356 16182 4384 20470
rect 4434 19952 4490 19961
rect 4434 19887 4490 19896
rect 4448 19854 4476 19887
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4528 19780 4580 19786
rect 4528 19722 4580 19728
rect 4540 19666 4568 19722
rect 4448 19638 4568 19666
rect 4448 17134 4476 19638
rect 4632 19174 4660 22442
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4526 18864 4582 18873
rect 4526 18799 4582 18808
rect 4540 18766 4568 18799
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 17678 4660 18702
rect 4724 18630 4752 23122
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4816 22166 4844 22578
rect 4804 22160 4856 22166
rect 4804 22102 4856 22108
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4816 18630 4844 19722
rect 4712 18624 4764 18630
rect 4710 18592 4712 18601
rect 4804 18624 4856 18630
rect 4764 18592 4766 18601
rect 4804 18566 4856 18572
rect 4710 18527 4766 18536
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4724 17048 4752 18090
rect 4802 17640 4858 17649
rect 4802 17575 4858 17584
rect 4816 17542 4844 17575
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4632 17020 4752 17048
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4448 15570 4476 15914
rect 4436 15564 4488 15570
rect 4264 15524 4436 15552
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4264 14498 4292 15524
rect 4436 15506 4488 15512
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4172 14470 4292 14498
rect 4172 13818 4200 14470
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4264 13938 4292 14350
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4080 13790 4200 13818
rect 4080 12850 4108 13790
rect 4264 13682 4292 13874
rect 4172 13654 4292 13682
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4080 10146 4108 12679
rect 4172 12617 4200 13654
rect 4356 12918 4384 15302
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4448 13530 4476 14418
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 14113 4568 14214
rect 4526 14104 4582 14113
rect 4526 14039 4582 14048
rect 4526 13696 4582 13705
rect 4526 13631 4582 13640
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4158 12608 4214 12617
rect 4158 12543 4214 12552
rect 4158 12336 4214 12345
rect 4264 12306 4292 12718
rect 4356 12442 4384 12854
rect 4434 12608 4490 12617
rect 4434 12543 4490 12552
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4158 12271 4214 12280
rect 4252 12300 4304 12306
rect 4172 12238 4200 12271
rect 4252 12242 4304 12248
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4172 11830 4200 12174
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4080 10118 4200 10146
rect 4264 10130 4292 12242
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 10441 4384 12038
rect 4448 10810 4476 12543
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4342 10432 4398 10441
rect 4342 10367 4398 10376
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 4080 9110 4108 9959
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4172 8922 4200 10118
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4080 8894 4200 8922
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3804 7478 3832 8026
rect 3896 7857 3924 8026
rect 3882 7848 3938 7857
rect 3882 7783 3938 7792
rect 4080 7546 4108 8894
rect 4264 8498 4292 8910
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4264 8090 4292 8434
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3330 6896 3386 6905
rect 3330 6831 3332 6840
rect 3384 6831 3386 6840
rect 3332 6802 3384 6808
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3988 6390 4016 6598
rect 4356 6458 4384 10367
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4448 8294 4476 10202
rect 4540 10130 4568 13631
rect 4632 12918 4660 17020
rect 4710 16960 4766 16969
rect 4710 16895 4766 16904
rect 4724 15094 4752 16895
rect 4908 16590 4936 24346
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 5000 22094 5028 23462
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26330 7434 27000
rect 8022 26330 8078 27000
rect 6932 26302 7434 26330
rect 5460 23662 5488 26200
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5000 22066 5120 22094
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4816 14958 4844 15098
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4724 14074 4752 14214
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4816 13870 4844 14894
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4908 13716 4936 16186
rect 4724 13688 4936 13716
rect 4724 13258 4752 13688
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4804 13184 4856 13190
rect 5000 13138 5028 19178
rect 5092 17270 5120 22066
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 5078 17096 5134 17105
rect 5078 17031 5134 17040
rect 5092 16794 5120 17031
rect 5184 16998 5212 22986
rect 5368 22778 5396 23054
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5276 21486 5304 22374
rect 6012 22137 6040 23802
rect 6104 23186 6132 26200
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6564 24410 6592 24754
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6564 23526 6592 23666
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6472 22234 6500 22374
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 5998 22128 6054 22137
rect 6564 22094 6592 23462
rect 6656 23254 6684 23802
rect 6748 23474 6776 26200
rect 6932 24290 6960 26302
rect 7378 26200 7434 26302
rect 7852 26302 8078 26330
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 7288 24676 7340 24682
rect 7288 24618 7340 24624
rect 6840 24274 6960 24290
rect 6828 24268 6960 24274
rect 6880 24262 6960 24268
rect 6828 24210 6880 24216
rect 6748 23446 7052 23474
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 5998 22063 6054 22072
rect 6472 22066 6592 22094
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5828 21690 5856 21830
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5356 21480 5408 21486
rect 5644 21457 5672 21490
rect 5356 21422 5408 21428
rect 5630 21448 5686 21457
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5276 18057 5304 19450
rect 5368 19242 5396 21422
rect 5630 21383 5686 21392
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5460 20058 5488 20878
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5460 18170 5488 19178
rect 5368 18142 5488 18170
rect 5262 18048 5318 18057
rect 5262 17983 5318 17992
rect 5368 17082 5396 18142
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5276 17054 5396 17082
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5276 15994 5304 17054
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 4804 13126 4856 13132
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4632 8090 4660 9930
rect 4724 8906 4752 12854
rect 4816 12782 4844 13126
rect 4908 13110 5028 13138
rect 5092 15966 5304 15994
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 12238 4844 12718
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4908 11626 4936 13110
rect 5092 12170 5120 15966
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 14521 5212 15302
rect 5170 14512 5226 14521
rect 5170 14447 5226 14456
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5184 13394 5212 14350
rect 5276 13938 5304 15846
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5184 12306 5212 13330
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5276 11762 5304 13670
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 10130 4844 11086
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4908 9110 4936 11562
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 5000 7342 5028 11494
rect 5368 11064 5396 16934
rect 5460 16182 5488 18022
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5460 15094 5488 15642
rect 5552 15570 5580 21286
rect 5630 20904 5686 20913
rect 5630 20839 5632 20848
rect 5684 20839 5686 20848
rect 5632 20810 5684 20816
rect 5630 20088 5686 20097
rect 5630 20023 5686 20032
rect 5644 18290 5672 20023
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 18057 5672 18226
rect 5630 18048 5686 18057
rect 5630 17983 5686 17992
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5644 16250 5672 17002
rect 5736 16794 5764 21626
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 5828 20806 5856 21422
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5828 17134 5856 20334
rect 5908 20324 5960 20330
rect 5908 20266 5960 20272
rect 5920 18426 5948 20266
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5446 14648 5502 14657
rect 5446 14583 5502 14592
rect 5460 14550 5488 14583
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5460 12918 5488 13398
rect 5644 13002 5672 16050
rect 5736 15094 5764 16458
rect 5828 15910 5856 17070
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5736 14346 5764 14894
rect 5828 14822 5856 15506
rect 5920 15162 5948 18158
rect 6012 16250 6040 22063
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6104 20466 6132 21830
rect 6184 21616 6236 21622
rect 6184 21558 6236 21564
rect 6276 21616 6328 21622
rect 6276 21558 6328 21564
rect 6196 21350 6224 21558
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 20874 6224 21286
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6196 19802 6224 20810
rect 6288 19990 6316 21558
rect 6368 20800 6420 20806
rect 6472 20777 6500 22066
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6368 20742 6420 20748
rect 6458 20768 6514 20777
rect 6276 19984 6328 19990
rect 6276 19926 6328 19932
rect 6196 19786 6316 19802
rect 6196 19780 6328 19786
rect 6196 19774 6276 19780
rect 6276 19722 6328 19728
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6104 18737 6132 19110
rect 6090 18728 6146 18737
rect 6288 18698 6316 19722
rect 6090 18663 6146 18672
rect 6276 18692 6328 18698
rect 6104 18222 6132 18663
rect 6276 18634 6328 18640
rect 6182 18592 6238 18601
rect 6182 18527 6238 18536
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6090 18048 6146 18057
rect 6090 17983 6146 17992
rect 6104 17202 6132 17983
rect 6196 17814 6224 18527
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6288 17678 6316 18634
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14482 5856 14758
rect 5920 14618 5948 14962
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 5722 14104 5778 14113
rect 5722 14039 5778 14048
rect 5736 14006 5764 14039
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5552 12986 5672 13002
rect 5736 12986 5764 13806
rect 5828 13258 5856 14418
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5920 13190 5948 13738
rect 6012 13462 6040 16186
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 6104 15366 6132 15982
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 6104 14958 6132 15302
rect 6196 15162 6224 16662
rect 6288 15706 6316 17614
rect 6380 16046 6408 20742
rect 6458 20703 6514 20712
rect 6564 20097 6592 21966
rect 6550 20088 6606 20097
rect 6550 20023 6606 20032
rect 6552 19304 6604 19310
rect 6550 19272 6552 19281
rect 6604 19272 6606 19281
rect 6550 19207 6606 19216
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18290 6500 19110
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6472 17218 6500 18226
rect 6472 17190 6592 17218
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6472 16561 6500 16934
rect 6458 16552 6514 16561
rect 6458 16487 6514 16496
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6104 14822 6132 14894
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6104 13870 6132 14554
rect 6288 14346 6316 15642
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5540 12980 5672 12986
rect 5592 12974 5672 12980
rect 5724 12980 5776 12986
rect 5540 12922 5592 12928
rect 5724 12922 5776 12928
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5644 11898 5672 12582
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5632 11688 5684 11694
rect 5736 11642 5764 12106
rect 5684 11636 5764 11642
rect 5632 11630 5764 11636
rect 5540 11620 5592 11626
rect 5644 11614 5764 11630
rect 5540 11562 5592 11568
rect 5552 11218 5580 11562
rect 5736 11354 5764 11614
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5644 11218 5672 11290
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5276 11036 5396 11064
rect 5446 11112 5502 11121
rect 5446 11047 5502 11056
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 8634 5120 10610
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 9586 5212 10406
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5276 9178 5304 11036
rect 5354 10976 5410 10985
rect 5354 10911 5410 10920
rect 5368 10674 5396 10911
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5460 9586 5488 11047
rect 5630 10840 5686 10849
rect 5630 10775 5686 10784
rect 5644 10674 5672 10775
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5828 10062 5856 12854
rect 5920 11694 5948 13126
rect 6012 12782 6040 13194
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6104 12434 6132 13806
rect 6288 13326 6316 14282
rect 6380 14074 6408 15302
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6472 13954 6500 14894
rect 6564 14362 6592 17190
rect 6656 17066 6684 22578
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 6748 19514 6776 22374
rect 6840 22098 6868 22374
rect 7024 22098 7052 23446
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7208 22681 7236 23054
rect 7194 22672 7250 22681
rect 7194 22607 7250 22616
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6828 21412 6880 21418
rect 6828 21354 6880 21360
rect 6840 20602 6868 21354
rect 6932 21146 6960 21830
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 7024 21185 7052 21490
rect 7010 21176 7066 21185
rect 6920 21140 6972 21146
rect 7010 21111 7066 21120
rect 6920 21082 6972 21088
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 7024 20913 7052 21014
rect 7010 20904 7066 20913
rect 7010 20839 7066 20848
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6748 18426 6776 18634
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6840 16658 6868 20334
rect 6932 19242 6960 20470
rect 7024 19281 7052 20742
rect 7010 19272 7066 19281
rect 6920 19236 6972 19242
rect 7010 19207 7066 19216
rect 6920 19178 6972 19184
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6656 15502 6684 16118
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6656 14793 6684 14962
rect 6642 14784 6698 14793
rect 6642 14719 6698 14728
rect 6748 14482 6776 16390
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6564 14334 6776 14362
rect 6380 13926 6500 13954
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6288 12918 6316 13262
rect 6380 13190 6408 13926
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6012 12406 6132 12434
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5906 11112 5962 11121
rect 5906 11047 5962 11056
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5630 9888 5686 9897
rect 5630 9823 5686 9832
rect 5538 9616 5594 9625
rect 5448 9580 5500 9586
rect 5538 9551 5594 9560
rect 5448 9522 5500 9528
rect 5460 9178 5488 9522
rect 5552 9178 5580 9551
rect 5644 9382 5672 9823
rect 5920 9654 5948 11047
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5644 7750 5672 9318
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 6012 5778 6040 12406
rect 6288 12170 6316 12854
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6182 11248 6238 11257
rect 6182 11183 6238 11192
rect 6196 9042 6224 11183
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6380 7206 6408 13126
rect 6472 11898 6500 13738
rect 6550 13696 6606 13705
rect 6550 13631 6606 13640
rect 6564 13190 6592 13631
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6472 11801 6500 11834
rect 6458 11792 6514 11801
rect 6458 11727 6514 11736
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 10198 6500 11086
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6472 9722 6500 10134
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6458 8664 6514 8673
rect 6458 8599 6460 8608
rect 6512 8599 6514 8608
rect 6460 8570 6512 8576
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4146 2820 4422
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2884 1601 2912 3470
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2650 3372 2994
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3436 2514 3464 3334
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3804 2650 3832 2858
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 4080 800 4108 2450
rect 6564 2310 6592 13126
rect 6656 12986 6684 13806
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6748 12434 6776 14334
rect 6840 12850 6868 16594
rect 6932 16454 6960 19178
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 7116 16266 7144 22442
rect 7300 22094 7328 24618
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7208 22066 7328 22094
rect 7208 18222 7236 22066
rect 7286 21720 7342 21729
rect 7286 21655 7342 21664
rect 7300 20398 7328 21655
rect 7392 21622 7420 23598
rect 7484 23497 7512 23598
rect 7470 23488 7526 23497
rect 7470 23423 7526 23432
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7484 19938 7512 22918
rect 7576 22778 7604 22986
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7576 21457 7604 21966
rect 7562 21448 7618 21457
rect 7562 21383 7618 21392
rect 7668 20942 7696 22510
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7392 19910 7512 19938
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7194 17912 7250 17921
rect 7194 17847 7250 17856
rect 7208 17678 7236 17847
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 6932 16238 7144 16266
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6656 12406 6776 12434
rect 6656 10266 6684 12406
rect 6734 12336 6790 12345
rect 6734 12271 6790 12280
rect 6748 10742 6776 12271
rect 6840 11830 6868 12582
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6932 10606 6960 16238
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7024 11370 7052 16050
rect 7116 15473 7144 16118
rect 7208 15706 7236 17138
rect 7300 16522 7328 18362
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7392 16250 7420 19910
rect 7576 19514 7604 20742
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7470 19408 7526 19417
rect 7470 19343 7472 19352
rect 7524 19343 7526 19352
rect 7472 19314 7524 19320
rect 7576 18442 7604 19450
rect 7484 18414 7604 18442
rect 7484 17785 7512 18414
rect 7562 18320 7618 18329
rect 7562 18255 7618 18264
rect 7470 17776 7526 17785
rect 7470 17711 7526 17720
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7484 17513 7512 17546
rect 7470 17504 7526 17513
rect 7470 17439 7526 17448
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7286 16144 7342 16153
rect 7286 16079 7342 16088
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7300 15552 7328 16079
rect 7208 15524 7328 15552
rect 7102 15464 7158 15473
rect 7102 15399 7158 15408
rect 7116 13530 7144 15399
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7208 12442 7236 15524
rect 7380 15496 7432 15502
rect 7378 15464 7380 15473
rect 7432 15464 7434 15473
rect 7300 15422 7378 15450
rect 7300 14906 7328 15422
rect 7378 15399 7434 15408
rect 7484 15366 7512 17439
rect 7576 16153 7604 18255
rect 7668 17678 7696 20198
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7760 17338 7788 23666
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8312 24138 8340 26318
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26330 10654 27000
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8312 23769 8340 24074
rect 8298 23760 8354 23769
rect 7932 23724 7984 23730
rect 8298 23695 8354 23704
rect 7932 23666 7984 23672
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7944 23089 7972 23666
rect 7930 23080 7986 23089
rect 7930 23015 7986 23024
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 7852 17814 7880 22578
rect 8220 21894 8248 22578
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8206 20904 8262 20913
rect 8206 20839 8208 20848
rect 8260 20839 8262 20848
rect 8208 20810 8260 20816
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 19394 8340 19654
rect 8220 19366 8340 19394
rect 8220 18766 8248 19366
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8404 18442 8432 24142
rect 8576 23792 8628 23798
rect 8576 23734 8628 23740
rect 8484 23044 8536 23050
rect 8484 22986 8536 22992
rect 8496 21010 8524 22986
rect 8588 21010 8616 23734
rect 8680 22574 8708 26200
rect 9128 25220 9180 25226
rect 9128 25162 9180 25168
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8760 22024 8812 22030
rect 8758 21992 8760 22001
rect 8812 21992 8814 22001
rect 8758 21927 8814 21936
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8680 21622 8708 21830
rect 8668 21616 8720 21622
rect 8668 21558 8720 21564
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 19174 8524 20198
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8588 18902 8616 20810
rect 8680 20466 8708 21558
rect 8864 21536 8892 23054
rect 9048 22982 9076 23122
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9048 21894 9076 22918
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8944 21548 8996 21554
rect 8864 21508 8944 21536
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8680 19786 8708 20402
rect 8864 20398 8892 21508
rect 8944 21490 8996 21496
rect 8942 21448 8998 21457
rect 8942 21383 8998 21392
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8864 20058 8892 20334
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8956 19802 8984 21383
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 9048 19922 9076 20198
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 8668 19780 8720 19786
rect 8956 19774 9076 19802
rect 8668 19722 8720 19728
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8576 18896 8628 18902
rect 8576 18838 8628 18844
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8312 18414 8432 18442
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7944 17746 7972 18294
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7944 17626 7972 17682
rect 7852 17598 7972 17626
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7852 17134 7880 17598
rect 8036 17542 8064 17750
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8114 17232 8170 17241
rect 8114 17167 8170 17176
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 8128 16538 8156 17167
rect 8208 17128 8260 17134
rect 8206 17096 8208 17105
rect 8260 17096 8262 17105
rect 8206 17031 8262 17040
rect 8206 16688 8262 16697
rect 8206 16623 8208 16632
rect 8260 16623 8262 16632
rect 8208 16594 8260 16600
rect 8206 16552 8262 16561
rect 7748 16516 7800 16522
rect 8128 16510 8206 16538
rect 8206 16487 8262 16496
rect 7748 16458 7800 16464
rect 7562 16144 7618 16153
rect 7562 16079 7618 16088
rect 7564 16040 7616 16046
rect 7562 16008 7564 16017
rect 7616 16008 7618 16017
rect 7562 15943 7618 15952
rect 7654 15736 7710 15745
rect 7654 15671 7710 15680
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7392 15178 7420 15302
rect 7668 15178 7696 15671
rect 7392 15150 7696 15178
rect 7300 14878 7420 14906
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14074 7328 14758
rect 7392 14278 7420 14878
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7484 13870 7512 14486
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7484 13512 7512 13806
rect 7300 13484 7512 13512
rect 7300 13258 7328 13484
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7300 12374 7328 13194
rect 7392 12646 7420 13330
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7484 12889 7512 13194
rect 7470 12880 7526 12889
rect 7470 12815 7526 12824
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7392 11762 7420 12582
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7286 11384 7342 11393
rect 7024 11342 7236 11370
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7010 10704 7066 10713
rect 7010 10639 7066 10648
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 10470 6960 10542
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6642 8936 6698 8945
rect 6642 8871 6698 8880
rect 6656 8634 6684 8871
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6748 8022 6776 10406
rect 6918 10160 6974 10169
rect 6918 10095 6974 10104
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9110 6868 9454
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6932 8362 6960 10095
rect 7024 8430 7052 10639
rect 7116 9994 7144 11222
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7208 9330 7236 11342
rect 7484 11354 7512 12815
rect 7576 12306 7604 14826
rect 7668 14550 7696 15150
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7654 14376 7710 14385
rect 7760 14346 7788 16458
rect 8220 16454 8248 16487
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8208 16040 8260 16046
rect 8114 16008 8170 16017
rect 8208 15982 8260 15988
rect 8114 15943 8170 15952
rect 8128 15502 8156 15943
rect 8220 15706 8248 15982
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7840 14952 7892 14958
rect 7838 14920 7840 14929
rect 7892 14920 7894 14929
rect 7838 14855 7894 14864
rect 7852 14822 7880 14855
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7944 14550 7972 14962
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7654 14311 7710 14320
rect 7748 14340 7800 14346
rect 7668 14226 7696 14311
rect 7748 14282 7800 14288
rect 7840 14272 7892 14278
rect 7668 14198 7788 14226
rect 7840 14214 7892 14220
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7668 13190 7696 13738
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7576 11642 7604 12038
rect 7668 11830 7696 13126
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7576 11614 7696 11642
rect 7286 11319 7342 11328
rect 7472 11348 7524 11354
rect 7300 11218 7328 11319
rect 7472 11290 7524 11296
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7116 9302 7236 9330
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 4146 6868 7754
rect 7116 6730 7144 9302
rect 7194 9208 7250 9217
rect 7194 9143 7196 9152
rect 7248 9143 7250 9152
rect 7196 9114 7248 9120
rect 7300 7954 7328 11154
rect 7484 11150 7512 11290
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7668 10554 7696 11614
rect 7392 10538 7696 10554
rect 7380 10532 7696 10538
rect 7432 10526 7696 10532
rect 7380 10474 7432 10480
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7392 9382 7420 9930
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7484 8294 7512 10406
rect 7668 9722 7696 10526
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7760 9194 7788 14198
rect 7852 11642 7880 14214
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8312 12186 8340 18414
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8404 17882 8432 18226
rect 8496 18204 8524 18770
rect 8574 18728 8630 18737
rect 8574 18663 8630 18672
rect 8588 18630 8616 18663
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8576 18216 8628 18222
rect 8496 18176 8576 18204
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8404 17678 8432 17818
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8404 12764 8432 17206
rect 8496 16114 8524 18176
rect 8576 18158 8628 18164
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 17202 8616 17614
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8588 15638 8616 17002
rect 8680 15706 8708 19314
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8772 17134 8800 18634
rect 8864 17814 8892 19654
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 8956 18426 8984 18634
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8852 17808 8904 17814
rect 8852 17750 8904 17756
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8864 16640 8892 17750
rect 9048 17320 9076 19774
rect 9140 19446 9168 25162
rect 9324 24290 9352 26200
rect 9232 24274 9352 24290
rect 9220 24268 9352 24274
rect 9272 24262 9352 24268
rect 9220 24210 9272 24216
rect 9218 24168 9274 24177
rect 9218 24103 9274 24112
rect 9232 24070 9260 24103
rect 9220 24064 9272 24070
rect 9220 24006 9272 24012
rect 9232 20534 9260 24006
rect 9968 23798 9996 26200
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10048 25560 10100 25566
rect 10048 25502 10100 25508
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9402 22128 9458 22137
rect 9402 22063 9458 22072
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 9128 19440 9180 19446
rect 9232 19417 9260 20470
rect 9324 19825 9352 21830
rect 9416 21486 9444 22063
rect 9600 21622 9628 22986
rect 10060 22642 10088 25502
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 9864 22568 9916 22574
rect 9864 22510 9916 22516
rect 9876 22098 9904 22510
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9680 21888 9732 21894
rect 9678 21856 9680 21865
rect 9732 21856 9734 21865
rect 9678 21791 9734 21800
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9692 21350 9720 21626
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9404 20800 9456 20806
rect 9402 20768 9404 20777
rect 9456 20768 9458 20777
rect 9402 20703 9458 20712
rect 9404 20528 9456 20534
rect 9456 20476 9536 20482
rect 9404 20470 9536 20476
rect 9416 20454 9536 20470
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9310 19816 9366 19825
rect 9310 19751 9366 19760
rect 9128 19382 9180 19388
rect 9218 19408 9274 19417
rect 9218 19343 9274 19352
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9140 18737 9168 18770
rect 9126 18728 9182 18737
rect 9126 18663 9182 18672
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9140 18358 9168 18566
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 9232 17610 9260 18566
rect 9416 17746 9444 20334
rect 9508 20058 9536 20454
rect 9496 20052 9548 20058
rect 9496 19994 9548 20000
rect 9508 19786 9536 19994
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18222 9536 19110
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9600 18086 9628 20810
rect 9692 18329 9720 21286
rect 9784 18884 9812 21966
rect 10060 20262 10088 21966
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10140 19304 10192 19310
rect 10138 19272 10140 19281
rect 10192 19272 10194 19281
rect 10138 19207 10194 19216
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 9864 18896 9916 18902
rect 9784 18856 9864 18884
rect 9864 18838 9916 18844
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9864 18760 9916 18766
rect 9784 18720 9864 18748
rect 9678 18320 9734 18329
rect 9678 18255 9734 18264
rect 9588 18080 9640 18086
rect 9494 18048 9550 18057
rect 9588 18022 9640 18028
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9494 17983 9550 17992
rect 9508 17864 9536 17983
rect 9508 17836 9628 17864
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9310 17368 9366 17377
rect 8772 16612 8892 16640
rect 8956 17292 9076 17320
rect 9128 17332 9180 17338
rect 8772 16182 8800 16612
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8496 15434 8524 15506
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8588 15026 8616 15302
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8772 14940 8800 15846
rect 8956 15042 8984 17292
rect 9180 17292 9260 17320
rect 9416 17354 9444 17546
rect 9366 17326 9444 17354
rect 9494 17368 9550 17377
rect 9310 17303 9366 17312
rect 9494 17303 9496 17312
rect 9128 17274 9180 17280
rect 9232 17218 9260 17292
rect 9548 17303 9550 17312
rect 9496 17274 9548 17280
rect 9232 17202 9536 17218
rect 9232 17196 9548 17202
rect 9232 17190 9496 17196
rect 9600 17184 9628 17836
rect 9692 17184 9720 18022
rect 9600 17156 9720 17184
rect 9496 17138 9548 17144
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9416 16998 9444 17070
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9218 16824 9274 16833
rect 9218 16759 9220 16768
rect 9272 16759 9274 16768
rect 9220 16730 9272 16736
rect 9416 16726 9444 16934
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9232 15638 9260 16458
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 8680 14912 8800 14940
rect 8864 15014 8984 15042
rect 8574 14512 8630 14521
rect 8574 14447 8630 14456
rect 8588 14006 8616 14447
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8588 12918 8616 13398
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8404 12736 8616 12764
rect 8312 12158 8524 12186
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 7852 11614 7972 11642
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 10470 7880 11494
rect 7944 11218 7972 11614
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8128 11150 8156 11766
rect 8116 11144 8168 11150
rect 8168 11104 8340 11132
rect 8116 11086 8168 11092
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8312 10742 8340 11104
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 10130 7880 10406
rect 8128 10198 8156 10542
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7852 9518 7880 10066
rect 8220 9908 8248 10406
rect 8312 10130 8340 10678
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8392 9920 8444 9926
rect 8220 9880 8340 9908
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8312 9636 8340 9880
rect 8392 9862 8444 9868
rect 8220 9608 8340 9636
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7668 9166 7788 9194
rect 7668 8838 7696 9166
rect 7746 9072 7802 9081
rect 7746 9007 7802 9016
rect 7760 8974 7788 9007
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7576 8090 7604 8434
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7576 2650 7604 5782
rect 7852 3058 7880 9454
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 9042 8156 9318
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8220 8838 8248 9608
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8128 8430 8156 8570
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8312 8090 8340 8774
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8404 7274 8432 9862
rect 8496 9654 8524 12158
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8496 8294 8524 9590
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8588 7886 8616 12736
rect 8680 8974 8708 14912
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 12918 8800 13670
rect 8760 12912 8812 12918
rect 8758 12880 8760 12889
rect 8812 12880 8814 12889
rect 8758 12815 8814 12824
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 11082 8800 11494
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8864 9674 8892 15014
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8956 14278 8984 14894
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 12374 8984 14214
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 9048 11626 9076 12718
rect 9140 12170 9168 15574
rect 9218 15464 9274 15473
rect 9218 15399 9220 15408
rect 9272 15399 9274 15408
rect 9220 15370 9272 15376
rect 9324 15162 9352 16662
rect 9508 16232 9536 16934
rect 9416 16204 9536 16232
rect 9416 15570 9444 16204
rect 9494 16144 9550 16153
rect 9600 16130 9628 16934
rect 9692 16561 9720 17156
rect 9784 17134 9812 18720
rect 9864 18702 9916 18708
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17202 9904 18022
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9678 16552 9734 16561
rect 9678 16487 9734 16496
rect 9550 16102 9628 16130
rect 9494 16079 9550 16088
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9588 15360 9640 15366
rect 9692 15314 9720 16487
rect 9876 15910 9904 17138
rect 9968 16046 9996 18770
rect 10244 18698 10272 19178
rect 10336 18834 10364 19314
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10060 17746 10088 18634
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10152 17134 10180 18362
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9640 15308 9720 15314
rect 9588 15302 9720 15308
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9600 15286 9720 15302
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9402 15056 9458 15065
rect 9312 15020 9364 15026
rect 9402 14991 9458 15000
rect 9312 14962 9364 14968
rect 9324 13954 9352 14962
rect 9416 14618 9444 14991
rect 9508 14793 9536 15098
rect 9678 15056 9734 15065
rect 9678 14991 9734 15000
rect 9692 14958 9720 14991
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 14816 9640 14822
rect 9494 14784 9550 14793
rect 9588 14758 9640 14764
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9494 14719 9550 14728
rect 9600 14618 9628 14758
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9232 13926 9352 13954
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9140 11762 9168 12106
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 9048 11286 9076 11562
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9140 10266 9168 11698
rect 9232 11150 9260 13926
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9324 12646 9352 13806
rect 9404 13320 9456 13326
rect 9402 13288 9404 13297
rect 9456 13288 9458 13297
rect 9402 13223 9458 13232
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12306 9352 12582
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9312 11824 9364 11830
rect 9310 11792 9312 11801
rect 9364 11792 9366 11801
rect 9310 11727 9366 11736
rect 9416 11200 9444 12310
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9324 11172 9444 11200
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8772 9646 8892 9674
rect 9048 9654 9076 10066
rect 9036 9648 9088 9654
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8772 8498 8800 9646
rect 9036 9590 9088 9596
rect 9048 8838 9076 9590
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8498 9076 8774
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 9140 7546 9168 8842
rect 9324 8378 9352 11172
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 9042 9444 11018
rect 9508 10674 9536 11766
rect 9600 11218 9628 14010
rect 9692 12238 9720 14758
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 14385 9812 14418
rect 9770 14376 9826 14385
rect 9770 14311 9826 14320
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 13841 9812 14214
rect 9770 13832 9826 13841
rect 9770 13767 9826 13776
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9324 8350 9444 8378
rect 9310 8256 9366 8265
rect 9310 8191 9366 8200
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9324 7410 9352 8191
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 9416 5166 9444 8350
rect 9600 7478 9628 10950
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 9178 9720 9522
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 9692 3738 9720 8774
rect 9784 6866 9812 12106
rect 9876 8480 9904 15302
rect 9968 12782 9996 15982
rect 10060 15706 10088 16118
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10152 14482 10180 15982
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 10046 13832 10102 13841
rect 10046 13767 10102 13776
rect 10060 13734 10088 13767
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13530 10180 13670
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10048 12640 10100 12646
rect 9954 12608 10010 12617
rect 10048 12582 10100 12588
rect 9954 12543 10010 12552
rect 9968 11830 9996 12543
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10060 8566 10088 12582
rect 10152 9178 10180 12718
rect 10244 11558 10272 18226
rect 10428 18086 10456 25162
rect 10612 24206 10640 25638
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10704 22710 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10796 22030 10824 25434
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 11072 24313 11100 24346
rect 11058 24304 11114 24313
rect 11058 24239 11114 24248
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11164 22545 11192 23666
rect 11150 22536 11206 22545
rect 11150 22471 11206 22480
rect 11256 22098 11284 26200
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11716 24410 11744 24550
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11336 23588 11388 23594
rect 11336 23530 11388 23536
rect 11348 22982 11376 23530
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 11440 23186 11468 23462
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11336 22976 11388 22982
rect 11336 22918 11388 22924
rect 11900 22778 11928 26200
rect 12072 25764 12124 25770
rect 12072 25706 12124 25712
rect 11980 24336 12032 24342
rect 11980 24278 12032 24284
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10520 21593 10548 21966
rect 11520 21888 11572 21894
rect 10966 21856 11022 21865
rect 11520 21830 11572 21836
rect 10966 21791 11022 21800
rect 10980 21690 11008 21791
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 10506 21584 10562 21593
rect 10506 21519 10562 21528
rect 11532 21350 11560 21830
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10704 19514 10732 20266
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10796 19854 10824 19994
rect 10888 19922 10916 20198
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10796 19174 10824 19314
rect 10980 19310 11008 20334
rect 11072 19786 11100 21286
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 11164 19718 11192 20198
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10520 18442 10548 18770
rect 10520 18414 10640 18442
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10612 17882 10640 18414
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 10336 12646 10364 17750
rect 10796 17513 10824 19110
rect 10874 17776 10930 17785
rect 10874 17711 10930 17720
rect 10888 17678 10916 17711
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10782 17504 10838 17513
rect 10782 17439 10838 17448
rect 10414 17368 10470 17377
rect 10414 17303 10470 17312
rect 10428 16794 10456 17303
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10428 16590 10456 16730
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10428 15570 10456 15642
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10520 15042 10548 16390
rect 10598 16280 10654 16289
rect 10598 16215 10654 16224
rect 10612 16114 10640 16215
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10612 15094 10640 16050
rect 10428 15014 10548 15042
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10428 14958 10456 15014
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10520 14385 10548 14826
rect 10704 14482 10732 17070
rect 10888 16046 10916 17614
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10980 16114 11008 16526
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10966 16008 11022 16017
rect 10784 15972 10836 15978
rect 10966 15943 10968 15952
rect 10784 15914 10836 15920
rect 11020 15943 11022 15952
rect 10968 15914 11020 15920
rect 10796 15570 10824 15914
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10966 15328 11022 15337
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10796 14550 10824 14826
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10506 14376 10562 14385
rect 10506 14311 10562 14320
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10428 11150 10456 13126
rect 10520 12714 10548 14214
rect 10612 12986 10640 14214
rect 10704 13025 10732 14418
rect 10796 14278 10824 14486
rect 10888 14414 10916 15302
rect 10966 15263 11022 15272
rect 10980 15094 11008 15263
rect 10968 15088 11020 15094
rect 10966 15056 10968 15065
rect 11020 15056 11022 15065
rect 10966 14991 11022 15000
rect 10968 14952 11020 14958
rect 10966 14920 10968 14929
rect 11020 14920 11022 14929
rect 10966 14855 11022 14864
rect 11072 14657 11100 19246
rect 11164 18834 11192 19654
rect 11256 19281 11284 20946
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11242 19272 11298 19281
rect 11242 19207 11298 19216
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 18630 11284 18702
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11348 16538 11376 20810
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11440 19961 11468 20742
rect 11426 19952 11482 19961
rect 11426 19887 11482 19896
rect 11428 19440 11480 19446
rect 11426 19408 11428 19417
rect 11480 19408 11482 19417
rect 11426 19343 11482 19352
rect 11532 17814 11560 21286
rect 11610 21176 11666 21185
rect 11610 21111 11666 21120
rect 11624 20806 11652 21111
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11624 19378 11652 20198
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11716 18850 11744 22510
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 21078 11836 21286
rect 11796 21072 11848 21078
rect 11796 21014 11848 21020
rect 11992 20890 12020 24278
rect 12084 21010 12112 25706
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12268 23866 12296 25298
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 12360 23866 12388 24618
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12268 23050 12296 23462
rect 12452 23304 12480 23802
rect 12544 23798 12572 26200
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12636 24206 12664 24686
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13280 23633 13308 23666
rect 13266 23624 13322 23633
rect 13266 23559 13322 23568
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12360 23276 12480 23304
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12360 22642 12388 23276
rect 12820 23254 12848 23462
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12452 22574 12480 23122
rect 12544 22982 12572 23122
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12176 21146 12204 21490
rect 12452 21486 12480 22510
rect 12544 21570 12572 22714
rect 12728 22710 12756 22918
rect 12820 22710 12848 23190
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12716 22704 12768 22710
rect 12716 22646 12768 22652
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 12636 22098 12664 22646
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12544 21542 12664 21570
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12268 21078 12296 21422
rect 12346 21176 12402 21185
rect 12346 21111 12348 21120
rect 12400 21111 12402 21120
rect 12348 21082 12400 21088
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12636 21010 12664 21542
rect 12728 21418 12756 22646
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13372 22098 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 13728 25628 13780 25634
rect 13728 25570 13780 25576
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13556 23497 13584 24754
rect 13740 24750 13768 25570
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13832 24138 13860 26200
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13634 23760 13690 23769
rect 13634 23695 13690 23704
rect 13542 23488 13598 23497
rect 13542 23423 13598 23432
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13360 21480 13412 21486
rect 13464 21468 13492 22374
rect 13556 22098 13584 22918
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13412 21440 13492 21468
rect 13360 21422 13412 21428
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 11992 20862 12112 20890
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11794 20496 11850 20505
rect 11794 20431 11850 20440
rect 11808 20058 11836 20431
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11900 19666 11928 20742
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11992 20369 12020 20402
rect 11978 20360 12034 20369
rect 11978 20295 12034 20304
rect 12084 20058 12112 20862
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 13372 19922 13400 21422
rect 13544 20800 13596 20806
rect 13648 20788 13676 23695
rect 13924 21962 13952 25230
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14292 24410 14320 24754
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14476 24342 14504 26200
rect 14648 25424 14700 25430
rect 14648 25366 14700 25372
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14476 23361 14504 24142
rect 14186 23352 14242 23361
rect 14186 23287 14242 23296
rect 14462 23352 14518 23361
rect 14462 23287 14518 23296
rect 14200 22234 14228 23287
rect 14370 23080 14426 23089
rect 14370 23015 14372 23024
rect 14424 23015 14426 23024
rect 14372 22986 14424 22992
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14660 22001 14688 25366
rect 14740 24880 14792 24886
rect 14740 24822 14792 24828
rect 14646 21992 14702 22001
rect 13912 21956 13964 21962
rect 14646 21927 14648 21936
rect 13912 21898 13964 21904
rect 14700 21927 14702 21936
rect 14648 21898 14700 21904
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14108 21486 14136 21830
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13596 20760 13676 20788
rect 13544 20742 13596 20748
rect 13740 20466 13768 21286
rect 13910 21176 13966 21185
rect 13910 21111 13966 21120
rect 13924 20806 13952 21111
rect 14384 21078 14412 21354
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 13912 20800 13964 20806
rect 13910 20768 13912 20777
rect 13964 20768 13966 20777
rect 13910 20703 13966 20712
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13556 20233 13584 20402
rect 13636 20256 13688 20262
rect 13542 20224 13598 20233
rect 13636 20198 13688 20204
rect 13542 20159 13598 20168
rect 13544 19984 13596 19990
rect 13544 19926 13596 19932
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12990 19816 13046 19825
rect 12990 19751 13046 19760
rect 13268 19780 13320 19786
rect 13004 19718 13032 19751
rect 13268 19722 13320 19728
rect 11808 19638 11928 19666
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 11808 18986 11836 19638
rect 11900 19514 12204 19530
rect 11888 19508 12204 19514
rect 11940 19502 12204 19508
rect 11888 19450 11940 19456
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 12176 19394 12204 19502
rect 13280 19446 13308 19722
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13268 19440 13320 19446
rect 11808 18958 11928 18986
rect 11716 18822 11836 18850
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 17270 11468 17682
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11164 16510 11376 16538
rect 11164 15201 11192 16510
rect 11440 16402 11468 17206
rect 11624 16998 11652 18566
rect 11716 18086 11744 18634
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 17649 11744 18022
rect 11702 17640 11758 17649
rect 11702 17575 11758 17584
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11348 16374 11468 16402
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11150 15192 11206 15201
rect 11150 15127 11206 15136
rect 11058 14648 11114 14657
rect 11058 14583 11114 14592
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 11072 14414 11100 14447
rect 10876 14408 10928 14414
rect 11060 14408 11112 14414
rect 10876 14350 10928 14356
rect 10966 14376 11022 14385
rect 11060 14350 11112 14356
rect 10966 14311 11022 14320
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10876 13932 10928 13938
rect 10796 13892 10876 13920
rect 10796 13841 10824 13892
rect 10876 13874 10928 13880
rect 10980 13870 11008 14311
rect 11072 14226 11100 14350
rect 11072 14198 11192 14226
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10968 13864 11020 13870
rect 10782 13832 10838 13841
rect 10968 13806 11020 13812
rect 10782 13767 10838 13776
rect 10690 13016 10746 13025
rect 10600 12980 10652 12986
rect 10690 12951 10746 12960
rect 10600 12922 10652 12928
rect 10690 12880 10746 12889
rect 10690 12815 10692 12824
rect 10744 12815 10746 12824
rect 10692 12786 10744 12792
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11830 10640 12038
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9876 8452 9996 8480
rect 9862 8392 9918 8401
rect 9862 8327 9864 8336
rect 9916 8327 9918 8336
rect 9864 8298 9916 8304
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9968 4690 9996 8452
rect 10244 8294 10272 10474
rect 10336 9518 10364 10610
rect 10612 9654 10640 11290
rect 10704 10606 10732 12786
rect 10796 12714 10824 13767
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10888 12442 10916 13126
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10796 10266 10824 10950
rect 10980 10674 11008 13806
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10888 9518 10916 10134
rect 10980 10062 11008 10202
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10336 7954 10364 9454
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6748 800 6776 2450
rect 8312 2446 8340 2790
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9416 800 9444 2450
rect 9784 2446 9812 3130
rect 10428 3126 10456 8434
rect 10520 6866 10548 8434
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10612 3942 10640 8366
rect 11072 7886 11100 14010
rect 11164 13530 11192 14198
rect 11256 13802 11284 15982
rect 11348 15881 11376 16374
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11334 15872 11390 15881
rect 11334 15807 11390 15816
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 11348 13938 11376 15370
rect 11440 15366 11468 15982
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11532 13870 11560 16730
rect 11624 16658 11652 16934
rect 11702 16824 11758 16833
rect 11702 16759 11758 16768
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11334 13696 11390 13705
rect 11334 13631 11390 13640
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12170 11192 12582
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11150 11656 11206 11665
rect 11150 11591 11206 11600
rect 11164 11558 11192 11591
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11256 11370 11284 13330
rect 11348 12374 11376 13631
rect 11532 13394 11560 13806
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11348 11762 11376 12310
rect 11336 11756 11388 11762
rect 11440 11744 11468 12582
rect 11624 12434 11652 16594
rect 11716 16046 11744 16759
rect 11808 16522 11836 18822
rect 11900 16794 11928 18958
rect 11992 17678 12020 19382
rect 12176 19366 12572 19394
rect 13268 19382 13320 19388
rect 12070 19272 12126 19281
rect 12070 19207 12126 19216
rect 12084 18222 12112 19207
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12162 18184 12218 18193
rect 12162 18119 12164 18128
rect 12216 18119 12218 18128
rect 12164 18090 12216 18096
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11992 16114 12020 17614
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 12084 17066 12112 17478
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 12268 16182 12296 17546
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 13326 11744 15846
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11808 12986 11836 16050
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12072 15632 12124 15638
rect 12070 15600 12072 15609
rect 12124 15600 12126 15609
rect 12070 15535 12126 15544
rect 12268 15416 12296 15982
rect 12084 15388 12296 15416
rect 11886 15192 11942 15201
rect 11886 15127 11942 15136
rect 11900 15026 11928 15127
rect 11978 15056 12034 15065
rect 11888 15020 11940 15026
rect 11978 14991 11980 15000
rect 11888 14962 11940 14968
rect 12032 14991 12034 15000
rect 11980 14962 12032 14968
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11624 12406 11744 12434
rect 11440 11716 11652 11744
rect 11336 11698 11388 11704
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11256 11342 11468 11370
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11164 8634 11192 10678
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10062 11284 10542
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9518 11284 9998
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11348 8974 11376 11222
rect 11440 11098 11468 11342
rect 11532 11218 11560 11562
rect 11624 11354 11652 11716
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11440 11070 11652 11098
rect 11520 10464 11572 10470
rect 11518 10432 11520 10441
rect 11572 10432 11574 10441
rect 11518 10367 11574 10376
rect 11428 9920 11480 9926
rect 11480 9897 11560 9908
rect 11480 9888 11574 9897
rect 11480 9880 11518 9888
rect 11428 9862 11480 9868
rect 11518 9823 11574 9832
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11256 8566 11284 8774
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11440 7478 11468 9318
rect 11532 8634 11560 9823
rect 11624 8838 11652 11070
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11716 7546 11744 12406
rect 11900 12186 11928 14962
rect 12084 14929 12112 15388
rect 12360 15348 12388 18226
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12176 15320 12388 15348
rect 12070 14920 12126 14929
rect 12070 14855 12126 14864
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13394 12020 14350
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13938 12112 14010
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11900 12158 12020 12186
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11808 10470 11836 11562
rect 11796 10464 11848 10470
rect 11900 10441 11928 12038
rect 11992 10742 12020 12158
rect 12084 11558 12112 12242
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 10742 12112 11494
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11796 10406 11848 10412
rect 11886 10432 11942 10441
rect 11808 9994 11836 10406
rect 11886 10367 11942 10376
rect 12176 10266 12204 15320
rect 12452 15162 12480 18158
rect 12544 17338 12572 19366
rect 12714 19136 12770 19145
rect 12714 19071 12770 19080
rect 12728 18630 12756 19071
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12820 18358 12848 18634
rect 13372 18426 13400 19654
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 17746 12664 18158
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12544 16794 12572 17138
rect 12636 16794 12664 17682
rect 12728 17610 12756 18022
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13464 17882 13492 19314
rect 13556 18834 13584 19926
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13268 17808 13320 17814
rect 13266 17776 13268 17785
rect 13320 17776 13322 17785
rect 12808 17740 12860 17746
rect 13266 17711 13322 17720
rect 12808 17682 12860 17688
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12716 16992 12768 16998
rect 12820 16969 12848 17682
rect 12716 16934 12768 16940
rect 12806 16960 12862 16969
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12544 16250 12572 16594
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12636 15745 12664 15982
rect 12622 15736 12678 15745
rect 12622 15671 12678 15680
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12268 12646 12296 13806
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12360 12306 12388 13194
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12360 11354 12388 12242
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11888 9920 11940 9926
rect 11992 9908 12020 10066
rect 11940 9880 12020 9908
rect 11888 9862 11940 9868
rect 11992 9654 12020 9880
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 7546 11928 8842
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 12084 3738 12112 7754
rect 12268 6254 12296 11290
rect 12452 9382 12480 13466
rect 12544 12442 12572 15302
rect 12728 14464 12756 16934
rect 12806 16895 12862 16904
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13176 16448 13228 16454
rect 13174 16416 13176 16425
rect 13360 16448 13412 16454
rect 13228 16416 13230 16425
rect 13360 16390 13412 16396
rect 13174 16351 13230 16360
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15706 13400 16390
rect 13648 15722 13676 20198
rect 13740 19990 13768 20402
rect 13910 20360 13966 20369
rect 13910 20295 13966 20304
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13924 19718 13952 20295
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13924 19446 13952 19654
rect 14108 19514 14136 19926
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13740 17882 13768 19246
rect 13832 19174 13860 19382
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18086 13860 19110
rect 14108 18358 14136 19450
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 14200 17921 14228 21014
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14186 17912 14242 17921
rect 13728 17876 13780 17882
rect 14186 17847 14242 17856
rect 13728 17818 13780 17824
rect 13740 17134 13768 17818
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13832 17270 13860 17546
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13740 16250 13768 16730
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13924 15881 13952 17138
rect 14004 15904 14056 15910
rect 13910 15872 13966 15881
rect 14004 15846 14056 15852
rect 13910 15807 13966 15816
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13556 15694 13676 15722
rect 13726 15736 13782 15745
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12820 14482 12848 15506
rect 13556 15042 13584 15694
rect 13726 15671 13782 15680
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13464 15014 13584 15042
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14618 13400 14962
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 12636 14436 12756 14464
rect 12808 14476 12860 14482
rect 12636 13138 12664 14436
rect 12808 14418 12860 14424
rect 12820 13530 12848 14418
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13524 12860 13530
rect 13372 13512 13400 13670
rect 12808 13466 12860 13472
rect 13188 13484 13400 13512
rect 12636 13110 12756 13138
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12442 12664 12650
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12636 11626 12664 12174
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9654 12664 9998
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8498 12480 8774
rect 12728 8514 12756 13110
rect 13188 12918 13216 13484
rect 13268 13388 13320 13394
rect 13320 13348 13400 13376
rect 13268 13330 13320 13336
rect 13372 12918 13400 13348
rect 13464 12986 13492 15014
rect 13542 14920 13598 14929
rect 13542 14855 13598 14864
rect 13556 14618 13584 14855
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13176 12776 13228 12782
rect 13174 12744 13176 12753
rect 13228 12744 13230 12753
rect 13174 12679 13230 12688
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13176 12096 13228 12102
rect 13280 12073 13308 12310
rect 13176 12038 13228 12044
rect 13266 12064 13322 12073
rect 13188 11937 13216 12038
rect 13266 11999 13322 12008
rect 13174 11928 13230 11937
rect 13174 11863 13230 11872
rect 13372 11830 13400 12854
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13464 12646 13492 12786
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13176 11620 13228 11626
rect 13228 11580 13400 11608
rect 13176 11562 13228 11568
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13372 11354 13400 11580
rect 13464 11354 13492 12582
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13372 9450 13400 11154
rect 13556 10130 13584 13874
rect 13648 13190 13676 15574
rect 13740 15502 13768 15671
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13740 12986 13768 15302
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14618 13860 14962
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13924 14278 13952 15302
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13530 13860 13806
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13924 13258 13952 14214
rect 14016 14006 14044 15846
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13556 9042 13584 9318
rect 13648 9110 13676 12922
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 10810 13860 12718
rect 13924 12442 13952 13194
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12646 14044 13126
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13924 12102 13952 12378
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11354 13952 12038
rect 14108 11898 14136 17138
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14200 16697 14228 17070
rect 14186 16688 14242 16697
rect 14292 16658 14320 17206
rect 14186 16623 14242 16632
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14384 16454 14412 20742
rect 14568 20398 14596 21286
rect 14752 20584 14780 24822
rect 15014 22400 15070 22409
rect 15014 22335 15070 22344
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14936 21146 14964 21830
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 15028 21010 15056 22335
rect 15120 22166 15148 26200
rect 15660 25084 15712 25090
rect 15660 25026 15712 25032
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 15212 22030 15240 24890
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 14660 20556 14780 20584
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14568 19854 14596 19926
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14476 19446 14504 19790
rect 14660 19718 14688 20556
rect 15120 20482 15148 21082
rect 15212 20874 15240 21966
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 15304 21010 15332 21558
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 15304 20534 15332 20946
rect 15396 20618 15424 24142
rect 15566 21448 15622 21457
rect 15566 21383 15568 21392
rect 15620 21383 15622 21392
rect 15568 21354 15620 21360
rect 15396 20590 15608 20618
rect 14752 20454 15148 20482
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19514 14688 19654
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18873 14504 19110
rect 14462 18864 14518 18873
rect 14462 18799 14518 18808
rect 14568 16810 14596 19314
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14660 17338 14688 18294
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14568 16782 14688 16810
rect 14556 16720 14608 16726
rect 14554 16688 14556 16697
rect 14608 16688 14610 16697
rect 14464 16652 14516 16658
rect 14554 16623 14610 16632
rect 14464 16594 14516 16600
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14200 14074 14228 15030
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14414 14320 14894
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14200 12764 14228 13738
rect 14292 13326 14320 14350
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12918 14320 13262
rect 14384 13190 14412 15506
rect 14476 13870 14504 16594
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14200 12736 14412 12764
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14200 11694 14228 12582
rect 14384 12434 14412 12736
rect 14476 12442 14504 12922
rect 14292 12406 14412 12434
rect 14464 12436 14516 12442
rect 14292 11801 14320 12406
rect 14464 12378 14516 12384
rect 14370 11928 14426 11937
rect 14568 11914 14596 15642
rect 14660 13734 14688 16782
rect 14752 15706 14780 20454
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 14924 19304 14976 19310
rect 15028 19281 15056 20334
rect 14924 19246 14976 19252
rect 15014 19272 15070 19281
rect 14830 18456 14886 18465
rect 14830 18391 14886 18400
rect 14844 17490 14872 18391
rect 14936 17814 14964 19246
rect 15014 19207 15070 19216
rect 15212 18986 15240 20334
rect 15304 19786 15332 20470
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15304 19378 15332 19722
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15028 18970 15240 18986
rect 15016 18964 15240 18970
rect 15068 18958 15240 18964
rect 15016 18906 15068 18912
rect 15396 18630 15424 20402
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19922 15516 20198
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 15028 18329 15056 18362
rect 15014 18320 15070 18329
rect 15014 18255 15070 18264
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 14936 17490 14964 17546
rect 15028 17542 15056 17614
rect 15120 17542 15148 18158
rect 15382 18048 15438 18057
rect 15382 17983 15438 17992
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 14844 17462 14964 17490
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14844 15162 14872 17274
rect 14936 17202 14964 17462
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15028 17082 15056 17478
rect 14936 17054 15056 17082
rect 14936 16114 14964 17054
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14752 14618 14780 15030
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14936 14618 14964 14894
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14752 14056 14780 14554
rect 14832 14068 14884 14074
rect 14752 14028 14832 14056
rect 14832 14010 14884 14016
rect 14936 13870 14964 14554
rect 15028 14278 15056 16662
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 15120 12850 15148 17478
rect 15212 16810 15240 17478
rect 15304 17202 15332 17546
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15396 16946 15424 17983
rect 15488 17134 15516 18634
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15396 16918 15516 16946
rect 15212 16782 15424 16810
rect 15396 16590 15424 16782
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15304 14362 15332 16526
rect 15488 16130 15516 16918
rect 15580 16726 15608 20590
rect 15672 19378 15700 25026
rect 15764 23798 15792 26200
rect 15936 25016 15988 25022
rect 15936 24958 15988 24964
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15750 21720 15806 21729
rect 15750 21655 15806 21664
rect 15764 20913 15792 21655
rect 15750 20904 15806 20913
rect 15750 20839 15806 20848
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15672 18086 15700 19314
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 16454 15608 16526
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15212 14334 15332 14362
rect 15396 16102 15516 16130
rect 15212 13870 15240 14334
rect 15396 14226 15424 16102
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15488 15502 15516 15982
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15476 15360 15528 15366
rect 15474 15328 15476 15337
rect 15528 15328 15530 15337
rect 15474 15263 15530 15272
rect 15304 14198 15424 14226
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14660 12306 14688 12582
rect 14844 12306 14872 12786
rect 15212 12782 15240 13330
rect 15304 12986 15332 14198
rect 15580 13938 15608 15982
rect 15672 14521 15700 18022
rect 15764 16998 15792 20839
rect 15856 18737 15884 24074
rect 15948 21729 15976 24958
rect 16132 22710 16160 26302
rect 16394 26200 16450 26302
rect 17038 26330 17094 27000
rect 17038 26302 17356 26330
rect 17038 26200 17094 26302
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16302 24712 16358 24721
rect 16302 24647 16358 24656
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16212 22500 16264 22506
rect 16212 22442 16264 22448
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 15934 21720 15990 21729
rect 15934 21655 15990 21664
rect 15936 21616 15988 21622
rect 15934 21584 15936 21593
rect 15988 21584 15990 21593
rect 15934 21519 15990 21528
rect 16132 20602 16160 22170
rect 16224 21486 16252 22442
rect 16316 21690 16344 24647
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 16408 21010 16436 22170
rect 16592 21622 16620 23666
rect 16684 23118 16712 25094
rect 17132 24132 17184 24138
rect 17132 24074 17184 24080
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16776 23594 16804 24006
rect 17144 23730 17172 24074
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 16764 23588 16816 23594
rect 16764 23530 16816 23536
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16684 21690 16712 22646
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16776 22001 16804 22578
rect 16868 22574 16896 23054
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16762 21992 16818 22001
rect 16762 21927 16818 21936
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 16684 21434 16712 21626
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16592 21406 16712 21434
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 16026 19680 16082 19689
rect 16026 19615 16082 19624
rect 16040 19174 16068 19615
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 15842 18728 15898 18737
rect 15842 18663 15898 18672
rect 15936 18692 15988 18698
rect 15856 17882 15884 18663
rect 15936 18634 15988 18640
rect 15948 18290 15976 18634
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15948 17542 15976 18226
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15658 14512 15714 14521
rect 15658 14447 15714 14456
rect 15764 14464 15792 16594
rect 15856 14634 15884 17138
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15948 15706 15976 17070
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16040 15434 16068 19110
rect 16132 16266 16160 20266
rect 16592 20262 16620 21406
rect 16776 21332 16804 21558
rect 16684 21304 16804 21332
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16578 20088 16634 20097
rect 16578 20023 16634 20032
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16302 19136 16358 19145
rect 16302 19071 16358 19080
rect 16212 18828 16264 18834
rect 16316 18816 16344 19071
rect 16264 18788 16344 18816
rect 16212 18770 16264 18776
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16224 16454 16252 17818
rect 16316 17746 16344 18788
rect 16408 18630 16436 19654
rect 16592 19334 16620 20023
rect 16500 19306 16620 19334
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16500 18170 16528 19306
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16408 18154 16528 18170
rect 16396 18148 16528 18154
rect 16448 18142 16528 18148
rect 16396 18090 16448 18096
rect 16488 18080 16540 18086
rect 16486 18048 16488 18057
rect 16540 18048 16542 18057
rect 16486 17983 16542 17992
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 16658 16344 17478
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16132 16238 16252 16266
rect 16316 16250 16344 16594
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 15856 14606 16068 14634
rect 15936 14476 15988 14482
rect 15764 14436 15936 14464
rect 15936 14418 15988 14424
rect 15658 14376 15714 14385
rect 15658 14311 15714 14320
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15212 12345 15240 12378
rect 15198 12336 15254 12345
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14832 12300 14884 12306
rect 15198 12271 15254 12280
rect 14832 12242 14884 12248
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14568 11886 14688 11914
rect 14370 11863 14372 11872
rect 14424 11863 14426 11872
rect 14372 11834 14424 11840
rect 14278 11792 14334 11801
rect 14278 11727 14334 11736
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13924 11082 13952 11290
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13924 10742 13952 11018
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13726 10296 13782 10305
rect 13924 10266 13952 10678
rect 13726 10231 13782 10240
rect 13912 10260 13964 10266
rect 13740 9489 13768 10231
rect 13912 10202 13964 10208
rect 13924 9994 13952 10202
rect 14568 10130 14596 11018
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13924 9674 13952 9930
rect 14568 9674 14596 10066
rect 14660 10033 14688 11886
rect 14844 11830 14872 12038
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14936 11082 14964 12174
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15028 10266 15056 11018
rect 15304 10810 15332 11562
rect 15396 10810 15424 13806
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14646 10024 14702 10033
rect 14646 9959 14702 9968
rect 13832 9654 13952 9674
rect 13820 9648 13952 9654
rect 13872 9646 13952 9648
rect 14476 9646 14596 9674
rect 13820 9590 13872 9596
rect 14476 9518 14504 9646
rect 14464 9512 14516 9518
rect 13726 9480 13782 9489
rect 14464 9454 14516 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 13726 9415 13782 9424
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 14016 8634 14044 9318
rect 14752 8838 14780 9454
rect 15028 8974 15056 10202
rect 15212 10130 15240 10542
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9654 15240 9862
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 9042 15332 9454
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14752 8566 14780 8774
rect 15396 8634 15424 10610
rect 15672 9897 15700 14311
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15488 9042 15516 9658
rect 15764 9382 15792 13874
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15856 11830 15884 13194
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15856 11014 15884 11766
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15948 9110 15976 11698
rect 16040 10470 16068 14606
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16132 13190 16160 13806
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16224 12434 16252 16238
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16316 15094 16344 16186
rect 16408 16114 16436 17818
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16454 16528 16934
rect 16488 16448 16540 16454
rect 16592 16425 16620 18226
rect 16488 16390 16540 16396
rect 16578 16416 16634 16425
rect 16578 16351 16634 16360
rect 16684 16182 16712 21304
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16776 18834 16804 20742
rect 16868 19145 16896 22510
rect 16960 21865 16988 23666
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 16946 21856 17002 21865
rect 16946 21791 17002 21800
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 17144 20754 17172 21898
rect 17328 21486 17356 26302
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26330 21602 27000
rect 21546 26302 22048 26330
rect 21546 26200 21602 26302
rect 17590 24304 17646 24313
rect 17590 24239 17646 24248
rect 17604 24138 17632 24239
rect 17592 24132 17644 24138
rect 17512 24092 17592 24120
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17420 23662 17448 24006
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17420 23050 17448 23598
rect 17512 23050 17540 24092
rect 17592 24074 17644 24080
rect 17592 23588 17644 23594
rect 17592 23530 17644 23536
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17512 22438 17540 22986
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17316 21072 17368 21078
rect 17316 21014 17368 21020
rect 17328 20913 17356 21014
rect 17314 20904 17370 20913
rect 17314 20839 17370 20848
rect 16960 20602 16988 20742
rect 17144 20726 17356 20754
rect 17222 20632 17278 20641
rect 16948 20596 17000 20602
rect 17222 20567 17278 20576
rect 16948 20538 17000 20544
rect 17236 20534 17264 20567
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 17222 20360 17278 20369
rect 17222 20295 17278 20304
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17144 20058 17172 20198
rect 17236 20058 17264 20295
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16854 19136 16910 19145
rect 16854 19071 16910 19080
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16960 18766 16988 19246
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 17144 18630 17172 19382
rect 17328 19310 17356 20726
rect 17420 20330 17448 21898
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17512 20806 17540 21558
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 17512 19922 17540 20742
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17604 19802 17632 23530
rect 17696 22982 17724 26200
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23798 18368 26200
rect 18984 24410 19012 26200
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 18420 24336 18472 24342
rect 18420 24278 18472 24284
rect 18970 24304 19026 24313
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18432 23730 18460 24278
rect 18696 24268 18748 24274
rect 18970 24239 18972 24248
rect 18696 24210 18748 24216
rect 19024 24239 19026 24248
rect 18972 24210 19024 24216
rect 18708 23730 18736 24210
rect 19076 23798 19104 24686
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 19260 23798 19288 24210
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17880 23186 17908 23598
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 17972 23225 18000 23258
rect 17958 23216 18014 23225
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17868 23180 17920 23186
rect 17958 23151 18014 23160
rect 17868 23122 17920 23128
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17684 22704 17736 22710
rect 17788 22681 17816 23122
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17684 22646 17736 22652
rect 17774 22672 17830 22681
rect 17696 22438 17724 22646
rect 17774 22607 17830 22616
rect 17774 22536 17830 22545
rect 18432 22506 18460 23666
rect 18708 23526 18736 23666
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 19076 23254 19104 23734
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 17774 22471 17830 22480
rect 18420 22500 18472 22506
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17696 21962 17724 22374
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17788 21865 17816 22471
rect 18420 22442 18472 22448
rect 18524 22438 18552 22714
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 19156 22432 19208 22438
rect 19156 22374 19208 22380
rect 18524 22166 18552 22374
rect 18512 22160 18564 22166
rect 18512 22102 18564 22108
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17774 21856 17830 21865
rect 17774 21791 17830 21800
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17696 19922 17724 20742
rect 17774 20632 17830 20641
rect 17880 20618 17908 21898
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18696 21344 18748 21350
rect 18892 21332 18920 21966
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 18984 21690 19012 21830
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 19076 21622 19104 21830
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18748 21304 18920 21332
rect 18696 21286 18748 21292
rect 18602 21176 18658 21185
rect 18602 21111 18658 21120
rect 18616 21010 18644 21111
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17830 20590 17908 20618
rect 18512 20596 18564 20602
rect 17774 20567 17776 20576
rect 17828 20567 17830 20576
rect 17776 20538 17828 20544
rect 18512 20538 18564 20544
rect 18524 20233 18552 20538
rect 18510 20224 18566 20233
rect 18510 20159 18566 20168
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17512 19774 17632 19802
rect 18328 19780 18380 19786
rect 17406 19544 17462 19553
rect 17406 19479 17462 19488
rect 17316 19304 17368 19310
rect 17222 19272 17278 19281
rect 17316 19246 17368 19252
rect 17222 19207 17278 19216
rect 17236 18902 17264 19207
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17052 18340 17080 18566
rect 16960 18312 17080 18340
rect 16960 18222 16988 18312
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17377 16804 18022
rect 16762 17368 16818 17377
rect 16762 17303 16818 17312
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16408 14958 16436 15302
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 14482 16344 14758
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 13394 16436 14214
rect 16500 13394 16528 16118
rect 16776 15201 16804 16390
rect 16762 15192 16818 15201
rect 16868 15162 16896 18090
rect 16960 17746 16988 18158
rect 17144 18154 17172 18566
rect 17420 18306 17448 19479
rect 17512 19281 17540 19774
rect 18328 19722 18380 19728
rect 17592 19712 17644 19718
rect 17684 19712 17736 19718
rect 17592 19654 17644 19660
rect 17682 19680 17684 19689
rect 17868 19712 17920 19718
rect 17736 19680 17738 19689
rect 17498 19272 17554 19281
rect 17498 19207 17554 19216
rect 17328 18278 17448 18306
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17130 17776 17186 17785
rect 16948 17740 17000 17746
rect 17130 17711 17186 17720
rect 16948 17682 17000 17688
rect 16946 17640 17002 17649
rect 16946 17575 17002 17584
rect 16960 16969 16988 17575
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16946 16960 17002 16969
rect 16946 16895 17002 16904
rect 17052 15502 17080 17274
rect 17144 17202 17172 17711
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17236 16658 17264 17138
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17130 16280 17186 16289
rect 17130 16215 17132 16224
rect 17184 16215 17186 16224
rect 17132 16186 17184 16192
rect 17328 15586 17356 18278
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17512 18170 17540 19207
rect 17604 18290 17632 19654
rect 17868 19654 17920 19660
rect 17682 19615 17738 19624
rect 17682 19544 17738 19553
rect 17682 19479 17738 19488
rect 17880 19496 17908 19654
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17960 19508 18012 19514
rect 17696 19378 17724 19479
rect 17880 19468 17960 19496
rect 17960 19450 18012 19456
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17696 19145 17724 19178
rect 17788 19174 17816 19314
rect 17776 19168 17828 19174
rect 17682 19136 17738 19145
rect 17776 19110 17828 19116
rect 17682 19071 17738 19080
rect 18340 18902 18368 19722
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17774 18456 17830 18465
rect 17950 18459 18258 18468
rect 17684 18420 17736 18426
rect 17774 18391 17830 18400
rect 17684 18362 17736 18368
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17420 17082 17448 18158
rect 17512 18142 17632 18170
rect 17420 17054 17540 17082
rect 17512 16998 17540 17054
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17236 15558 17356 15586
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16762 15127 16818 15136
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16592 14414 16620 15030
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16592 14006 16620 14350
rect 16776 14074 16804 15030
rect 17052 14464 17080 15438
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 14929 17172 14962
rect 17130 14920 17186 14929
rect 17236 14890 17264 15558
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17130 14855 17186 14864
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17132 14476 17184 14482
rect 17052 14436 17132 14464
rect 17132 14418 17184 14424
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16592 13258 16620 13942
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16592 12986 16620 13194
rect 16960 12986 16988 13874
rect 17144 13870 17172 14418
rect 17328 14074 17356 15370
rect 17420 15366 17448 16934
rect 17604 16250 17632 18142
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17420 14346 17448 15302
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17144 13394 17172 13806
rect 17512 13734 17540 15914
rect 17604 15434 17632 16050
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17604 14482 17632 15370
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 14346 17632 14418
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17696 13852 17724 18362
rect 17788 17746 17816 18391
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 18068 18184 18158
rect 18328 18080 18380 18086
rect 18156 18040 18328 18068
rect 18328 18022 18380 18028
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17788 17134 17816 17274
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17788 15706 17816 16526
rect 17880 16250 17908 17274
rect 18340 17270 18368 17478
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17972 16522 18000 17002
rect 18236 16584 18288 16590
rect 18288 16544 18368 16572
rect 18236 16526 18288 16532
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18340 15094 18368 16544
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18432 15026 18460 19654
rect 18510 19544 18566 19553
rect 18510 19479 18566 19488
rect 18524 19378 18552 19479
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18708 19174 18736 20946
rect 18892 20806 18920 21304
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18892 20602 18920 20742
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 18800 19922 18828 20334
rect 18892 20262 18920 20334
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18984 19786 19012 21422
rect 19076 20942 19104 21422
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 19076 19514 19104 19790
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18510 18864 18566 18873
rect 18510 18799 18566 18808
rect 18524 17241 18552 18799
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18510 17232 18566 17241
rect 18510 17167 18566 17176
rect 18616 17105 18644 18702
rect 18696 18624 18748 18630
rect 18694 18592 18696 18601
rect 18748 18592 18750 18601
rect 18694 18527 18750 18536
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18892 17610 18920 18158
rect 18984 18057 19012 18158
rect 18970 18048 19026 18057
rect 18970 17983 19026 17992
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18602 17096 18658 17105
rect 18524 17054 18602 17082
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17776 13864 17828 13870
rect 17696 13824 17776 13852
rect 17776 13806 17828 13812
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13530 17540 13670
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17420 12850 17448 13466
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 16856 12776 16908 12782
rect 16578 12744 16634 12753
rect 16856 12718 16908 12724
rect 16578 12679 16634 12688
rect 16224 12406 16436 12434
rect 16212 12096 16264 12102
rect 16210 12064 16212 12073
rect 16264 12064 16266 12073
rect 16210 11999 16266 12008
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9722 16252 10066
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15856 8566 15884 8978
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12544 8486 12756 8514
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 12544 8362 12572 8486
rect 16040 8430 16068 9590
rect 16316 9382 16344 10542
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8906 16344 9318
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12452 5234 12480 7142
rect 12636 5846 12664 8366
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 8090 12848 8230
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 14200 7886 14228 8366
rect 16408 8294 16436 12406
rect 16592 12306 16620 12679
rect 16868 12646 16896 12718
rect 17512 12714 17540 13330
rect 17880 12866 17908 13330
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17880 12850 18000 12866
rect 17880 12844 18012 12850
rect 17880 12838 17960 12844
rect 17960 12786 18012 12792
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16592 11354 16620 12242
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 8362 16528 11018
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16592 8634 16620 10542
rect 16776 9518 16804 10678
rect 16868 10062 16896 11086
rect 17052 10810 17080 11630
rect 17236 11626 17264 12650
rect 17316 12300 17368 12306
rect 17368 12260 17448 12288
rect 17316 12242 17368 12248
rect 17420 11801 17448 12260
rect 17406 11792 17462 11801
rect 17406 11727 17408 11736
rect 17460 11727 17462 11736
rect 17408 11698 17460 11704
rect 17224 11620 17276 11626
rect 17224 11562 17276 11568
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17420 11082 17448 11290
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16868 9518 16896 9998
rect 17052 9994 17080 10746
rect 17512 10674 17540 12650
rect 17972 12442 18000 12786
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18144 12436 18196 12442
rect 18524 12434 18552 17054
rect 18602 17031 18658 17040
rect 18708 16250 18736 17478
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18786 16824 18842 16833
rect 18786 16759 18842 16768
rect 18880 16788 18932 16794
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18602 15192 18658 15201
rect 18602 15127 18658 15136
rect 18616 14822 18644 15127
rect 18604 14816 18656 14822
rect 18656 14776 18736 14804
rect 18604 14758 18656 14764
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18144 12378 18196 12384
rect 18432 12406 18552 12434
rect 18156 12238 18184 12378
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18432 12102 18460 12406
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18432 11830 18460 12038
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 16868 9042 16896 9454
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13372 7546 13400 7686
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12084 3466 12112 3674
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 11624 2582 11652 3334
rect 12636 3126 12664 5646
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13464 3466 13492 7686
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 5778 14044 7142
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 15212 4146 15240 7958
rect 16868 5778 16896 8978
rect 17236 8090 17264 9454
rect 17604 8838 17632 11630
rect 17788 10266 17816 11630
rect 18616 11354 18644 12718
rect 18708 11898 18736 14776
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18800 11830 18828 16759
rect 18880 16730 18932 16736
rect 18892 16182 18920 16730
rect 18984 16454 19012 17070
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 12918 18920 14962
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18892 12374 18920 12854
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18892 12102 18920 12310
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18604 11348 18656 11354
rect 18656 11308 18736 11336
rect 18604 11290 18656 11296
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10742 17908 11018
rect 18708 11014 18736 11308
rect 18892 11150 18920 12038
rect 18984 11354 19012 13194
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18892 9722 18920 10202
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18524 9450 18552 9590
rect 19076 9450 19104 19314
rect 19168 16114 19196 22374
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 14482 19196 14758
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19168 13530 19196 14418
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19168 13326 19196 13466
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19168 12442 19196 13262
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19260 12186 19288 22578
rect 19352 20058 19380 24074
rect 19628 23254 19656 26200
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19798 23624 19854 23633
rect 19798 23559 19854 23568
rect 19432 23248 19484 23254
rect 19430 23216 19432 23225
rect 19616 23248 19668 23254
rect 19484 23216 19486 23225
rect 19616 23190 19668 23196
rect 19430 23151 19486 23160
rect 19614 22808 19670 22817
rect 19614 22743 19670 22752
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19444 22098 19472 22578
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19444 21350 19472 22034
rect 19628 22030 19656 22743
rect 19812 22438 19840 23559
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 20942 19472 21286
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20602 19472 20878
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19352 19514 19380 19722
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19444 17746 19472 19382
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19432 16584 19484 16590
rect 19338 16552 19394 16561
rect 19432 16526 19484 16532
rect 19338 16487 19394 16496
rect 19352 15366 19380 16487
rect 19444 16114 19472 16526
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19338 14920 19394 14929
rect 19338 14855 19394 14864
rect 19352 14822 19380 14855
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19168 12158 19288 12186
rect 19168 11558 19196 12158
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 18524 8838 18552 9386
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 12084 800 12112 2450
rect 12452 2446 12480 2858
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14752 800 14780 2450
rect 15028 2446 15056 3878
rect 15488 3126 15516 5102
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 17052 3058 17080 5510
rect 17420 4826 17448 5578
rect 17512 5234 17540 7142
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18524 5710 18552 8774
rect 19260 7954 19288 9930
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19352 6866 19380 14758
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19444 13433 19472 14282
rect 19536 13977 19564 19994
rect 19628 15502 19656 21626
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 21010 19748 21286
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19720 20777 19748 20810
rect 19706 20768 19762 20777
rect 19706 20703 19762 20712
rect 19812 20097 19840 21898
rect 19798 20088 19854 20097
rect 19798 20023 19854 20032
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19720 19310 19748 19790
rect 19904 19786 19932 24210
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19720 18834 19748 19246
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19720 18154 19748 18634
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19720 16794 19748 17614
rect 19812 17513 19840 18158
rect 19892 17536 19944 17542
rect 19798 17504 19854 17513
rect 19892 17478 19944 17484
rect 19798 17439 19854 17448
rect 19904 16998 19932 17478
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19996 16522 20024 24142
rect 20166 23896 20222 23905
rect 20166 23831 20222 23840
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23186 20116 23462
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20088 22710 20116 23122
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 20180 22556 20208 23831
rect 20088 22528 20208 22556
rect 20088 18850 20116 22528
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 20180 21418 20208 22374
rect 20272 22234 20300 26200
rect 20810 24304 20866 24313
rect 20916 24274 20944 26200
rect 21560 24954 21956 24970
rect 21560 24948 21968 24954
rect 21560 24942 21916 24948
rect 21560 24886 21588 24942
rect 21916 24890 21968 24896
rect 21548 24880 21600 24886
rect 21178 24848 21234 24857
rect 21548 24822 21600 24828
rect 21178 24783 21234 24792
rect 20810 24239 20812 24248
rect 20864 24239 20866 24248
rect 20904 24268 20956 24274
rect 20812 24210 20864 24216
rect 20904 24210 20956 24216
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20364 22778 20392 22986
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20456 22094 20484 24006
rect 21192 23798 21220 24783
rect 21732 24608 21784 24614
rect 21732 24550 21784 24556
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21638 24440 21694 24449
rect 21638 24375 21694 24384
rect 21180 23792 21232 23798
rect 21180 23734 21232 23740
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20364 22066 20484 22094
rect 20364 22030 20392 22066
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20272 21622 20300 21966
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20168 21412 20220 21418
rect 20168 21354 20220 21360
rect 20088 18822 20208 18850
rect 20074 17912 20130 17921
rect 20074 17847 20130 17856
rect 20088 17270 20116 17847
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19890 16144 19946 16153
rect 20088 16114 20116 16730
rect 19890 16079 19946 16088
rect 20076 16108 20128 16114
rect 19904 15638 19932 16079
rect 20076 16050 20128 16056
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 20088 15570 20116 16050
rect 20180 15910 20208 18822
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18290 20300 18566
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20272 16810 20300 18226
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20364 16998 20392 17070
rect 20352 16992 20404 16998
rect 20350 16960 20352 16969
rect 20404 16960 20406 16969
rect 20350 16895 20406 16904
rect 20272 16782 20392 16810
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 20260 15428 20312 15434
rect 20260 15370 20312 15376
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19522 13968 19578 13977
rect 19522 13903 19578 13912
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19430 13424 19486 13433
rect 19430 13359 19486 13368
rect 19536 13326 19564 13466
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 11762 19472 12582
rect 19720 12170 19748 14962
rect 20168 14952 20220 14958
rect 20166 14920 20168 14929
rect 20220 14920 20222 14929
rect 19984 14884 20036 14890
rect 20166 14855 20222 14864
rect 19984 14826 20036 14832
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19720 11082 19748 11630
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 10606 19748 11018
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10130 19748 10542
rect 19812 10266 19840 14418
rect 19996 13870 20024 14826
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 12986 20208 13670
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20088 12306 20116 12718
rect 20272 12345 20300 15370
rect 20364 15201 20392 16782
rect 20456 16658 20484 17614
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20350 15192 20406 15201
rect 20350 15127 20406 15136
rect 20548 14822 20576 22918
rect 20640 22574 20668 23462
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20640 19310 20668 20334
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20732 17082 20760 23666
rect 21548 22500 21600 22506
rect 21548 22442 21600 22448
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21284 22030 21312 22170
rect 21560 22098 21588 22442
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 21008 21350 21036 21558
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21008 20874 21036 21286
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21192 19922 21220 20742
rect 21548 19984 21600 19990
rect 21376 19932 21548 19938
rect 21376 19926 21600 19932
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21376 19910 21588 19926
rect 21376 19553 21404 19910
rect 21548 19848 21600 19854
rect 21468 19808 21548 19836
rect 21362 19544 21418 19553
rect 21362 19479 21418 19488
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21100 18612 21128 18838
rect 21100 18584 21220 18612
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 21008 17746 21036 18090
rect 21100 17814 21128 18226
rect 21192 18222 21220 18584
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20996 17740 21048 17746
rect 20996 17682 21048 17688
rect 20994 17640 21050 17649
rect 20994 17575 21050 17584
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20732 17054 20852 17082
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16658 20760 16934
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20824 15722 20852 17054
rect 20916 15745 20944 17206
rect 20732 15694 20852 15722
rect 20902 15736 20958 15745
rect 20732 15178 20760 15694
rect 20902 15671 20958 15680
rect 20640 15150 20760 15178
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20258 12336 20314 12345
rect 20076 12300 20128 12306
rect 20258 12271 20314 12280
rect 20076 12242 20128 12248
rect 20364 12170 20392 13126
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 20364 8430 20392 12106
rect 20456 8498 20484 13874
rect 20548 10470 20576 14214
rect 20640 14074 20668 15150
rect 21008 15026 21036 17575
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 21100 16522 21128 17002
rect 21088 16516 21140 16522
rect 21088 16458 21140 16464
rect 21100 15570 21128 16458
rect 21192 16250 21220 18158
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21272 15904 21324 15910
rect 21270 15872 21272 15881
rect 21324 15872 21326 15881
rect 21270 15807 21326 15816
rect 21088 15564 21140 15570
rect 21140 15524 21220 15552
rect 21088 15506 21140 15512
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20640 11257 20668 12854
rect 20732 12442 20760 13738
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13530 21036 13670
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21100 12986 21128 14010
rect 21192 13258 21220 15524
rect 21376 14550 21404 19479
rect 21468 18834 21496 19808
rect 21548 19790 21600 19796
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21454 18456 21510 18465
rect 21454 18391 21456 18400
rect 21508 18391 21510 18400
rect 21456 18362 21508 18368
rect 21560 16998 21588 18770
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21468 14906 21496 16186
rect 21560 15094 21588 16390
rect 21652 16046 21680 24375
rect 21744 24206 21772 24550
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21928 23866 21956 24550
rect 22020 24256 22048 26302
rect 22190 26200 22246 27000
rect 22834 26330 22890 27000
rect 23388 26376 23440 26382
rect 22834 26302 23336 26330
rect 23478 26330 23534 27000
rect 23440 26324 23534 26330
rect 23388 26318 23534 26324
rect 23400 26302 23534 26318
rect 22834 26200 22890 26302
rect 22100 24268 22152 24274
rect 22020 24228 22100 24256
rect 22100 24210 22152 24216
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21836 22982 21864 23666
rect 22100 23520 22152 23526
rect 21914 23488 21970 23497
rect 22204 23497 22232 26200
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22282 23896 22338 23905
rect 23308 23882 23336 26302
rect 23478 26200 23534 26302
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26330 25466 27000
rect 24964 26302 25466 26330
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 23308 23854 23428 23882
rect 22282 23831 22338 23840
rect 22296 23633 22324 23831
rect 22376 23656 22428 23662
rect 22282 23624 22338 23633
rect 22376 23598 22428 23604
rect 22282 23559 22338 23568
rect 22100 23462 22152 23468
rect 22190 23488 22246 23497
rect 21914 23423 21970 23432
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21836 22409 21864 22918
rect 21822 22400 21878 22409
rect 21822 22335 21878 22344
rect 21928 22250 21956 23423
rect 22112 23050 22140 23462
rect 22190 23423 22246 23432
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 22112 22438 22140 22986
rect 22296 22642 22324 23054
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22296 22506 22324 22578
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 21928 22222 22232 22250
rect 22008 22160 22060 22166
rect 22008 22102 22060 22108
rect 22020 21894 22048 22102
rect 22204 22030 22232 22222
rect 22388 22094 22416 23598
rect 22836 23520 22888 23526
rect 22836 23462 22888 23468
rect 22742 23352 22798 23361
rect 22742 23287 22798 23296
rect 22756 22953 22784 23287
rect 22742 22944 22798 22953
rect 22742 22879 22798 22888
rect 22848 22642 22876 23462
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22296 22066 22416 22094
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21928 21350 21956 21422
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21824 20868 21876 20874
rect 21824 20810 21876 20816
rect 21836 20262 21864 20810
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21928 20534 21956 20742
rect 21916 20528 21968 20534
rect 21916 20470 21968 20476
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21928 19786 21956 20470
rect 22112 20466 22140 21830
rect 22296 21078 22324 22066
rect 22848 21690 22876 22578
rect 23216 22522 23244 22918
rect 23400 22522 23428 23854
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 23254 23796 23462
rect 23756 23248 23808 23254
rect 23756 23190 23808 23196
rect 23860 23050 23888 23802
rect 23848 23044 23900 23050
rect 23848 22986 23900 22992
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 23480 22568 23532 22574
rect 23124 22506 23336 22522
rect 23112 22500 23336 22506
rect 23164 22494 23336 22500
rect 23400 22516 23480 22522
rect 23400 22510 23532 22516
rect 23400 22494 23520 22510
rect 23112 22442 23164 22448
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22234 23336 22494
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 23676 22030 23704 22646
rect 23860 22438 23888 22986
rect 23952 22681 23980 24142
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 23938 22672 23994 22681
rect 23938 22607 23994 22616
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23754 22264 23810 22273
rect 23754 22199 23810 22208
rect 23768 22166 23796 22199
rect 23756 22160 23808 22166
rect 23756 22102 23808 22108
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23296 21888 23348 21894
rect 23294 21856 23296 21865
rect 23348 21856 23350 21865
rect 23294 21791 23350 21800
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22376 21412 22428 21418
rect 22376 21354 22428 21360
rect 22284 21072 22336 21078
rect 22284 21014 22336 21020
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 21916 19780 21968 19786
rect 21916 19722 21968 19728
rect 21928 19378 21956 19722
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21928 17542 21956 19314
rect 22112 19242 22140 20402
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22020 18970 22048 19178
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22112 18630 22140 19178
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21822 17232 21878 17241
rect 21822 17167 21878 17176
rect 21836 17066 21864 17167
rect 21916 17128 21968 17134
rect 21914 17096 21916 17105
rect 21968 17096 21970 17105
rect 21824 17060 21876 17066
rect 21914 17031 21970 17040
rect 21824 17002 21876 17008
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21652 15706 21680 15982
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21468 14878 21588 14906
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21376 14385 21404 14486
rect 21362 14376 21418 14385
rect 21362 14311 21418 14320
rect 21376 14278 21404 14311
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 14006 21404 14214
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21192 12986 21220 13194
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 21088 12164 21140 12170
rect 21192 12152 21220 12922
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21140 12124 21220 12152
rect 21088 12106 21140 12112
rect 21192 11694 21220 12124
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21468 11558 21496 12718
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 20626 11248 20682 11257
rect 20626 11183 20682 11192
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9382 20760 9998
rect 21192 9926 21220 11018
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 10538 21404 10950
rect 21468 10810 21496 11494
rect 21560 11218 21588 14878
rect 21744 14550 21772 16934
rect 21836 15094 21864 17002
rect 21914 16824 21970 16833
rect 21914 16759 21970 16768
rect 21928 16425 21956 16759
rect 22020 16726 22048 17614
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 21914 16416 21970 16425
rect 21914 16351 21970 16360
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21652 13462 21680 13874
rect 21836 13530 21864 15030
rect 21928 14890 21956 15302
rect 22020 15026 22048 16662
rect 22112 15570 22140 18566
rect 22204 15994 22232 20198
rect 22296 19854 22324 21014
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22296 17270 22324 17750
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22388 16114 22416 21354
rect 22480 21146 22508 21422
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22664 20890 22692 20946
rect 22664 20862 22784 20890
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22480 20602 22508 20742
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22572 20330 22600 20742
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22664 19446 22692 20742
rect 22756 19990 22784 20862
rect 23400 20466 23428 21490
rect 23584 20874 23612 21966
rect 23952 21622 23980 22374
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23572 20868 23624 20874
rect 23572 20810 23624 20816
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 20641 23704 20742
rect 23662 20632 23718 20641
rect 23662 20567 23718 20576
rect 23756 20596 23808 20602
rect 23756 20538 23808 20544
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 23768 19854 23796 20538
rect 23860 19922 23888 20946
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22572 18970 22600 19246
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22664 17202 22692 18362
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22204 15966 22324 15994
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22112 15162 22140 15506
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21928 14346 21956 14826
rect 22020 14482 22048 14962
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 22204 13546 22232 15846
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 22112 13518 22232 13546
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 22112 12850 22140 13518
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22204 12850 22232 13330
rect 22296 12889 22324 15966
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22388 15366 22416 15438
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22374 13968 22430 13977
rect 22374 13903 22376 13912
rect 22428 13903 22430 13912
rect 22376 13874 22428 13880
rect 22388 13530 22416 13874
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22282 12880 22338 12889
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22192 12844 22244 12850
rect 22282 12815 22338 12824
rect 22192 12786 22244 12792
rect 22204 12238 22232 12786
rect 22480 12714 22508 16390
rect 22572 13734 22600 17070
rect 22664 16833 22692 17138
rect 22650 16824 22706 16833
rect 22650 16759 22706 16768
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22664 15434 22692 16594
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22756 14362 22784 19722
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23308 19514 23336 19654
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22848 15978 22876 19314
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23386 18728 23442 18737
rect 22928 18692 22980 18698
rect 23386 18663 23442 18672
rect 22928 18634 22980 18640
rect 22940 18426 22968 18634
rect 23400 18630 23428 18663
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 23032 18358 23060 18566
rect 23492 18426 23520 19110
rect 23584 18766 23612 19110
rect 23676 18834 23704 19654
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23020 18352 23072 18358
rect 23020 18294 23072 18300
rect 23386 18048 23442 18057
rect 22950 17980 23258 17989
rect 23386 17983 23442 17992
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23400 17354 23428 17983
rect 23480 17536 23532 17542
rect 23676 17513 23704 18566
rect 23768 18465 23796 19654
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23754 18456 23810 18465
rect 23754 18391 23810 18400
rect 23860 18358 23888 18634
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23860 17610 23888 18294
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23480 17478 23532 17484
rect 23662 17504 23718 17513
rect 23124 17326 23428 17354
rect 23124 17270 23152 17326
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16590 23336 16934
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22664 14334 22784 14362
rect 22664 14278 22692 14334
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22650 13968 22706 13977
rect 22650 13903 22706 13912
rect 22664 13870 22692 13903
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22204 11694 22232 12174
rect 22756 11830 22784 14214
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21560 10266 21588 10678
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21560 10062 21588 10202
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21192 9518 21220 9862
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 22204 7410 22232 11630
rect 22848 11354 22876 13806
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 13530 23336 15438
rect 23400 15178 23428 16458
rect 23492 15366 23520 17478
rect 23662 17439 23718 17448
rect 23676 17116 23704 17439
rect 23952 17338 23980 20742
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 23846 17232 23902 17241
rect 24044 17218 24072 24006
rect 24136 23322 24164 26200
rect 24124 23316 24176 23322
rect 24124 23258 24176 23264
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24136 21350 24164 22918
rect 24412 22166 24440 23258
rect 24492 23044 24544 23050
rect 24492 22986 24544 22992
rect 24504 22642 24532 22986
rect 24780 22953 24808 26200
rect 24964 24206 24992 26302
rect 25410 26200 25466 26302
rect 26054 26330 26110 27000
rect 26698 26330 26754 27000
rect 27342 26330 27398 27000
rect 27986 26330 28042 27000
rect 26054 26302 26188 26330
rect 26054 26200 26110 26302
rect 26160 24936 26188 26302
rect 26698 26302 27016 26330
rect 26698 26200 26754 26302
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26160 24908 26280 24936
rect 26252 24818 26280 24908
rect 26148 24812 26200 24818
rect 26148 24754 26200 24760
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 25780 24676 25832 24682
rect 25780 24618 25832 24624
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 25792 24410 25820 24618
rect 25136 24404 25188 24410
rect 25780 24404 25832 24410
rect 25188 24364 25268 24392
rect 25136 24346 25188 24352
rect 25240 24274 25268 24364
rect 25780 24346 25832 24352
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 26068 24206 26096 24618
rect 26160 24206 26188 24754
rect 26424 24744 26476 24750
rect 26424 24686 26476 24692
rect 26436 24274 26464 24686
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 24964 23866 24992 24006
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25780 23860 25832 23866
rect 25780 23802 25832 23808
rect 25412 23792 25464 23798
rect 25412 23734 25464 23740
rect 25424 23497 25452 23734
rect 25410 23488 25466 23497
rect 25410 23423 25466 23432
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 24952 22976 25004 22982
rect 24766 22944 24822 22953
rect 24952 22918 25004 22924
rect 24766 22879 24822 22888
rect 24964 22817 24992 22918
rect 24950 22808 25006 22817
rect 25148 22778 25176 23122
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 24950 22743 25006 22752
rect 25136 22772 25188 22778
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24400 22160 24452 22166
rect 24400 22102 24452 22108
rect 24308 21888 24360 21894
rect 24308 21830 24360 21836
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24216 20936 24268 20942
rect 24216 20878 24268 20884
rect 24228 20466 24256 20878
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24124 19168 24176 19174
rect 24124 19110 24176 19116
rect 24136 18766 24164 19110
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24214 18592 24270 18601
rect 24214 18527 24270 18536
rect 24228 17338 24256 18527
rect 24320 17785 24348 21830
rect 24504 21690 24532 22578
rect 24688 22030 24716 22646
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24492 21684 24544 21690
rect 24964 21672 24992 22743
rect 25136 22714 25188 22720
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25044 21684 25096 21690
rect 24964 21644 25044 21672
rect 24492 21626 24544 21632
rect 25044 21626 25096 21632
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24688 20398 24716 21422
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24780 21078 24808 21354
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 24306 17776 24362 17785
rect 24306 17711 24362 17720
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24044 17190 24164 17218
rect 23846 17167 23902 17176
rect 23860 17134 23888 17167
rect 23756 17128 23808 17134
rect 23676 17088 23756 17116
rect 23756 17070 23808 17076
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 23768 16794 23796 17070
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23846 16688 23902 16697
rect 23756 16652 23808 16658
rect 23846 16623 23902 16632
rect 23756 16594 23808 16600
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23676 16114 23704 16526
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23400 15150 23520 15178
rect 23584 15162 23612 15370
rect 23492 14906 23520 15150
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23400 14878 23520 14906
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23032 12850 23060 13262
rect 23308 13240 23336 13466
rect 23400 13462 23428 14878
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23388 13252 23440 13258
rect 23308 13212 23388 13240
rect 23388 13194 23440 13200
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23124 12986 23152 13126
rect 23492 12986 23520 13330
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23584 12918 23612 13330
rect 23572 12912 23624 12918
rect 23572 12854 23624 12860
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 23676 12782 23704 14486
rect 23768 13870 23796 16594
rect 23860 16454 23888 16623
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23860 16046 23888 16390
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23860 15162 23888 15302
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23860 14346 23888 15098
rect 23952 15026 23980 15370
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23952 14482 23980 14962
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23848 14340 23900 14346
rect 23900 14300 23980 14328
rect 23848 14282 23900 14288
rect 23848 14000 23900 14006
rect 23846 13968 23848 13977
rect 23900 13968 23902 13977
rect 23846 13903 23902 13912
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23860 13462 23888 13903
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23952 12918 23980 14300
rect 24044 13870 24072 15982
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 23952 12782 23980 12854
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23952 12238 23980 12718
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 23952 11830 23980 12174
rect 24044 12102 24072 13806
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11898 24072 12038
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22296 10810 22324 11086
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22848 10606 22876 11290
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23400 9994 23428 11494
rect 23952 11354 23980 11766
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23400 7750 23428 9454
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17420 2990 17448 4762
rect 17696 4486 17724 5102
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 3126 17724 4422
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17880 3058 17908 4966
rect 20272 4826 20300 5646
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20272 4622 20300 4762
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 20548 3058 20576 4966
rect 20732 3466 20760 6802
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21744 5846 21772 6734
rect 22480 5914 22508 7278
rect 22848 6458 22876 7686
rect 23584 7410 23612 11290
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23768 6934 23796 9522
rect 24136 9081 24164 17190
rect 24228 16590 24256 17274
rect 24412 17202 24440 17478
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24504 16590 24532 19314
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24688 17746 24716 18022
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24596 17134 24624 17682
rect 24688 17202 24716 17682
rect 24872 17218 24900 19246
rect 24950 18456 25006 18465
rect 24950 18391 25006 18400
rect 24964 17354 24992 18391
rect 25056 18290 25084 19314
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25148 18329 25176 18566
rect 25134 18320 25190 18329
rect 25044 18284 25096 18290
rect 25134 18255 25190 18264
rect 25044 18226 25096 18232
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 24964 17326 25084 17354
rect 24676 17196 24728 17202
rect 24872 17190 24992 17218
rect 24728 17156 24808 17184
rect 24676 17138 24728 17144
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24596 16454 24624 16934
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24596 16114 24624 16390
rect 24584 16108 24636 16114
rect 24780 16096 24808 17156
rect 24964 16250 24992 17190
rect 25056 16998 25084 17326
rect 25148 16998 25176 17546
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24860 16108 24912 16114
rect 24780 16068 24860 16096
rect 24584 16050 24636 16056
rect 24860 16050 24912 16056
rect 24596 15706 24624 16050
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24964 15162 24992 16186
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 25056 14482 25084 16594
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25148 14929 25176 16390
rect 25240 15910 25268 21286
rect 25332 21146 25360 22374
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25332 19446 25360 20946
rect 25424 20777 25452 22918
rect 25792 22778 25820 23802
rect 26068 22982 26096 24006
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 26148 23656 26200 23662
rect 26148 23598 26200 23604
rect 26160 23254 26188 23598
rect 26148 23248 26200 23254
rect 26148 23190 26200 23196
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 26436 22574 26464 23734
rect 26608 23520 26660 23526
rect 26792 23520 26844 23526
rect 26608 23462 26660 23468
rect 26790 23488 26792 23497
rect 26844 23488 26846 23497
rect 26620 23322 26648 23462
rect 26790 23423 26846 23432
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 26516 22976 26568 22982
rect 26516 22918 26568 22924
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 25872 22568 25924 22574
rect 25700 22516 25872 22522
rect 25700 22510 25924 22516
rect 26424 22568 26476 22574
rect 26424 22510 26476 22516
rect 25700 22506 25912 22510
rect 25688 22500 25912 22506
rect 25740 22494 25912 22500
rect 25688 22442 25740 22448
rect 26528 22438 26556 22918
rect 26804 22642 26832 22918
rect 26792 22636 26844 22642
rect 26792 22578 26844 22584
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 26528 22273 26556 22374
rect 26514 22264 26570 22273
rect 26240 22228 26292 22234
rect 26292 22188 26372 22216
rect 26514 22199 26570 22208
rect 26240 22170 26292 22176
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25688 21616 25740 21622
rect 25688 21558 25740 21564
rect 25410 20768 25466 20777
rect 25410 20703 25466 20712
rect 25700 20466 25728 21558
rect 25792 20942 25820 21966
rect 26344 21962 26372 22188
rect 26700 22092 26752 22098
rect 26700 22034 26752 22040
rect 26792 22094 26844 22098
rect 26896 22094 26924 25638
rect 26988 24070 27016 26302
rect 27342 26302 27568 26330
rect 27342 26200 27398 26302
rect 27252 24744 27304 24750
rect 27158 24712 27214 24721
rect 27252 24686 27304 24692
rect 27158 24647 27214 24656
rect 27172 24410 27200 24647
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27068 23316 27120 23322
rect 27068 23258 27120 23264
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 26792 22092 26924 22094
rect 26844 22066 26924 22092
rect 26792 22034 26844 22040
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25976 21554 26004 21830
rect 25964 21548 26016 21554
rect 25964 21490 26016 21496
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26252 21321 26280 21422
rect 26238 21312 26294 21321
rect 26238 21247 26294 21256
rect 26344 21146 26372 21898
rect 26712 21486 26740 22034
rect 26700 21480 26752 21486
rect 26700 21422 26752 21428
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26068 20602 26096 20878
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25700 20262 25728 20402
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25596 19780 25648 19786
rect 25596 19722 25648 19728
rect 25320 19440 25372 19446
rect 25320 19382 25372 19388
rect 25608 16590 25636 19722
rect 25700 19514 25728 20198
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25792 19310 25820 19790
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25792 18834 25820 19246
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25792 17746 25820 18770
rect 25976 18698 26004 20334
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 26068 18358 26096 20538
rect 26148 19916 26200 19922
rect 26148 19858 26200 19864
rect 26160 19224 26188 19858
rect 26252 19514 26280 20810
rect 26606 20632 26662 20641
rect 26606 20567 26608 20576
rect 26660 20567 26662 20576
rect 26608 20538 26660 20544
rect 26424 19780 26476 19786
rect 26424 19722 26476 19728
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26160 19196 26280 19224
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 26252 18222 26280 19196
rect 26436 18834 26464 19722
rect 26804 19666 26832 22034
rect 26988 22012 27016 22510
rect 27080 22386 27108 23258
rect 27172 23186 27200 23598
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 27264 22574 27292 24686
rect 27540 23662 27568 26302
rect 27986 26302 28488 26330
rect 27986 26200 28042 26302
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27344 23316 27396 23322
rect 27632 23304 27660 24278
rect 27712 24132 27764 24138
rect 27712 24074 27764 24080
rect 27396 23276 27660 23304
rect 27344 23258 27396 23264
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27632 22710 27660 23122
rect 27528 22704 27580 22710
rect 27434 22672 27490 22681
rect 27528 22646 27580 22652
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27434 22607 27436 22616
rect 27488 22607 27490 22616
rect 27436 22578 27488 22584
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27344 22500 27396 22506
rect 27344 22442 27396 22448
rect 27356 22386 27384 22442
rect 27080 22358 27384 22386
rect 27066 22264 27122 22273
rect 27122 22222 27200 22250
rect 27356 22234 27384 22358
rect 27066 22199 27122 22208
rect 27068 22024 27120 22030
rect 26988 21984 27068 22012
rect 27068 21966 27120 21972
rect 26804 19638 26924 19666
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26804 18766 26832 19450
rect 26896 19310 26924 19638
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 26804 18426 26832 18702
rect 27068 18692 27120 18698
rect 26988 18652 27068 18680
rect 26792 18420 26844 18426
rect 26792 18362 26844 18368
rect 26240 18216 26292 18222
rect 26240 18158 26292 18164
rect 26252 17814 26280 18158
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25686 17640 25742 17649
rect 26804 17610 26832 18362
rect 25686 17575 25742 17584
rect 26792 17604 26844 17610
rect 25700 16726 25728 17575
rect 26792 17546 26844 17552
rect 26804 17270 26832 17546
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 26792 17264 26844 17270
rect 26792 17206 26844 17212
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25976 16726 26004 16934
rect 25688 16720 25740 16726
rect 25688 16662 25740 16668
rect 25964 16720 26016 16726
rect 25964 16662 26016 16668
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25424 15434 25452 16118
rect 25792 15570 25820 16594
rect 25884 16454 25912 16594
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 26252 16114 26280 17206
rect 26988 16658 27016 18652
rect 27068 18634 27120 18640
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 27080 16658 27108 18158
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26976 15632 27028 15638
rect 26976 15574 27028 15580
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25412 15428 25464 15434
rect 25412 15370 25464 15376
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25134 14920 25190 14929
rect 25134 14855 25190 14864
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24596 14006 24624 14214
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 25056 13988 25084 14418
rect 25148 14346 25176 14855
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25136 14000 25188 14006
rect 25056 13960 25136 13988
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24504 12442 24532 12718
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24596 9654 24624 13670
rect 25056 12170 25084 13960
rect 25136 13942 25188 13948
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 25148 11558 25176 13806
rect 25240 13190 25268 15302
rect 25608 15201 25636 15438
rect 25594 15192 25650 15201
rect 25594 15127 25650 15136
rect 25792 14550 25820 15506
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 25780 14544 25832 14550
rect 25780 14486 25832 14492
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25792 14074 25820 14214
rect 25884 14074 25912 14282
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 26160 13297 26188 14894
rect 26344 14346 26372 15370
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26620 14482 26648 14758
rect 26988 14618 27016 15574
rect 27080 15162 27108 16050
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 26896 14074 26924 14554
rect 26988 14414 27016 14554
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 26146 13288 26202 13297
rect 26146 13223 26202 13232
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 25228 13184 25280 13190
rect 25228 13126 25280 13132
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 26896 11218 26924 13194
rect 27172 12434 27200 22222
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27448 22094 27476 22578
rect 27540 22273 27568 22646
rect 27526 22264 27582 22273
rect 27526 22199 27582 22208
rect 27264 22066 27476 22094
rect 27724 22080 27752 24074
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 28368 22982 28396 24006
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 28460 22778 28488 26302
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29918 26330 29974 27000
rect 29918 26302 30144 26330
rect 29918 26200 29974 26302
rect 28540 25152 28592 25158
rect 28540 25094 28592 25100
rect 28552 23882 28580 25094
rect 28644 24052 28672 26200
rect 29184 24812 29236 24818
rect 29184 24754 29236 24760
rect 29092 24404 29144 24410
rect 29092 24346 29144 24352
rect 29104 24154 29132 24346
rect 29196 24206 29224 24754
rect 29288 24274 29316 26200
rect 30012 24608 30064 24614
rect 30012 24550 30064 24556
rect 30024 24274 30052 24550
rect 29276 24268 29328 24274
rect 29276 24210 29328 24216
rect 30012 24268 30064 24274
rect 30012 24210 30064 24216
rect 29012 24126 29132 24154
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 28644 24024 28856 24052
rect 28552 23854 28672 23882
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28552 23118 28580 23666
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28264 22432 28316 22438
rect 28264 22374 28316 22380
rect 27264 20466 27292 22066
rect 27632 22052 27752 22080
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27356 20874 27384 21966
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27540 21078 27568 21626
rect 27528 21072 27580 21078
rect 27528 21014 27580 21020
rect 27344 20868 27396 20874
rect 27344 20810 27396 20816
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27252 20256 27304 20262
rect 27356 20244 27384 20810
rect 27528 20596 27580 20602
rect 27632 20584 27660 22052
rect 28276 22030 28304 22374
rect 28356 22228 28408 22234
rect 28356 22170 28408 22176
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28368 21486 28396 22170
rect 28644 22094 28672 23854
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 28736 23322 28764 23462
rect 28724 23316 28776 23322
rect 28724 23258 28776 23264
rect 28736 22574 28764 23258
rect 28828 23050 28856 24024
rect 29012 23322 29040 24126
rect 29092 24064 29144 24070
rect 29092 24006 29144 24012
rect 29000 23316 29052 23322
rect 29000 23258 29052 23264
rect 28816 23044 28868 23050
rect 28816 22986 28868 22992
rect 28908 22976 28960 22982
rect 28908 22918 28960 22924
rect 28920 22710 28948 22918
rect 28908 22704 28960 22710
rect 28908 22646 28960 22652
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 29000 22160 29052 22166
rect 28552 22066 28672 22094
rect 28920 22108 29000 22114
rect 28920 22102 29052 22108
rect 28920 22086 29040 22102
rect 28448 21888 28500 21894
rect 28448 21830 28500 21836
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 27816 21010 27844 21422
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 27580 20556 27660 20584
rect 27528 20538 27580 20544
rect 27632 20466 27660 20556
rect 27712 20528 27764 20534
rect 27712 20470 27764 20476
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27304 20216 27384 20244
rect 27252 20198 27304 20204
rect 27264 19854 27292 20198
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27264 19514 27292 19790
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 27632 19334 27660 20402
rect 27724 19514 27752 20470
rect 27816 19990 27844 20946
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28368 20466 28396 21422
rect 28460 21350 28488 21830
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28552 21010 28580 22066
rect 28724 21480 28776 21486
rect 28724 21422 28776 21428
rect 28736 21321 28764 21422
rect 28722 21312 28778 21321
rect 28722 21247 28778 21256
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 28540 21004 28592 21010
rect 28540 20946 28592 20952
rect 28448 20936 28500 20942
rect 28500 20884 28580 20890
rect 28448 20878 28580 20884
rect 28460 20862 28580 20878
rect 28446 20768 28502 20777
rect 28446 20703 28502 20712
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 27804 19984 27856 19990
rect 27804 19926 27856 19932
rect 28460 19854 28488 20703
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28000 19718 28028 19790
rect 27988 19712 28040 19718
rect 27988 19654 28040 19660
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27804 19508 27856 19514
rect 27804 19450 27856 19456
rect 27816 19334 27844 19450
rect 27436 19304 27488 19310
rect 27632 19306 27844 19334
rect 27434 19272 27436 19281
rect 27488 19272 27490 19281
rect 27434 19207 27490 19216
rect 27816 19174 27844 19306
rect 28264 19304 28316 19310
rect 28316 19264 28396 19292
rect 28264 19246 28316 19252
rect 27804 19168 27856 19174
rect 27804 19110 27856 19116
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27356 17610 27384 18022
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 27264 16658 27292 16934
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27264 16046 27292 16594
rect 27632 16590 27660 17070
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27172 12406 27292 12434
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24122 9072 24178 9081
rect 24122 9007 24178 9016
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23952 7002 23980 7482
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23756 6928 23808 6934
rect 23756 6870 23808 6876
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 22756 5778 22784 6054
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 23400 5642 23428 6598
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5234 21404 5510
rect 22204 5234 22232 5578
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 17420 800 17448 2450
rect 17512 2446 17540 2790
rect 20088 2446 20116 2790
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 1170 20208 2450
rect 22020 2446 22048 2790
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 25516 2650 25544 5578
rect 27172 5370 27200 5578
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 25976 4554 26004 4966
rect 27264 4622 27292 12406
rect 27632 11200 27660 16186
rect 27724 12209 27752 18702
rect 27816 17082 27844 19110
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 28264 18352 28316 18358
rect 28368 18340 28396 19264
rect 28316 18312 28396 18340
rect 28264 18294 28316 18300
rect 28368 17746 28396 18312
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 28368 17270 28396 17682
rect 28356 17264 28408 17270
rect 28356 17206 28408 17212
rect 27816 17054 28396 17082
rect 28262 16688 28318 16697
rect 27804 16652 27856 16658
rect 28262 16623 28264 16632
rect 27804 16594 27856 16600
rect 28316 16623 28318 16632
rect 28264 16594 28316 16600
rect 27816 16250 27844 16594
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27804 16244 27856 16250
rect 27804 16186 27856 16192
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27710 12200 27766 12209
rect 27710 12135 27766 12144
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27632 11172 27752 11200
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 27632 7546 27660 11018
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27724 7426 27752 11172
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27804 9648 27856 9654
rect 27804 9590 27856 9596
rect 27816 9382 27844 9590
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27632 7398 27752 7426
rect 27632 5574 27660 7398
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 25964 4548 26016 4554
rect 25964 4490 26016 4496
rect 27264 3602 27292 4558
rect 27252 3596 27304 3602
rect 27252 3538 27304 3544
rect 27632 3534 27660 5510
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 28368 5302 28396 17054
rect 28460 16522 28488 17750
rect 28552 17105 28580 20862
rect 28828 20788 28856 21014
rect 28920 20942 28948 22086
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 29012 21622 29040 21830
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 28828 20760 28948 20788
rect 28816 20256 28868 20262
rect 28816 20198 28868 20204
rect 28630 19952 28686 19961
rect 28630 19887 28632 19896
rect 28684 19887 28686 19896
rect 28632 19858 28684 19864
rect 28828 19446 28856 20198
rect 28816 19440 28868 19446
rect 28816 19382 28868 19388
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28644 18358 28672 19110
rect 28632 18352 28684 18358
rect 28632 18294 28684 18300
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28828 17542 28856 17614
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 17338 28856 17478
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28538 17096 28594 17105
rect 28538 17031 28594 17040
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 28920 5778 28948 20760
rect 29000 20596 29052 20602
rect 29104 20584 29132 24006
rect 29184 22976 29236 22982
rect 29184 22918 29236 22924
rect 29196 22166 29224 22918
rect 29932 22710 29960 24142
rect 30116 23798 30144 26302
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26330 33838 27000
rect 33782 26302 34100 26330
rect 33782 26200 33838 26302
rect 30196 25220 30248 25226
rect 30196 25162 30248 25168
rect 30208 23866 30236 25162
rect 30380 25084 30432 25090
rect 30380 25026 30432 25032
rect 30392 24614 30420 25026
rect 30472 24676 30524 24682
rect 30472 24618 30524 24624
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 30196 23860 30248 23866
rect 30196 23802 30248 23808
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 30116 23202 30144 23734
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 30116 23174 30236 23202
rect 29920 22704 29972 22710
rect 29920 22646 29972 22652
rect 30104 22432 30156 22438
rect 30104 22374 30156 22380
rect 29184 22160 29236 22166
rect 29184 22102 29236 22108
rect 29828 22092 29880 22098
rect 29828 22034 29880 22040
rect 29840 21554 29868 22034
rect 30010 21992 30066 22001
rect 29920 21956 29972 21962
rect 30010 21927 30066 21936
rect 29920 21898 29972 21904
rect 29932 21865 29960 21898
rect 29918 21856 29974 21865
rect 29918 21791 29974 21800
rect 29828 21548 29880 21554
rect 29748 21508 29828 21536
rect 29184 21072 29236 21078
rect 29184 21014 29236 21020
rect 29052 20556 29132 20584
rect 29000 20538 29052 20544
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 29012 16658 29040 19858
rect 29196 19825 29224 21014
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29564 20346 29592 20878
rect 29748 20466 29776 21508
rect 29828 21490 29880 21496
rect 30024 21010 30052 21927
rect 30116 21486 30144 22374
rect 30208 21842 30236 23174
rect 30392 22778 30420 23666
rect 30484 22778 30512 24618
rect 30576 24206 30604 26200
rect 31116 25424 31168 25430
rect 31116 25366 31168 25372
rect 30656 24336 30708 24342
rect 30656 24278 30708 24284
rect 30564 24200 30616 24206
rect 30564 24142 30616 24148
rect 30668 23594 30696 24278
rect 31024 23860 31076 23866
rect 31024 23802 31076 23808
rect 30656 23588 30708 23594
rect 30656 23530 30708 23536
rect 30748 23588 30800 23594
rect 30748 23530 30800 23536
rect 30564 23520 30616 23526
rect 30616 23468 30696 23474
rect 30564 23462 30696 23468
rect 30576 23446 30696 23462
rect 30564 23316 30616 23322
rect 30564 23258 30616 23264
rect 30380 22772 30432 22778
rect 30380 22714 30432 22720
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30288 22160 30340 22166
rect 30340 22108 30420 22114
rect 30288 22102 30420 22108
rect 30300 22098 30420 22102
rect 30300 22092 30432 22098
rect 30300 22086 30380 22092
rect 30380 22034 30432 22040
rect 30472 22024 30524 22030
rect 30392 21972 30472 21978
rect 30392 21966 30524 21972
rect 30392 21950 30512 21966
rect 30208 21814 30328 21842
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 30300 21418 30328 21814
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29564 20330 29684 20346
rect 29564 20324 29696 20330
rect 29564 20318 29644 20324
rect 29182 19816 29238 19825
rect 29182 19751 29238 19760
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 29564 16017 29592 20318
rect 29644 20266 29696 20272
rect 29748 19718 29776 20402
rect 30208 20398 30236 21286
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29644 19372 29696 19378
rect 29748 19360 29776 19654
rect 29696 19332 29776 19360
rect 29644 19314 29696 19320
rect 29748 18902 29776 19332
rect 29736 18896 29788 18902
rect 29736 18838 29788 18844
rect 29748 18714 29776 18838
rect 29656 18686 29776 18714
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29656 18358 29684 18686
rect 29736 18624 29788 18630
rect 29736 18566 29788 18572
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 29656 17746 29684 18294
rect 29644 17740 29696 17746
rect 29644 17682 29696 17688
rect 29656 17338 29684 17682
rect 29644 17332 29696 17338
rect 29644 17274 29696 17280
rect 29550 16008 29606 16017
rect 29550 15943 29606 15952
rect 29748 15706 29776 18566
rect 29840 18086 29868 18702
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29932 15609 29960 19790
rect 30208 18834 30236 20198
rect 30300 19174 30328 20334
rect 30392 19854 30420 21950
rect 30576 21690 30604 23258
rect 30668 22273 30696 23446
rect 30760 23186 30788 23530
rect 30748 23180 30800 23186
rect 30748 23122 30800 23128
rect 30930 22672 30986 22681
rect 31036 22642 31064 23802
rect 31128 23526 31156 25366
rect 31116 23520 31168 23526
rect 31116 23462 31168 23468
rect 30930 22607 30932 22616
rect 30984 22607 30986 22616
rect 31024 22636 31076 22642
rect 30932 22578 30984 22584
rect 31024 22578 31076 22584
rect 30944 22438 30972 22578
rect 31220 22574 31248 26200
rect 31300 24744 31352 24750
rect 31300 24686 31352 24692
rect 31208 22568 31260 22574
rect 31208 22510 31260 22516
rect 30932 22432 30984 22438
rect 30932 22374 30984 22380
rect 30654 22264 30710 22273
rect 30654 22199 30710 22208
rect 30668 22094 30696 22199
rect 30944 22094 30972 22374
rect 30668 22066 30880 22094
rect 30944 22066 31064 22094
rect 30564 21684 30616 21690
rect 30564 21626 30616 21632
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30564 21004 30616 21010
rect 30564 20946 30616 20952
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 30392 19718 30420 19790
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30392 19514 30420 19654
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30116 18426 30144 18566
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30392 18034 30420 18090
rect 30300 18006 30420 18034
rect 30300 17746 30328 18006
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 17338 30236 17478
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30208 17066 30236 17274
rect 30300 17134 30328 17682
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30196 17060 30248 17066
rect 30196 17002 30248 17008
rect 30208 16794 30236 17002
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 29918 15600 29974 15609
rect 29918 15535 29974 15544
rect 30576 14958 30604 20946
rect 30668 20874 30696 21286
rect 30656 20868 30708 20874
rect 30656 20810 30708 20816
rect 30852 20602 30880 22066
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 30654 19408 30710 19417
rect 30654 19343 30656 19352
rect 30708 19343 30710 19352
rect 30656 19314 30708 19320
rect 30932 19304 30984 19310
rect 30932 19246 30984 19252
rect 30748 18964 30800 18970
rect 30748 18906 30800 18912
rect 30760 18426 30788 18906
rect 30944 18902 30972 19246
rect 30932 18896 30984 18902
rect 30932 18838 30984 18844
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30656 18352 30708 18358
rect 30656 18294 30708 18300
rect 30668 18057 30696 18294
rect 30654 18048 30710 18057
rect 30654 17983 30710 17992
rect 31036 17678 31064 22066
rect 31116 22092 31168 22098
rect 31116 22034 31168 22040
rect 31128 21865 31156 22034
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31114 21856 31170 21865
rect 31114 21791 31170 21800
rect 31114 21448 31170 21457
rect 31114 21383 31170 21392
rect 31128 20942 31156 21383
rect 31220 21010 31248 21898
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31220 18873 31248 20742
rect 31206 18864 31262 18873
rect 31206 18799 31262 18808
rect 31312 18358 31340 24686
rect 31668 24676 31720 24682
rect 31668 24618 31720 24624
rect 31680 24410 31708 24618
rect 31576 24404 31628 24410
rect 31576 24346 31628 24352
rect 31668 24404 31720 24410
rect 31668 24346 31720 24352
rect 31588 24290 31616 24346
rect 31588 24262 31708 24290
rect 31680 24138 31708 24262
rect 31864 24206 31892 26200
rect 32508 25378 32536 26200
rect 32312 25356 32364 25362
rect 32312 25298 32364 25304
rect 32416 25350 32536 25378
rect 31852 24200 31904 24206
rect 31852 24142 31904 24148
rect 31576 24132 31628 24138
rect 31576 24074 31628 24080
rect 31668 24132 31720 24138
rect 31668 24074 31720 24080
rect 31392 23724 31444 23730
rect 31392 23666 31444 23672
rect 31404 21418 31432 23666
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31496 22506 31524 22918
rect 31484 22500 31536 22506
rect 31484 22442 31536 22448
rect 31496 22166 31524 22442
rect 31484 22160 31536 22166
rect 31484 22102 31536 22108
rect 31588 21622 31616 24074
rect 31852 24064 31904 24070
rect 31852 24006 31904 24012
rect 31668 23588 31720 23594
rect 31760 23588 31812 23594
rect 31720 23548 31760 23576
rect 31668 23530 31720 23536
rect 31760 23530 31812 23536
rect 31668 22772 31720 22778
rect 31668 22714 31720 22720
rect 31680 22642 31708 22714
rect 31772 22710 31800 23530
rect 31864 23322 31892 24006
rect 32324 23798 32352 25298
rect 32312 23792 32364 23798
rect 32312 23734 32364 23740
rect 32128 23656 32180 23662
rect 32128 23598 32180 23604
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 31864 23118 31892 23258
rect 31852 23112 31904 23118
rect 31852 23054 31904 23060
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 31760 22704 31812 22710
rect 31760 22646 31812 22652
rect 31668 22636 31720 22642
rect 31668 22578 31720 22584
rect 31864 22234 31892 23054
rect 31944 22976 31996 22982
rect 31944 22918 31996 22924
rect 31852 22228 31904 22234
rect 31852 22170 31904 22176
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31392 21412 31444 21418
rect 31392 21354 31444 21360
rect 31680 21010 31708 21830
rect 31864 21350 31892 22170
rect 31956 21554 31984 22918
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 31852 21344 31904 21350
rect 31852 21286 31904 21292
rect 31668 21004 31720 21010
rect 31864 20992 31892 21286
rect 31956 21146 31984 21490
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31668 20946 31720 20952
rect 31772 20964 31892 20992
rect 31680 19854 31708 20946
rect 31772 20602 31800 20964
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 31772 20074 31800 20538
rect 31864 20369 31892 20810
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31850 20360 31906 20369
rect 31850 20295 31906 20304
rect 31772 20046 31892 20074
rect 31760 19984 31812 19990
rect 31760 19926 31812 19932
rect 31668 19848 31720 19854
rect 31668 19790 31720 19796
rect 31772 19009 31800 19926
rect 31864 19378 31892 20046
rect 31852 19372 31904 19378
rect 31852 19314 31904 19320
rect 31758 19000 31814 19009
rect 31758 18935 31814 18944
rect 31300 18352 31352 18358
rect 31300 18294 31352 18300
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 30932 17604 30984 17610
rect 30932 17546 30984 17552
rect 30944 17338 30972 17546
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 31036 17270 31064 17614
rect 31024 17264 31076 17270
rect 31024 17206 31076 17212
rect 31036 16697 31064 17206
rect 31022 16688 31078 16697
rect 31022 16623 31078 16632
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 31864 11354 31892 19314
rect 31956 15473 31984 20742
rect 32048 19922 32076 23054
rect 32036 19916 32088 19922
rect 32036 19858 32088 19864
rect 32140 19514 32168 23598
rect 32312 23316 32364 23322
rect 32312 23258 32364 23264
rect 32324 22794 32352 23258
rect 32416 22964 32444 25350
rect 32496 25288 32548 25294
rect 32496 25230 32548 25236
rect 32508 23322 32536 25230
rect 32864 25016 32916 25022
rect 32864 24958 32916 24964
rect 32680 24200 32732 24206
rect 32680 24142 32732 24148
rect 32588 23588 32640 23594
rect 32588 23530 32640 23536
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 32496 22976 32548 22982
rect 32416 22936 32496 22964
rect 32496 22918 32548 22924
rect 32324 22766 32536 22794
rect 32508 22642 32536 22766
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32232 21049 32260 22170
rect 32416 21894 32444 22578
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32508 22137 32536 22374
rect 32494 22128 32550 22137
rect 32494 22063 32550 22072
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32218 21040 32274 21049
rect 32218 20975 32274 20984
rect 32324 20505 32352 21490
rect 32310 20496 32366 20505
rect 32310 20431 32366 20440
rect 32128 19508 32180 19514
rect 32128 19450 32180 19456
rect 31942 15464 31998 15473
rect 31942 15399 31998 15408
rect 31852 11348 31904 11354
rect 31852 11290 31904 11296
rect 31864 11150 31892 11290
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31312 9654 31340 11018
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 28356 5296 28408 5302
rect 28356 5238 28408 5244
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27816 2650 27844 4626
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28736 2650 28764 5714
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 28828 4826 28856 5102
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 28920 3670 28948 5714
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 31588 2514 31616 9318
rect 32416 9178 32444 21830
rect 32496 21344 32548 21350
rect 32496 21286 32548 21292
rect 32508 13394 32536 21286
rect 32600 21146 32628 23530
rect 32692 22098 32720 24142
rect 32876 23798 32904 24958
rect 33152 24664 33180 26200
rect 33968 25764 34020 25770
rect 33968 25706 34020 25712
rect 33600 25560 33652 25566
rect 33600 25502 33652 25508
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33152 24636 33364 24664
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 33336 24206 33364 24636
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 32864 23792 32916 23798
rect 32864 23734 32916 23740
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33336 23202 33364 24142
rect 33416 24064 33468 24070
rect 33416 24006 33468 24012
rect 33428 23769 33456 24006
rect 33414 23760 33470 23769
rect 33414 23695 33470 23704
rect 33520 23322 33548 24822
rect 33612 23798 33640 25502
rect 33876 24336 33928 24342
rect 33876 24278 33928 24284
rect 33600 23792 33652 23798
rect 33600 23734 33652 23740
rect 33888 23526 33916 24278
rect 33876 23520 33928 23526
rect 33876 23462 33928 23468
rect 33980 23322 34008 25706
rect 34072 24342 34100 26302
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26330 37058 27000
rect 37002 26302 37228 26330
rect 37002 26200 37058 26302
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34164 24410 34192 24550
rect 34152 24404 34204 24410
rect 34152 24346 34204 24352
rect 34060 24336 34112 24342
rect 34060 24278 34112 24284
rect 34072 24206 34100 24278
rect 34060 24200 34112 24206
rect 34440 24188 34468 26200
rect 34888 25628 34940 25634
rect 34888 25570 34940 25576
rect 34520 24200 34572 24206
rect 34440 24160 34520 24188
rect 34060 24142 34112 24148
rect 34520 24142 34572 24148
rect 34900 23798 34928 25570
rect 34980 25492 35032 25498
rect 34980 25434 35032 25440
rect 34992 23798 35020 25434
rect 35084 24290 35112 26200
rect 35084 24262 35204 24290
rect 35070 24168 35126 24177
rect 35176 24138 35204 24262
rect 35624 24200 35676 24206
rect 35728 24188 35756 26200
rect 35898 24984 35954 24993
rect 35898 24919 35954 24928
rect 35912 24342 35940 24919
rect 35900 24336 35952 24342
rect 35900 24278 35952 24284
rect 35900 24200 35952 24206
rect 35728 24160 35900 24188
rect 35624 24142 35676 24148
rect 35900 24142 35952 24148
rect 35070 24103 35126 24112
rect 35164 24132 35216 24138
rect 35084 24070 35112 24103
rect 35164 24074 35216 24080
rect 35072 24064 35124 24070
rect 35072 24006 35124 24012
rect 35256 24064 35308 24070
rect 35256 24006 35308 24012
rect 34888 23792 34940 23798
rect 34888 23734 34940 23740
rect 34980 23792 35032 23798
rect 34980 23734 35032 23740
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 33508 23316 33560 23322
rect 33508 23258 33560 23264
rect 33968 23316 34020 23322
rect 33968 23258 34020 23264
rect 34428 23316 34480 23322
rect 34428 23258 34480 23264
rect 33598 23216 33654 23225
rect 33336 23174 33456 23202
rect 32864 23044 32916 23050
rect 32864 22986 32916 22992
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 32876 22234 32904 22986
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32864 22228 32916 22234
rect 32864 22170 32916 22176
rect 32680 22092 32732 22098
rect 32680 22034 32732 22040
rect 33336 22030 33364 22986
rect 33428 22506 33456 23174
rect 33598 23151 33654 23160
rect 33612 22642 33640 23151
rect 33874 22672 33930 22681
rect 33600 22636 33652 22642
rect 33874 22607 33876 22616
rect 33600 22578 33652 22584
rect 33928 22607 33930 22616
rect 33876 22578 33928 22584
rect 34440 22574 34468 23258
rect 34716 22778 34744 23666
rect 35072 23248 35124 23254
rect 35072 23190 35124 23196
rect 34980 23112 35032 23118
rect 34886 23080 34942 23089
rect 34980 23054 35032 23060
rect 34886 23015 34942 23024
rect 34900 22982 34928 23015
rect 34888 22976 34940 22982
rect 34888 22918 34940 22924
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34992 22642 35020 23054
rect 35084 22982 35112 23190
rect 35072 22976 35124 22982
rect 35072 22918 35124 22924
rect 35072 22772 35124 22778
rect 35072 22714 35124 22720
rect 34980 22636 35032 22642
rect 34980 22578 35032 22584
rect 34428 22568 34480 22574
rect 34428 22510 34480 22516
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 33416 22500 33468 22506
rect 33416 22442 33468 22448
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 32784 21350 32812 21966
rect 32772 21344 32824 21350
rect 32772 21286 32824 21292
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32784 21078 32812 21286
rect 32772 21072 32824 21078
rect 32772 21014 32824 21020
rect 32680 20936 32732 20942
rect 32680 20878 32732 20884
rect 32692 18193 32720 20878
rect 32678 18184 32734 18193
rect 32678 18119 32734 18128
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32876 8401 32904 21966
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 33336 15065 33364 21966
rect 34520 21412 34572 21418
rect 34520 21354 34572 21360
rect 34532 17678 34560 21354
rect 34624 18222 34652 22510
rect 34612 18216 34664 18222
rect 34612 18158 34664 18164
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34520 17264 34572 17270
rect 34520 17206 34572 17212
rect 34532 15638 34560 17206
rect 34520 15632 34572 15638
rect 34520 15574 34572 15580
rect 33322 15056 33378 15065
rect 33322 14991 33378 15000
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 35084 14074 35112 22714
rect 35268 21962 35296 24006
rect 35636 23254 35664 24142
rect 36268 24132 36320 24138
rect 36268 24074 36320 24080
rect 36280 23905 36308 24074
rect 36266 23896 36322 23905
rect 36266 23831 36322 23840
rect 36372 23730 36400 26200
rect 36636 24744 36688 24750
rect 36636 24686 36688 24692
rect 36648 24138 36676 24686
rect 36912 24336 36964 24342
rect 36912 24278 36964 24284
rect 36820 24200 36872 24206
rect 36820 24142 36872 24148
rect 36636 24132 36688 24138
rect 36636 24074 36688 24080
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 35624 23248 35676 23254
rect 35624 23190 35676 23196
rect 35716 23112 35768 23118
rect 35716 23054 35768 23060
rect 35728 22438 35756 23054
rect 36280 23050 36308 23666
rect 36268 23044 36320 23050
rect 36268 22986 36320 22992
rect 36176 22976 36228 22982
rect 36176 22918 36228 22924
rect 35716 22432 35768 22438
rect 35716 22374 35768 22380
rect 35256 21956 35308 21962
rect 35256 21898 35308 21904
rect 36188 21593 36216 22918
rect 36174 21584 36230 21593
rect 36174 21519 36230 21528
rect 36464 21010 36492 24006
rect 36542 23896 36598 23905
rect 36542 23831 36598 23840
rect 36556 23798 36584 23831
rect 36544 23792 36596 23798
rect 36544 23734 36596 23740
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36740 21690 36768 23462
rect 36832 23322 36860 24142
rect 36820 23316 36872 23322
rect 36820 23258 36872 23264
rect 36728 21684 36780 21690
rect 36728 21626 36780 21632
rect 36452 21004 36504 21010
rect 36452 20946 36504 20952
rect 36924 20466 36952 24278
rect 37200 24188 37228 26302
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38934 26330 38990 27000
rect 38290 26302 38516 26330
rect 38290 26200 38346 26302
rect 37280 24200 37332 24206
rect 37200 24160 37280 24188
rect 37280 24142 37332 24148
rect 37188 23588 37240 23594
rect 37188 23530 37240 23536
rect 36912 20460 36964 20466
rect 36912 20402 36964 20408
rect 37200 19718 37228 23530
rect 37292 23322 37320 24142
rect 37660 23730 37688 26200
rect 38488 24206 38516 26302
rect 38934 26302 39252 26330
rect 38934 26200 38990 26302
rect 39224 24206 39252 26302
rect 39578 26200 39634 27000
rect 40222 26330 40278 27000
rect 40222 26302 40356 26330
rect 40222 26200 40278 26302
rect 39304 24948 39356 24954
rect 39304 24890 39356 24896
rect 39316 24410 39344 24890
rect 39304 24404 39356 24410
rect 39304 24346 39356 24352
rect 39592 24274 39620 26200
rect 40130 24304 40186 24313
rect 39580 24268 39632 24274
rect 40130 24239 40132 24248
rect 39580 24210 39632 24216
rect 40184 24239 40186 24248
rect 40132 24210 40184 24216
rect 38476 24200 38528 24206
rect 38476 24142 38528 24148
rect 38660 24200 38712 24206
rect 38660 24142 38712 24148
rect 39212 24200 39264 24206
rect 39212 24142 39264 24148
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38488 23866 38516 24142
rect 38476 23860 38528 23866
rect 38476 23802 38528 23808
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 38672 23633 38700 24142
rect 39224 23866 39252 24142
rect 39592 23866 39620 24210
rect 40328 23866 40356 26302
rect 40866 26200 40922 27000
rect 41510 26200 41566 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26330 43498 27000
rect 43442 26302 43760 26330
rect 43442 26200 43498 26302
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 39580 23860 39632 23866
rect 39580 23802 39632 23808
rect 40316 23860 40368 23866
rect 40316 23802 40368 23808
rect 40880 23746 40908 26200
rect 41524 24206 41552 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 41512 24200 41564 24206
rect 41512 24142 41564 24148
rect 43260 24200 43312 24206
rect 43260 24142 43312 24148
rect 41524 23866 41552 24142
rect 42064 24064 42116 24070
rect 42064 24006 42116 24012
rect 42616 24064 42668 24070
rect 42616 24006 42668 24012
rect 41512 23860 41564 23866
rect 41512 23802 41564 23808
rect 40880 23730 41000 23746
rect 42076 23730 42104 24006
rect 40880 23724 41012 23730
rect 40880 23718 40960 23724
rect 40960 23666 41012 23672
rect 42064 23724 42116 23730
rect 42064 23666 42116 23672
rect 38658 23624 38714 23633
rect 38658 23559 38714 23568
rect 40776 23588 40828 23594
rect 40776 23530 40828 23536
rect 37740 23520 37792 23526
rect 37740 23462 37792 23468
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 37752 21418 37780 23462
rect 39948 22976 40000 22982
rect 39948 22918 40000 22924
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 39960 22710 39988 22918
rect 39948 22704 40000 22710
rect 39948 22646 40000 22652
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37740 21412 37792 21418
rect 37740 21354 37792 21360
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37188 19712 37240 19718
rect 37188 19654 37240 19660
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 40788 15366 40816 23530
rect 41420 23520 41472 23526
rect 41420 23462 41472 23468
rect 41432 18154 41460 23462
rect 42628 23118 42656 24006
rect 43272 23866 43300 24142
rect 43260 23860 43312 23866
rect 43260 23802 43312 23808
rect 43732 23730 43760 26302
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26330 45430 27000
rect 45374 26302 45508 26330
rect 45374 26200 45430 26302
rect 44100 23746 44128 26200
rect 44744 24410 44772 26200
rect 44732 24404 44784 24410
rect 44732 24346 44784 24352
rect 44744 24206 44772 24346
rect 45480 24290 45508 26302
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26330 48006 27000
rect 47872 26302 48006 26330
rect 45480 24262 45600 24290
rect 45572 24206 45600 24262
rect 46032 24206 46060 26200
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 46020 24200 46072 24206
rect 46020 24142 46072 24148
rect 45376 24064 45428 24070
rect 45376 24006 45428 24012
rect 44100 23730 44220 23746
rect 43720 23724 43772 23730
rect 44100 23724 44232 23730
rect 44100 23718 44180 23724
rect 43720 23666 43772 23672
rect 44180 23666 44232 23672
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 43732 23322 43760 23666
rect 44640 23520 44692 23526
rect 44640 23462 44692 23468
rect 43720 23316 43772 23322
rect 43720 23258 43772 23264
rect 42616 23112 42668 23118
rect 42616 23054 42668 23060
rect 44548 22976 44600 22982
rect 44548 22918 44600 22924
rect 44560 22778 44588 22918
rect 44548 22772 44600 22778
rect 44548 22714 44600 22720
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 41420 18148 41472 18154
rect 41420 18090 41472 18096
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 44652 17649 44680 23462
rect 45388 18737 45416 24006
rect 45572 23866 45600 24142
rect 45560 23860 45612 23866
rect 45560 23802 45612 23808
rect 46676 23730 46704 26200
rect 47320 24206 47348 26200
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 46848 24064 46900 24070
rect 46848 24006 46900 24012
rect 47032 24064 47084 24070
rect 47032 24006 47084 24012
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 46860 18834 46888 24006
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 46952 19990 46980 23462
rect 46940 19984 46992 19990
rect 46940 19926 46992 19932
rect 46848 18828 46900 18834
rect 46848 18770 46900 18776
rect 45374 18728 45430 18737
rect 45374 18663 45430 18672
rect 44638 17640 44694 17649
rect 44638 17575 44694 17584
rect 47044 16998 47072 24006
rect 47320 23866 47348 24142
rect 47872 23866 47900 26302
rect 47950 26200 48006 26302
rect 48594 26200 48650 27000
rect 48318 24848 48374 24857
rect 48318 24783 48374 24792
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 47860 23860 47912 23866
rect 47860 23802 47912 23808
rect 48332 23730 48360 24783
rect 48608 24206 48636 26200
rect 48596 24200 48648 24206
rect 48596 24142 48648 24148
rect 48320 23724 48372 23730
rect 48320 23666 48372 23672
rect 48504 23520 48556 23526
rect 48504 23462 48556 23468
rect 47216 22976 47268 22982
rect 47216 22918 47268 22924
rect 47228 17066 47256 22918
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48320 22432 48372 22438
rect 48320 22374 48372 22380
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 47872 21350 47900 21490
rect 47860 21344 47912 21350
rect 47860 21286 47912 21292
rect 47216 17060 47268 17066
rect 47216 17002 47268 17008
rect 47032 16992 47084 16998
rect 47032 16934 47084 16940
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 40776 15360 40828 15366
rect 40776 15302 40828 15308
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 35072 14068 35124 14074
rect 35072 14010 35124 14016
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 47872 11082 47900 21286
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48332 17270 48360 22374
rect 48516 18970 48544 23462
rect 48608 22778 48636 24142
rect 48688 24064 48740 24070
rect 48688 24006 48740 24012
rect 48700 23118 48728 24006
rect 49238 23896 49294 23905
rect 49238 23831 49294 23840
rect 48688 23112 48740 23118
rect 48688 23054 48740 23060
rect 49056 23112 49108 23118
rect 49056 23054 49108 23060
rect 49068 22953 49096 23054
rect 49054 22944 49110 22953
rect 49054 22879 49110 22888
rect 48596 22772 48648 22778
rect 48596 22714 48648 22720
rect 49252 22642 49280 23831
rect 49240 22636 49292 22642
rect 49240 22578 49292 22584
rect 49056 22024 49108 22030
rect 49054 21992 49056 22001
rect 49108 21992 49110 22001
rect 49054 21927 49110 21936
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21049 49188 21422
rect 49146 21040 49202 21049
rect 49146 20975 49202 20984
rect 49252 20058 49280 21830
rect 49240 20052 49292 20058
rect 49240 19994 49292 20000
rect 48504 18964 48556 18970
rect 48504 18906 48556 18912
rect 48320 17264 48372 17270
rect 48320 17206 48372 17212
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47860 11076 47912 11082
rect 47860 11018 47912 11024
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 32862 8392 32918 8401
rect 32862 8327 32918 8336
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 41420 5160 41472 5166
rect 41420 5102 41472 5108
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33520 2650 33548 5034
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 31576 2508 31628 2514
rect 31576 2450 31628 2456
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 20088 1142 20208 1170
rect 20088 800 20116 1142
rect 22756 800 22784 2450
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 25424 800 25452 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28092 870 28212 898
rect 28092 800 28120 870
rect 1398 0 1454 800
rect 4066 0 4122 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 17406 0 17462 800
rect 20074 0 20130 800
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 28078 0 28134 800
rect 28184 762 28212 870
rect 28368 762 28396 2382
rect 30760 800 30788 2382
rect 33428 800 33456 2382
rect 36096 800 36124 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38764 800 38792 3402
rect 41432 800 41460 5102
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 44088 3664 44140 3670
rect 44088 3606 44140 3612
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 44100 800 44128 3606
rect 46756 3596 46808 3602
rect 46756 3538 46808 3544
rect 46768 800 46796 3538
rect 49424 3528 49476 3534
rect 49424 3470 49476 3476
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49436 800 49464 3470
rect 28184 734 28396 762
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< via2 >>
rect 938 17040 994 17096
rect 938 12180 940 12200
rect 940 12180 992 12200
rect 992 12180 994 12200
rect 938 12144 994 12180
rect 1122 16632 1178 16688
rect 1490 23160 1546 23216
rect 1306 20712 1362 20768
rect 1490 19352 1546 19408
rect 1398 17856 1454 17912
rect 1214 16224 1270 16280
rect 1122 15816 1178 15872
rect 1490 16632 1546 16688
rect 1122 15000 1178 15056
rect 1306 15408 1362 15464
rect 1306 14592 1362 14648
rect 1306 14184 1362 14240
rect 1214 13368 1270 13424
rect 1306 10920 1362 10976
rect 2134 23432 2190 23488
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2778 24404 2834 24440
rect 2778 24384 2780 24404
rect 2780 24384 2832 24404
rect 2832 24384 2834 24404
rect 1766 19760 1822 19816
rect 2042 17448 2098 17504
rect 1858 13932 1914 13968
rect 1858 13912 1860 13932
rect 1860 13912 1912 13932
rect 1912 13912 1914 13932
rect 2042 13776 2098 13832
rect 1950 13368 2006 13424
rect 1766 11892 1822 11928
rect 1766 11872 1768 11892
rect 1768 11872 1820 11892
rect 1820 11872 1822 11892
rect 1674 11600 1730 11656
rect 1582 9696 1638 9752
rect 1306 7656 1362 7712
rect 1766 8880 1822 8936
rect 1306 6432 1362 6488
rect 1306 6024 1362 6080
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 1306 5228 1362 5264
rect 1306 5208 1308 5228
rect 1308 5208 1360 5228
rect 1360 5208 1362 5228
rect 1306 4800 1362 4856
rect 1766 4392 1822 4448
rect 1306 4020 1308 4040
rect 1308 4020 1360 4040
rect 1360 4020 1362 4040
rect 1306 3984 1362 4020
rect 1214 3576 1270 3632
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2686 21528 2742 21584
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3238 21528 3294 21584
rect 3606 25608 3662 25664
rect 2870 21392 2926 21448
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2778 19896 2834 19952
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2778 19624 2834 19680
rect 2686 19080 2742 19136
rect 3330 19624 3386 19680
rect 2962 19488 3018 19544
rect 3330 19080 3386 19136
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18672 2926 18728
rect 2778 18264 2834 18320
rect 2778 18128 2834 18184
rect 3330 18128 3386 18184
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3422 17876 3478 17912
rect 3422 17856 3424 17876
rect 3424 17856 3476 17876
rect 3476 17856 3478 17876
rect 4066 25220 4122 25256
rect 4066 25200 4068 25220
rect 4068 25200 4120 25220
rect 4120 25200 4122 25220
rect 4066 24792 4122 24848
rect 3882 23976 3938 24032
rect 4802 24792 4858 24848
rect 4066 23604 4068 23624
rect 4068 23604 4120 23624
rect 4120 23604 4122 23624
rect 4066 23568 4122 23604
rect 3606 22752 3662 22808
rect 3790 22344 3846 22400
rect 4250 23160 4306 23216
rect 4158 22616 4214 22672
rect 4066 22480 4122 22536
rect 3606 21664 3662 21720
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2778 16496 2834 16552
rect 2594 11056 2650 11112
rect 2778 10512 2834 10568
rect 1306 3168 1362 3224
rect 1306 2760 1362 2816
rect 1214 2352 1270 2408
rect 1306 1944 1362 2000
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 3422 16652 3478 16688
rect 3422 16632 3424 16652
rect 3424 16632 3476 16652
rect 3476 16632 3478 16652
rect 3330 13640 3386 13696
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2870 10104 2926 10160
rect 2778 9288 2834 9344
rect 3238 9596 3240 9616
rect 3240 9596 3292 9616
rect 3292 9596 3294 9616
rect 3238 9560 3294 9596
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2870 8472 2926 8528
rect 3974 20712 4030 20768
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 3698 16768 3754 16824
rect 3790 16224 3846 16280
rect 3514 12144 3570 12200
rect 3514 11600 3570 11656
rect 3882 13268 3884 13288
rect 3884 13268 3936 13288
rect 3936 13268 3938 13288
rect 3882 13232 3938 13268
rect 3882 12960 3938 13016
rect 3790 11464 3846 11520
rect 3698 11192 3754 11248
rect 3422 10004 3424 10024
rect 3424 10004 3476 10024
rect 3476 10004 3478 10024
rect 3422 9968 3478 10004
rect 3606 9444 3662 9480
rect 3606 9424 3608 9444
rect 3608 9424 3660 9444
rect 3660 9424 3662 9444
rect 3790 11056 3846 11112
rect 3790 9424 3846 9480
rect 2778 8064 2834 8120
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3330 7812 3386 7848
rect 3330 7792 3332 7812
rect 3332 7792 3384 7812
rect 3384 7792 3386 7812
rect 2870 7248 2926 7304
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 4250 21936 4306 21992
rect 4250 21004 4306 21040
rect 4250 20984 4252 21004
rect 4252 20984 4304 21004
rect 4304 20984 4306 21004
rect 4066 15444 4068 15464
rect 4068 15444 4120 15464
rect 4120 15444 4122 15464
rect 4066 15408 4122 15444
rect 4250 17448 4306 17504
rect 4434 19896 4490 19952
rect 4526 18808 4582 18864
rect 4710 18572 4712 18592
rect 4712 18572 4764 18592
rect 4764 18572 4766 18592
rect 4710 18536 4766 18572
rect 4802 17584 4858 17640
rect 4066 12688 4122 12744
rect 4526 14048 4582 14104
rect 4526 13640 4582 13696
rect 4158 12552 4214 12608
rect 4158 12280 4214 12336
rect 4434 12552 4490 12608
rect 4342 10376 4398 10432
rect 4066 9968 4122 10024
rect 3882 7792 3938 7848
rect 3330 6860 3386 6896
rect 3330 6840 3332 6860
rect 3332 6840 3384 6860
rect 3384 6840 3386 6860
rect 4710 16904 4766 16960
rect 5078 17040 5134 17096
rect 5998 22072 6054 22128
rect 5630 21392 5686 21448
rect 5262 17992 5318 18048
rect 5170 14456 5226 14512
rect 5630 20868 5686 20904
rect 5630 20848 5632 20868
rect 5632 20848 5684 20868
rect 5684 20848 5686 20868
rect 5630 20032 5686 20088
rect 5630 17992 5686 18048
rect 5446 14592 5502 14648
rect 6090 18672 6146 18728
rect 6182 18536 6238 18592
rect 6090 17992 6146 18048
rect 5722 14048 5778 14104
rect 6458 20712 6514 20768
rect 6550 20032 6606 20088
rect 6550 19252 6552 19272
rect 6552 19252 6604 19272
rect 6604 19252 6606 19272
rect 6550 19216 6606 19252
rect 6458 16496 6514 16552
rect 5446 11056 5502 11112
rect 5354 10920 5410 10976
rect 5630 10784 5686 10840
rect 7194 22616 7250 22672
rect 7010 21120 7066 21176
rect 7010 20848 7066 20904
rect 7010 19216 7066 19272
rect 6642 14728 6698 14784
rect 5906 11056 5962 11112
rect 5630 9832 5686 9888
rect 5538 9560 5594 9616
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 6182 11192 6238 11248
rect 6550 13640 6606 13696
rect 6458 11736 6514 11792
rect 6458 8628 6514 8664
rect 6458 8608 6460 8628
rect 6460 8608 6512 8628
rect 6512 8608 6514 8628
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2870 1536 2926 1592
rect 7286 21664 7342 21720
rect 7470 23432 7526 23488
rect 7562 21392 7618 21448
rect 7194 17856 7250 17912
rect 6734 12280 6790 12336
rect 7470 19372 7526 19408
rect 7470 19352 7472 19372
rect 7472 19352 7524 19372
rect 7524 19352 7526 19372
rect 7562 18264 7618 18320
rect 7470 17720 7526 17776
rect 7470 17448 7526 17504
rect 7286 16088 7342 16144
rect 7102 15408 7158 15464
rect 7378 15444 7380 15464
rect 7380 15444 7432 15464
rect 7432 15444 7434 15464
rect 7378 15408 7434 15444
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 8298 23704 8354 23760
rect 7930 23024 7986 23080
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8206 20868 8262 20904
rect 8206 20848 8208 20868
rect 8208 20848 8260 20868
rect 8260 20848 8262 20868
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8758 21972 8760 21992
rect 8760 21972 8812 21992
rect 8812 21972 8814 21992
rect 8758 21936 8814 21972
rect 8942 21392 8998 21448
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8114 17176 8170 17232
rect 8206 17076 8208 17096
rect 8208 17076 8260 17096
rect 8260 17076 8262 17096
rect 8206 17040 8262 17076
rect 8206 16652 8262 16688
rect 8206 16632 8208 16652
rect 8208 16632 8260 16652
rect 8260 16632 8262 16652
rect 8206 16496 8262 16552
rect 7562 16088 7618 16144
rect 7562 15988 7564 16008
rect 7564 15988 7616 16008
rect 7616 15988 7618 16008
rect 7562 15952 7618 15988
rect 7654 15680 7710 15736
rect 7470 12824 7526 12880
rect 7010 10648 7066 10704
rect 6642 8880 6698 8936
rect 6918 10104 6974 10160
rect 7286 11328 7342 11384
rect 7654 14320 7710 14376
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8114 15952 8170 16008
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7838 14900 7840 14920
rect 7840 14900 7892 14920
rect 7892 14900 7894 14920
rect 7838 14864 7894 14900
rect 7194 9172 7250 9208
rect 7194 9152 7196 9172
rect 7196 9152 7248 9172
rect 7248 9152 7250 9172
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 8574 18672 8630 18728
rect 9218 24112 9274 24168
rect 9402 22072 9458 22128
rect 9678 21836 9680 21856
rect 9680 21836 9732 21856
rect 9732 21836 9734 21856
rect 9678 21800 9734 21836
rect 9402 20748 9404 20768
rect 9404 20748 9456 20768
rect 9456 20748 9458 20768
rect 9402 20712 9458 20748
rect 9310 19760 9366 19816
rect 9218 19352 9274 19408
rect 9126 18672 9182 18728
rect 10138 19252 10140 19272
rect 10140 19252 10192 19272
rect 10192 19252 10194 19272
rect 10138 19216 10194 19252
rect 9678 18264 9734 18320
rect 9494 17992 9550 18048
rect 9310 17312 9366 17368
rect 9494 17332 9550 17368
rect 9494 17312 9496 17332
rect 9496 17312 9548 17332
rect 9548 17312 9550 17332
rect 9218 16788 9274 16824
rect 9218 16768 9220 16788
rect 9220 16768 9272 16788
rect 9272 16768 9274 16788
rect 8574 14456 8630 14512
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7746 9016 7802 9072
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 8758 12860 8760 12880
rect 8760 12860 8812 12880
rect 8812 12860 8814 12880
rect 8758 12824 8814 12860
rect 9218 15428 9274 15464
rect 9218 15408 9220 15428
rect 9220 15408 9272 15428
rect 9272 15408 9274 15428
rect 9494 16088 9550 16144
rect 9678 16496 9734 16552
rect 9402 15000 9458 15056
rect 9678 15000 9734 15056
rect 9494 14728 9550 14784
rect 9402 13268 9404 13288
rect 9404 13268 9456 13288
rect 9456 13268 9458 13288
rect 9402 13232 9458 13268
rect 9310 11772 9312 11792
rect 9312 11772 9364 11792
rect 9364 11772 9366 11792
rect 9310 11736 9366 11772
rect 9770 14320 9826 14376
rect 9770 13776 9826 13832
rect 9310 8200 9366 8256
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 10046 13776 10102 13832
rect 9954 12552 10010 12608
rect 11058 24248 11114 24304
rect 11150 22480 11206 22536
rect 10966 21800 11022 21856
rect 10506 21528 10562 21584
rect 10874 17720 10930 17776
rect 10782 17448 10838 17504
rect 10414 17312 10470 17368
rect 10598 16224 10654 16280
rect 10966 15972 11022 16008
rect 10966 15952 10968 15972
rect 10968 15952 11020 15972
rect 11020 15952 11022 15972
rect 10506 14320 10562 14376
rect 10966 15272 11022 15328
rect 10966 15036 10968 15056
rect 10968 15036 11020 15056
rect 11020 15036 11022 15056
rect 10966 15000 11022 15036
rect 10966 14900 10968 14920
rect 10968 14900 11020 14920
rect 11020 14900 11022 14920
rect 10966 14864 11022 14900
rect 11242 19216 11298 19272
rect 11426 19896 11482 19952
rect 11426 19388 11428 19408
rect 11428 19388 11480 19408
rect 11480 19388 11482 19408
rect 11426 19352 11482 19388
rect 11610 21120 11666 21176
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 13266 23568 13322 23624
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12346 21140 12402 21176
rect 12346 21120 12348 21140
rect 12348 21120 12400 21140
rect 12400 21120 12402 21140
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 13634 23704 13690 23760
rect 13542 23432 13598 23488
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 11794 20440 11850 20496
rect 11978 20304 12034 20360
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 14186 23296 14242 23352
rect 14462 23296 14518 23352
rect 14370 23044 14426 23080
rect 14370 23024 14372 23044
rect 14372 23024 14424 23044
rect 14424 23024 14426 23044
rect 14646 21956 14702 21992
rect 14646 21936 14648 21956
rect 14648 21936 14700 21956
rect 14700 21936 14702 21956
rect 13910 21120 13966 21176
rect 13910 20748 13912 20768
rect 13912 20748 13964 20768
rect 13964 20748 13966 20768
rect 13910 20712 13966 20748
rect 13542 20168 13598 20224
rect 12990 19760 13046 19816
rect 11702 17584 11758 17640
rect 11150 15136 11206 15192
rect 11058 14592 11114 14648
rect 11058 14456 11114 14512
rect 10966 14320 11022 14376
rect 10782 13776 10838 13832
rect 10690 12960 10746 13016
rect 10690 12844 10746 12880
rect 10690 12824 10692 12844
rect 10692 12824 10744 12844
rect 10744 12824 10746 12844
rect 9862 8356 9918 8392
rect 9862 8336 9864 8356
rect 9864 8336 9916 8356
rect 9916 8336 9918 8356
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 11334 15816 11390 15872
rect 11702 16768 11758 16824
rect 11334 13640 11390 13696
rect 11150 11600 11206 11656
rect 12070 19216 12126 19272
rect 12162 18148 12218 18184
rect 12162 18128 12164 18148
rect 12164 18128 12216 18148
rect 12216 18128 12218 18148
rect 12070 15580 12072 15600
rect 12072 15580 12124 15600
rect 12124 15580 12126 15600
rect 12070 15544 12126 15580
rect 11886 15136 11942 15192
rect 11978 15020 12034 15056
rect 11978 15000 11980 15020
rect 11980 15000 12032 15020
rect 12032 15000 12034 15020
rect 11518 10412 11520 10432
rect 11520 10412 11572 10432
rect 11572 10412 11574 10432
rect 11518 10376 11574 10412
rect 11518 9832 11574 9888
rect 12070 14864 12126 14920
rect 11886 10376 11942 10432
rect 12714 19080 12770 19136
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13266 17756 13268 17776
rect 13268 17756 13320 17776
rect 13320 17756 13322 17776
rect 13266 17720 13322 17756
rect 12622 15680 12678 15736
rect 12806 16904 12862 16960
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13174 16396 13176 16416
rect 13176 16396 13228 16416
rect 13228 16396 13230 16416
rect 13174 16360 13230 16396
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13910 20304 13966 20360
rect 14186 17856 14242 17912
rect 13910 15816 13966 15872
rect 13726 15680 13782 15736
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13542 14864 13598 14920
rect 13174 12724 13176 12744
rect 13176 12724 13228 12744
rect 13228 12724 13230 12744
rect 13174 12688 13230 12724
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13266 12008 13322 12064
rect 13174 11872 13230 11928
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 14186 16632 14242 16688
rect 15014 22344 15070 22400
rect 15566 21412 15622 21448
rect 15566 21392 15568 21412
rect 15568 21392 15620 21412
rect 15620 21392 15622 21412
rect 14462 18808 14518 18864
rect 14554 16668 14556 16688
rect 14556 16668 14608 16688
rect 14608 16668 14610 16688
rect 14554 16632 14610 16668
rect 14370 11892 14426 11928
rect 14370 11872 14372 11892
rect 14372 11872 14424 11892
rect 14424 11872 14426 11892
rect 14830 18400 14886 18456
rect 15014 19216 15070 19272
rect 15014 18264 15070 18320
rect 15382 17992 15438 18048
rect 15750 21664 15806 21720
rect 15750 20848 15806 20904
rect 15474 15308 15476 15328
rect 15476 15308 15528 15328
rect 15528 15308 15530 15328
rect 15474 15272 15530 15308
rect 16302 24656 16358 24712
rect 15934 21664 15990 21720
rect 15934 21564 15936 21584
rect 15936 21564 15988 21584
rect 15988 21564 15990 21584
rect 15934 21528 15990 21564
rect 16762 21936 16818 21992
rect 16026 19624 16082 19680
rect 15842 18672 15898 18728
rect 15658 14456 15714 14512
rect 16578 20032 16634 20088
rect 16302 19080 16358 19136
rect 16486 18028 16488 18048
rect 16488 18028 16540 18048
rect 16540 18028 16542 18048
rect 16486 17992 16542 18028
rect 15658 14320 15714 14376
rect 15198 12280 15254 12336
rect 14278 11736 14334 11792
rect 13726 10240 13782 10296
rect 14646 9968 14702 10024
rect 13726 9424 13782 9480
rect 15658 9832 15714 9888
rect 16578 16360 16634 16416
rect 16946 21800 17002 21856
rect 17590 24248 17646 24304
rect 17314 20848 17370 20904
rect 17222 20576 17278 20632
rect 17222 20304 17278 20360
rect 16854 19080 16910 19136
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 18970 24268 19026 24304
rect 18970 24248 18972 24268
rect 18972 24248 19024 24268
rect 19024 24248 19026 24268
rect 17958 23160 18014 23216
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17774 22616 17830 22672
rect 17774 22480 17830 22536
rect 17774 21800 17830 21856
rect 17774 20596 17830 20632
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18602 21120 18658 21176
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17774 20576 17776 20596
rect 17776 20576 17828 20596
rect 17828 20576 17830 20596
rect 18510 20168 18566 20224
rect 17406 19488 17462 19544
rect 17222 19216 17278 19272
rect 16762 17312 16818 17368
rect 16762 15136 16818 15192
rect 17682 19660 17684 19680
rect 17684 19660 17736 19680
rect 17736 19660 17738 19680
rect 17498 19216 17554 19272
rect 17130 17720 17186 17776
rect 16946 17584 17002 17640
rect 16946 16904 17002 16960
rect 17130 16244 17186 16280
rect 17130 16224 17132 16244
rect 17132 16224 17184 16244
rect 17184 16224 17186 16244
rect 17682 19624 17738 19660
rect 17682 19488 17738 19544
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17682 19080 17738 19136
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17774 18400 17830 18456
rect 17130 14864 17186 14920
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18510 19488 18566 19544
rect 18510 18808 18566 18864
rect 18510 17176 18566 17232
rect 18694 18572 18696 18592
rect 18696 18572 18748 18592
rect 18748 18572 18750 18592
rect 18694 18536 18750 18572
rect 18970 17992 19026 18048
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 16578 12688 16634 12744
rect 16210 12044 16212 12064
rect 16212 12044 16264 12064
rect 16264 12044 16266 12064
rect 16210 12008 16266 12044
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17406 11756 17462 11792
rect 17406 11736 17408 11756
rect 17408 11736 17460 11756
rect 17460 11736 17462 11756
rect 18602 17040 18658 17096
rect 18786 16768 18842 16824
rect 18602 15136 18658 15192
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 19798 23568 19854 23624
rect 19430 23196 19432 23216
rect 19432 23196 19484 23216
rect 19484 23196 19486 23216
rect 19430 23160 19486 23196
rect 19614 22752 19670 22808
rect 19338 16496 19394 16552
rect 19338 14864 19394 14920
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 19706 20712 19762 20768
rect 19798 20032 19854 20088
rect 19798 17448 19854 17504
rect 20166 23840 20222 23896
rect 20810 24268 20866 24304
rect 21178 24792 21234 24848
rect 20810 24248 20812 24268
rect 20812 24248 20864 24268
rect 20864 24248 20866 24268
rect 21638 24384 21694 24440
rect 20074 17856 20130 17912
rect 19890 16088 19946 16144
rect 20350 16940 20352 16960
rect 20352 16940 20404 16960
rect 20404 16940 20406 16960
rect 20350 16904 20406 16940
rect 19522 13912 19578 13968
rect 19430 13368 19486 13424
rect 20166 14900 20168 14920
rect 20168 14900 20220 14920
rect 20220 14900 20222 14920
rect 20166 14864 20222 14900
rect 20350 15136 20406 15192
rect 21362 19488 21418 19544
rect 20994 17584 21050 17640
rect 20902 15680 20958 15736
rect 20258 12280 20314 12336
rect 21270 15852 21272 15872
rect 21272 15852 21324 15872
rect 21324 15852 21326 15872
rect 21270 15816 21326 15852
rect 21454 18420 21510 18456
rect 21454 18400 21456 18420
rect 21456 18400 21508 18420
rect 21508 18400 21510 18420
rect 21914 23432 21970 23488
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22282 23840 22338 23896
rect 22282 23568 22338 23624
rect 21822 22344 21878 22400
rect 22190 23432 22246 23488
rect 22742 23296 22798 23352
rect 22742 22888 22798 22944
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23938 22616 23994 22672
rect 23754 22208 23810 22264
rect 23294 21836 23296 21856
rect 23296 21836 23348 21856
rect 23348 21836 23350 21856
rect 23294 21800 23350 21836
rect 21822 17176 21878 17232
rect 21914 17076 21916 17096
rect 21916 17076 21968 17096
rect 21968 17076 21970 17096
rect 21914 17040 21970 17076
rect 21362 14320 21418 14376
rect 20626 11192 20682 11248
rect 21914 16768 21970 16824
rect 21914 16360 21970 16416
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23662 20576 23718 20632
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22374 13932 22430 13968
rect 22374 13912 22376 13932
rect 22376 13912 22428 13932
rect 22428 13912 22430 13932
rect 22282 12824 22338 12880
rect 22650 16768 22706 16824
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23386 18672 23442 18728
rect 23386 17992 23442 18048
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23754 18400 23810 18456
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22650 13912 22706 13968
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23662 17448 23718 17504
rect 23846 17176 23902 17232
rect 25410 23432 25466 23488
rect 24766 22888 24822 22944
rect 24950 22752 25006 22808
rect 24214 18536 24270 18592
rect 24306 17720 24362 17776
rect 23846 16632 23902 16688
rect 23846 13948 23848 13968
rect 23848 13948 23900 13968
rect 23900 13948 23902 13968
rect 23846 13912 23902 13948
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 24950 18400 25006 18456
rect 25134 18264 25190 18320
rect 26790 23468 26792 23488
rect 26792 23468 26844 23488
rect 26844 23468 26846 23488
rect 26790 23432 26846 23468
rect 26514 22208 26570 22264
rect 25410 20712 25466 20768
rect 27158 24656 27214 24712
rect 26238 21256 26294 21312
rect 26606 20596 26662 20632
rect 26606 20576 26608 20596
rect 26608 20576 26660 20596
rect 26660 20576 26662 20596
rect 27434 22636 27490 22672
rect 27434 22616 27436 22636
rect 27436 22616 27488 22636
rect 27488 22616 27490 22636
rect 27066 22208 27122 22264
rect 25686 17584 25742 17640
rect 25134 14864 25190 14920
rect 25594 15136 25650 15192
rect 26146 13232 26202 13288
rect 27526 22208 27582 22264
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 28722 21256 28778 21312
rect 28446 20712 28502 20768
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27434 19252 27436 19272
rect 27436 19252 27488 19272
rect 27488 19252 27490 19272
rect 27434 19216 27490 19252
rect 24122 9016 24178 9072
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 28262 16652 28318 16688
rect 28262 16632 28264 16652
rect 28264 16632 28316 16652
rect 28316 16632 28318 16652
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27710 12144 27766 12200
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 28630 19916 28686 19952
rect 28630 19896 28632 19916
rect 28632 19896 28684 19916
rect 28684 19896 28686 19916
rect 28538 17040 28594 17096
rect 30010 21936 30066 21992
rect 29918 21800 29974 21856
rect 29182 19760 29238 19816
rect 29550 15952 29606 16008
rect 30930 22636 30986 22672
rect 30930 22616 30932 22636
rect 30932 22616 30984 22636
rect 30984 22616 30986 22636
rect 30654 22208 30710 22264
rect 29918 15544 29974 15600
rect 30654 19372 30710 19408
rect 30654 19352 30656 19372
rect 30656 19352 30708 19372
rect 30708 19352 30710 19372
rect 30654 17992 30710 18048
rect 31114 21800 31170 21856
rect 31114 21392 31170 21448
rect 31206 18808 31262 18864
rect 31850 20304 31906 20360
rect 31758 18944 31814 19000
rect 31022 16632 31078 16688
rect 32494 22072 32550 22128
rect 32218 20984 32274 21040
rect 32310 20440 32366 20496
rect 31942 15408 31998 15464
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33414 23704 33470 23760
rect 35070 24112 35126 24168
rect 35898 24928 35954 24984
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 33598 23160 33654 23216
rect 33874 22636 33930 22672
rect 33874 22616 33876 22636
rect 33876 22616 33928 22636
rect 33928 22616 33930 22636
rect 34886 23024 34942 23080
rect 32678 18128 32734 18184
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 33322 15000 33378 15056
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 36266 23840 36322 23896
rect 36174 21528 36230 21584
rect 36542 23840 36598 23896
rect 40130 24268 40186 24304
rect 40130 24248 40132 24268
rect 40132 24248 40184 24268
rect 40184 24248 40186 24268
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 38658 23568 38714 23624
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 45374 18672 45430 18728
rect 44638 17584 44694 17640
rect 48318 24792 48374 24848
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49238 23840 49294 23896
rect 49054 22888 49110 22944
rect 49054 21972 49056 21992
rect 49056 21972 49108 21992
rect 49108 21972 49110 21992
rect 49054 21936 49110 21972
rect 49146 20984 49202 21040
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 32862 8336 32918 8392
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3601 25666 3667 25669
rect 0 25664 3667 25666
rect 0 25608 3606 25664
rect 3662 25608 3667 25664
rect 0 25606 3667 25608
rect 0 25576 800 25606
rect 3601 25603 3667 25606
rect 0 25258 800 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 800 25198
rect 4061 25195 4127 25198
rect 11646 24924 11652 24988
rect 11716 24986 11722 24988
rect 35893 24986 35959 24989
rect 11716 24984 35959 24986
rect 11716 24928 35898 24984
rect 35954 24928 35959 24984
rect 11716 24926 35959 24928
rect 11716 24924 11722 24926
rect 35893 24923 35959 24926
rect 0 24850 800 24880
rect 4061 24850 4127 24853
rect 0 24848 4127 24850
rect 0 24792 4066 24848
rect 4122 24792 4127 24848
rect 0 24790 4127 24792
rect 0 24760 800 24790
rect 4061 24787 4127 24790
rect 4797 24850 4863 24853
rect 21173 24850 21239 24853
rect 4797 24848 21239 24850
rect 4797 24792 4802 24848
rect 4858 24792 21178 24848
rect 21234 24792 21239 24848
rect 4797 24790 21239 24792
rect 4797 24787 4863 24790
rect 21173 24787 21239 24790
rect 48313 24850 48379 24853
rect 50200 24850 51000 24880
rect 48313 24848 51000 24850
rect 48313 24792 48318 24848
rect 48374 24792 51000 24848
rect 48313 24790 51000 24792
rect 48313 24787 48379 24790
rect 50200 24760 51000 24790
rect 16297 24714 16363 24717
rect 27153 24714 27219 24717
rect 16297 24712 27219 24714
rect 16297 24656 16302 24712
rect 16358 24656 27158 24712
rect 27214 24656 27219 24712
rect 16297 24654 27219 24656
rect 16297 24651 16363 24654
rect 27153 24651 27219 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 21633 24442 21699 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 16990 24440 21699 24442
rect 16990 24384 21638 24440
rect 21694 24384 21699 24440
rect 16990 24382 21699 24384
rect 11053 24306 11119 24309
rect 16990 24306 17050 24382
rect 21633 24379 21699 24382
rect 11053 24304 17050 24306
rect 11053 24248 11058 24304
rect 11114 24248 17050 24304
rect 11053 24246 17050 24248
rect 17585 24306 17651 24309
rect 18965 24306 19031 24309
rect 17585 24304 19031 24306
rect 17585 24248 17590 24304
rect 17646 24248 18970 24304
rect 19026 24248 19031 24304
rect 17585 24246 19031 24248
rect 11053 24243 11119 24246
rect 17585 24243 17651 24246
rect 18965 24243 19031 24246
rect 20805 24306 20871 24309
rect 40125 24306 40191 24309
rect 20805 24304 40191 24306
rect 20805 24248 20810 24304
rect 20866 24248 40130 24304
rect 40186 24248 40191 24304
rect 20805 24246 40191 24248
rect 20805 24243 20871 24246
rect 40125 24243 40191 24246
rect 9213 24170 9279 24173
rect 35065 24170 35131 24173
rect 9213 24168 35131 24170
rect 9213 24112 9218 24168
rect 9274 24112 35070 24168
rect 35126 24112 35131 24168
rect 9213 24110 35131 24112
rect 9213 24107 9279 24110
rect 35065 24107 35131 24110
rect 0 24034 800 24064
rect 3877 24034 3943 24037
rect 0 24032 3943 24034
rect 0 23976 3882 24032
rect 3938 23976 3943 24032
rect 0 23974 3943 23976
rect 0 23944 800 23974
rect 3877 23971 3943 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 20161 23898 20227 23901
rect 22277 23898 22343 23901
rect 20161 23896 22343 23898
rect 20161 23840 20166 23896
rect 20222 23840 22282 23896
rect 22338 23840 22343 23896
rect 20161 23838 22343 23840
rect 20161 23835 20227 23838
rect 22277 23835 22343 23838
rect 36261 23898 36327 23901
rect 36537 23898 36603 23901
rect 36261 23896 36603 23898
rect 36261 23840 36266 23896
rect 36322 23840 36542 23896
rect 36598 23840 36603 23896
rect 36261 23838 36603 23840
rect 36261 23835 36327 23838
rect 36537 23835 36603 23838
rect 49233 23898 49299 23901
rect 50200 23898 51000 23928
rect 49233 23896 51000 23898
rect 49233 23840 49238 23896
rect 49294 23840 51000 23896
rect 49233 23838 51000 23840
rect 49233 23835 49299 23838
rect 50200 23808 51000 23838
rect 8293 23762 8359 23765
rect 9806 23762 9812 23764
rect 8293 23760 9812 23762
rect 8293 23704 8298 23760
rect 8354 23704 9812 23760
rect 8293 23702 9812 23704
rect 8293 23699 8359 23702
rect 9806 23700 9812 23702
rect 9876 23700 9882 23764
rect 13629 23762 13695 23765
rect 33409 23762 33475 23765
rect 13629 23760 33475 23762
rect 13629 23704 13634 23760
rect 13690 23704 33414 23760
rect 33470 23704 33475 23760
rect 13629 23702 33475 23704
rect 13629 23699 13695 23702
rect 33409 23699 33475 23702
rect 0 23626 800 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 800 23566
rect 4061 23563 4127 23566
rect 13261 23626 13327 23629
rect 19793 23626 19859 23629
rect 13261 23624 19859 23626
rect 13261 23568 13266 23624
rect 13322 23568 19798 23624
rect 19854 23568 19859 23624
rect 13261 23566 19859 23568
rect 13261 23563 13327 23566
rect 19793 23563 19859 23566
rect 22277 23626 22343 23629
rect 38653 23626 38719 23629
rect 22277 23624 38719 23626
rect 22277 23568 22282 23624
rect 22338 23568 38658 23624
rect 38714 23568 38719 23624
rect 22277 23566 38719 23568
rect 22277 23563 22343 23566
rect 38653 23563 38719 23566
rect 2129 23490 2195 23493
rect 2262 23490 2268 23492
rect 2129 23488 2268 23490
rect 2129 23432 2134 23488
rect 2190 23432 2268 23488
rect 2129 23430 2268 23432
rect 2129 23427 2195 23430
rect 2262 23428 2268 23430
rect 2332 23428 2338 23492
rect 4286 23428 4292 23492
rect 4356 23490 4362 23492
rect 7465 23490 7531 23493
rect 4356 23488 7531 23490
rect 4356 23432 7470 23488
rect 7526 23432 7531 23488
rect 4356 23430 7531 23432
rect 4356 23428 4362 23430
rect 7465 23427 7531 23430
rect 13537 23490 13603 23493
rect 21909 23490 21975 23493
rect 22185 23492 22251 23493
rect 22134 23490 22140 23492
rect 13537 23488 21975 23490
rect 13537 23432 13542 23488
rect 13598 23432 21914 23488
rect 21970 23432 21975 23488
rect 13537 23430 21975 23432
rect 22094 23430 22140 23490
rect 22204 23488 22251 23492
rect 22246 23432 22251 23488
rect 13537 23427 13603 23430
rect 21909 23427 21975 23430
rect 22134 23428 22140 23430
rect 22204 23428 22251 23432
rect 22185 23427 22251 23428
rect 25405 23490 25471 23493
rect 26785 23490 26851 23493
rect 25405 23488 26851 23490
rect 25405 23432 25410 23488
rect 25466 23432 26790 23488
rect 26846 23432 26851 23488
rect 25405 23430 26851 23432
rect 25405 23427 25471 23430
rect 26785 23427 26851 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 14181 23354 14247 23357
rect 14457 23354 14523 23357
rect 22737 23354 22803 23357
rect 14181 23352 22803 23354
rect 14181 23296 14186 23352
rect 14242 23296 14462 23352
rect 14518 23296 22742 23352
rect 22798 23296 22803 23352
rect 14181 23294 22803 23296
rect 14181 23291 14247 23294
rect 14457 23291 14523 23294
rect 22737 23291 22803 23294
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 4245 23218 4311 23221
rect 5574 23218 5580 23220
rect 4245 23216 5580 23218
rect 4245 23160 4250 23216
rect 4306 23160 5580 23216
rect 4245 23158 5580 23160
rect 4245 23155 4311 23158
rect 5574 23156 5580 23158
rect 5644 23218 5650 23220
rect 17953 23218 18019 23221
rect 5644 23216 18019 23218
rect 5644 23160 17958 23216
rect 18014 23160 18019 23216
rect 5644 23158 18019 23160
rect 5644 23156 5650 23158
rect 17953 23155 18019 23158
rect 19425 23218 19491 23221
rect 33593 23218 33659 23221
rect 19425 23216 33659 23218
rect 19425 23160 19430 23216
rect 19486 23160 33598 23216
rect 33654 23160 33659 23216
rect 19425 23158 33659 23160
rect 19425 23155 19491 23158
rect 33593 23155 33659 23158
rect 7414 23020 7420 23084
rect 7484 23082 7490 23084
rect 7925 23082 7991 23085
rect 7484 23080 7991 23082
rect 7484 23024 7930 23080
rect 7986 23024 7991 23080
rect 7484 23022 7991 23024
rect 7484 23020 7490 23022
rect 7925 23019 7991 23022
rect 14365 23082 14431 23085
rect 34881 23082 34947 23085
rect 14365 23080 34947 23082
rect 14365 23024 14370 23080
rect 14426 23024 34886 23080
rect 34942 23024 34947 23080
rect 14365 23022 34947 23024
rect 14365 23019 14431 23022
rect 34881 23019 34947 23022
rect 22737 22946 22803 22949
rect 24761 22946 24827 22949
rect 22737 22944 24827 22946
rect 22737 22888 22742 22944
rect 22798 22888 24766 22944
rect 24822 22888 24827 22944
rect 22737 22886 24827 22888
rect 22737 22883 22803 22886
rect 24761 22883 24827 22886
rect 49049 22946 49115 22949
rect 50200 22946 51000 22976
rect 49049 22944 51000 22946
rect 49049 22888 49054 22944
rect 49110 22888 51000 22944
rect 49049 22886 51000 22888
rect 49049 22883 49115 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 50200 22856 51000 22886
rect 47946 22815 48262 22816
rect 3601 22810 3667 22813
rect 0 22808 3667 22810
rect 0 22752 3606 22808
rect 3662 22752 3667 22808
rect 0 22750 3667 22752
rect 0 22720 800 22750
rect 3601 22747 3667 22750
rect 19609 22810 19675 22813
rect 24945 22810 25011 22813
rect 19609 22808 25011 22810
rect 19609 22752 19614 22808
rect 19670 22752 24950 22808
rect 25006 22752 25011 22808
rect 19609 22750 25011 22752
rect 19609 22747 19675 22750
rect 24945 22747 25011 22750
rect 4153 22674 4219 22677
rect 7189 22676 7255 22677
rect 5390 22674 5396 22676
rect 4153 22672 5396 22674
rect 4153 22616 4158 22672
rect 4214 22616 5396 22672
rect 4153 22614 5396 22616
rect 4153 22611 4219 22614
rect 5390 22612 5396 22614
rect 5460 22612 5466 22676
rect 7189 22672 7236 22676
rect 7300 22674 7306 22676
rect 17769 22674 17835 22677
rect 23933 22674 23999 22677
rect 7189 22616 7194 22672
rect 7189 22612 7236 22616
rect 7300 22614 7346 22674
rect 17769 22672 23999 22674
rect 17769 22616 17774 22672
rect 17830 22616 23938 22672
rect 23994 22616 23999 22672
rect 17769 22614 23999 22616
rect 7300 22612 7306 22614
rect 7189 22611 7255 22612
rect 17769 22611 17835 22614
rect 23933 22611 23999 22614
rect 27429 22674 27495 22677
rect 30925 22674 30991 22677
rect 33869 22674 33935 22677
rect 27429 22672 30991 22674
rect 27429 22616 27434 22672
rect 27490 22616 30930 22672
rect 30986 22616 30991 22672
rect 27429 22614 30991 22616
rect 27429 22611 27495 22614
rect 30925 22611 30991 22614
rect 31710 22672 33935 22674
rect 31710 22616 33874 22672
rect 33930 22616 33935 22672
rect 31710 22614 33935 22616
rect 4061 22538 4127 22541
rect 2270 22536 4127 22538
rect 2270 22480 4066 22536
rect 4122 22480 4127 22536
rect 2270 22478 4127 22480
rect 0 22402 800 22432
rect 2270 22402 2330 22478
rect 4061 22475 4127 22478
rect 11145 22538 11211 22541
rect 17166 22538 17172 22540
rect 11145 22536 17172 22538
rect 11145 22480 11150 22536
rect 11206 22480 17172 22536
rect 11145 22478 17172 22480
rect 11145 22475 11211 22478
rect 17166 22476 17172 22478
rect 17236 22476 17242 22540
rect 17769 22538 17835 22541
rect 31710 22538 31770 22614
rect 33869 22611 33935 22614
rect 17769 22536 31770 22538
rect 17769 22480 17774 22536
rect 17830 22480 31770 22536
rect 17769 22478 31770 22480
rect 17769 22475 17835 22478
rect 0 22342 2330 22402
rect 3785 22402 3851 22405
rect 3918 22402 3924 22404
rect 3785 22400 3924 22402
rect 3785 22344 3790 22400
rect 3846 22344 3924 22400
rect 3785 22342 3924 22344
rect 0 22312 800 22342
rect 3785 22339 3851 22342
rect 3918 22340 3924 22342
rect 3988 22340 3994 22404
rect 15009 22402 15075 22405
rect 21817 22402 21883 22405
rect 15009 22400 21883 22402
rect 15009 22344 15014 22400
rect 15070 22344 21822 22400
rect 21878 22344 21883 22400
rect 15009 22342 21883 22344
rect 15009 22339 15075 22342
rect 21817 22339 21883 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 17166 22204 17172 22268
rect 17236 22266 17242 22268
rect 23749 22266 23815 22269
rect 26509 22266 26575 22269
rect 27061 22266 27127 22269
rect 27521 22266 27587 22269
rect 30649 22266 30715 22269
rect 17236 22206 22110 22266
rect 17236 22204 17242 22206
rect 5993 22130 6059 22133
rect 9397 22130 9463 22133
rect 5993 22128 9463 22130
rect 5993 22072 5998 22128
rect 6054 22072 9402 22128
rect 9458 22072 9463 22128
rect 5993 22070 9463 22072
rect 22050 22130 22110 22206
rect 23749 22264 30715 22266
rect 23749 22208 23754 22264
rect 23810 22208 26514 22264
rect 26570 22208 27066 22264
rect 27122 22208 27526 22264
rect 27582 22208 30654 22264
rect 30710 22208 30715 22264
rect 23749 22206 30715 22208
rect 23749 22203 23815 22206
rect 26509 22203 26575 22206
rect 27061 22203 27127 22206
rect 27521 22203 27587 22206
rect 30649 22203 30715 22206
rect 32489 22130 32555 22133
rect 22050 22128 32555 22130
rect 22050 22072 32494 22128
rect 32550 22072 32555 22128
rect 22050 22070 32555 22072
rect 5993 22067 6059 22070
rect 9397 22067 9463 22070
rect 32489 22067 32555 22070
rect 0 21994 800 22024
rect 4245 21994 4311 21997
rect 0 21992 4311 21994
rect 0 21936 4250 21992
rect 4306 21936 4311 21992
rect 0 21934 4311 21936
rect 0 21904 800 21934
rect 4245 21931 4311 21934
rect 8753 21994 8819 21997
rect 14641 21994 14707 21997
rect 8753 21992 14707 21994
rect 8753 21936 8758 21992
rect 8814 21936 14646 21992
rect 14702 21936 14707 21992
rect 8753 21934 14707 21936
rect 8753 21931 8819 21934
rect 14641 21931 14707 21934
rect 16757 21994 16823 21997
rect 30005 21994 30071 21997
rect 16757 21992 30071 21994
rect 16757 21936 16762 21992
rect 16818 21936 30010 21992
rect 30066 21936 30071 21992
rect 16757 21934 30071 21936
rect 16757 21931 16823 21934
rect 30005 21931 30071 21934
rect 49049 21994 49115 21997
rect 50200 21994 51000 22024
rect 49049 21992 51000 21994
rect 49049 21936 49054 21992
rect 49110 21936 51000 21992
rect 49049 21934 51000 21936
rect 49049 21931 49115 21934
rect 50200 21904 51000 21934
rect 9673 21858 9739 21861
rect 10542 21858 10548 21860
rect 9673 21856 10548 21858
rect 9673 21800 9678 21856
rect 9734 21800 10548 21856
rect 9673 21798 10548 21800
rect 9673 21795 9739 21798
rect 10542 21796 10548 21798
rect 10612 21796 10618 21860
rect 10961 21858 11027 21861
rect 16941 21858 17007 21861
rect 17769 21858 17835 21861
rect 10961 21856 17835 21858
rect 10961 21800 10966 21856
rect 11022 21800 16946 21856
rect 17002 21800 17774 21856
rect 17830 21800 17835 21856
rect 10961 21798 17835 21800
rect 10961 21795 11027 21798
rect 16941 21795 17007 21798
rect 17769 21795 17835 21798
rect 22686 21796 22692 21860
rect 22756 21858 22762 21860
rect 23289 21858 23355 21861
rect 22756 21856 23355 21858
rect 22756 21800 23294 21856
rect 23350 21800 23355 21856
rect 22756 21798 23355 21800
rect 22756 21796 22762 21798
rect 23289 21795 23355 21798
rect 29913 21858 29979 21861
rect 31109 21858 31175 21861
rect 29913 21856 31175 21858
rect 29913 21800 29918 21856
rect 29974 21800 31114 21856
rect 31170 21800 31175 21856
rect 29913 21798 31175 21800
rect 29913 21795 29979 21798
rect 31109 21795 31175 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 3601 21722 3667 21725
rect 7281 21722 7347 21725
rect 3601 21720 7347 21722
rect 3601 21664 3606 21720
rect 3662 21664 7286 21720
rect 7342 21664 7347 21720
rect 3601 21662 7347 21664
rect 3601 21659 3667 21662
rect 7281 21659 7347 21662
rect 15745 21722 15811 21725
rect 15929 21722 15995 21725
rect 15745 21720 15995 21722
rect 15745 21664 15750 21720
rect 15806 21664 15934 21720
rect 15990 21664 15995 21720
rect 15745 21662 15995 21664
rect 15745 21659 15811 21662
rect 15929 21659 15995 21662
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 3233 21586 3299 21589
rect 10501 21586 10567 21589
rect 3233 21584 10567 21586
rect 3233 21528 3238 21584
rect 3294 21528 10506 21584
rect 10562 21528 10567 21584
rect 3233 21526 10567 21528
rect 3233 21523 3299 21526
rect 10501 21523 10567 21526
rect 15929 21586 15995 21589
rect 36169 21586 36235 21589
rect 15929 21584 36235 21586
rect 15929 21528 15934 21584
rect 15990 21528 36174 21584
rect 36230 21528 36235 21584
rect 15929 21526 36235 21528
rect 15929 21523 15995 21526
rect 36169 21523 36235 21526
rect 2865 21450 2931 21453
rect 2730 21448 2931 21450
rect 2730 21392 2870 21448
rect 2926 21392 2931 21448
rect 2730 21390 2931 21392
rect 0 21178 800 21208
rect 2730 21178 2790 21390
rect 2865 21387 2931 21390
rect 5625 21450 5691 21453
rect 5758 21450 5764 21452
rect 5625 21448 5764 21450
rect 5625 21392 5630 21448
rect 5686 21392 5764 21448
rect 5625 21390 5764 21392
rect 5625 21387 5691 21390
rect 5758 21388 5764 21390
rect 5828 21388 5834 21452
rect 7557 21450 7623 21453
rect 8937 21450 9003 21453
rect 7557 21448 9003 21450
rect 7557 21392 7562 21448
rect 7618 21392 8942 21448
rect 8998 21392 9003 21448
rect 7557 21390 9003 21392
rect 5766 21314 5826 21388
rect 7557 21387 7623 21390
rect 8937 21387 9003 21390
rect 15561 21450 15627 21453
rect 31109 21450 31175 21453
rect 15561 21448 31175 21450
rect 15561 21392 15566 21448
rect 15622 21392 31114 21448
rect 31170 21392 31175 21448
rect 15561 21390 31175 21392
rect 15561 21387 15627 21390
rect 31109 21387 31175 21390
rect 26233 21314 26299 21317
rect 28717 21314 28783 21317
rect 5766 21254 12266 21314
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 0 21118 2790 21178
rect 7005 21178 7071 21181
rect 11605 21178 11671 21181
rect 7005 21176 11671 21178
rect 7005 21120 7010 21176
rect 7066 21120 11610 21176
rect 11666 21120 11671 21176
rect 7005 21118 11671 21120
rect 12206 21178 12266 21254
rect 26233 21312 28783 21314
rect 26233 21256 26238 21312
rect 26294 21256 28722 21312
rect 28778 21256 28783 21312
rect 26233 21254 28783 21256
rect 26233 21251 26299 21254
rect 28717 21251 28783 21254
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 12341 21178 12407 21181
rect 12206 21176 12407 21178
rect 12206 21120 12346 21176
rect 12402 21120 12407 21176
rect 12206 21118 12407 21120
rect 0 21088 800 21118
rect 7005 21115 7071 21118
rect 11605 21115 11671 21118
rect 12341 21115 12407 21118
rect 13905 21178 13971 21181
rect 18597 21178 18663 21181
rect 13905 21176 18663 21178
rect 13905 21120 13910 21176
rect 13966 21120 18602 21176
rect 18658 21120 18663 21176
rect 13905 21118 18663 21120
rect 13905 21115 13971 21118
rect 18597 21115 18663 21118
rect 4245 21042 4311 21045
rect 32213 21042 32279 21045
rect 4245 21040 32279 21042
rect 4245 20984 4250 21040
rect 4306 20984 32218 21040
rect 32274 20984 32279 21040
rect 4245 20982 32279 20984
rect 4245 20979 4311 20982
rect 32213 20979 32279 20982
rect 49141 21042 49207 21045
rect 50200 21042 51000 21072
rect 49141 21040 51000 21042
rect 49141 20984 49146 21040
rect 49202 20984 51000 21040
rect 49141 20982 51000 20984
rect 49141 20979 49207 20982
rect 50200 20952 51000 20982
rect 5625 20906 5691 20909
rect 7005 20906 7071 20909
rect 5625 20904 7071 20906
rect 5625 20848 5630 20904
rect 5686 20848 7010 20904
rect 7066 20848 7071 20904
rect 5625 20846 7071 20848
rect 5625 20843 5691 20846
rect 7005 20843 7071 20846
rect 8201 20906 8267 20909
rect 15745 20906 15811 20909
rect 8201 20904 15811 20906
rect 8201 20848 8206 20904
rect 8262 20848 15750 20904
rect 15806 20848 15811 20904
rect 8201 20846 15811 20848
rect 8201 20843 8267 20846
rect 15745 20843 15811 20846
rect 17309 20906 17375 20909
rect 17309 20904 28458 20906
rect 17309 20848 17314 20904
rect 17370 20848 28458 20904
rect 17309 20846 28458 20848
rect 17309 20843 17375 20846
rect 0 20770 800 20800
rect 28398 20773 28458 20846
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 3734 20708 3740 20772
rect 3804 20770 3810 20772
rect 3969 20770 4035 20773
rect 3804 20768 4035 20770
rect 3804 20712 3974 20768
rect 4030 20712 4035 20768
rect 3804 20710 4035 20712
rect 3804 20708 3810 20710
rect 3969 20707 4035 20710
rect 6310 20708 6316 20772
rect 6380 20770 6386 20772
rect 6453 20770 6519 20773
rect 6380 20768 6519 20770
rect 6380 20712 6458 20768
rect 6514 20712 6519 20768
rect 6380 20710 6519 20712
rect 6380 20708 6386 20710
rect 6453 20707 6519 20710
rect 9397 20772 9463 20773
rect 13905 20772 13971 20773
rect 9397 20768 9444 20772
rect 9508 20770 9514 20772
rect 9397 20712 9402 20768
rect 9397 20708 9444 20712
rect 9508 20710 9554 20770
rect 9508 20708 9514 20710
rect 13854 20708 13860 20772
rect 13924 20770 13971 20772
rect 19701 20770 19767 20773
rect 25405 20770 25471 20773
rect 13924 20768 14016 20770
rect 13966 20712 14016 20768
rect 13924 20710 14016 20712
rect 19701 20768 25471 20770
rect 19701 20712 19706 20768
rect 19762 20712 25410 20768
rect 25466 20712 25471 20768
rect 19701 20710 25471 20712
rect 28398 20768 28507 20773
rect 28398 20712 28446 20768
rect 28502 20712 28507 20768
rect 28398 20710 28507 20712
rect 13924 20708 13971 20710
rect 9397 20707 9463 20708
rect 13905 20707 13971 20708
rect 19701 20707 19767 20710
rect 25405 20707 25471 20710
rect 28441 20707 28507 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 17217 20634 17283 20637
rect 17769 20634 17835 20637
rect 17217 20632 17835 20634
rect 17217 20576 17222 20632
rect 17278 20576 17774 20632
rect 17830 20576 17835 20632
rect 17217 20574 17835 20576
rect 17217 20571 17283 20574
rect 17769 20571 17835 20574
rect 23657 20634 23723 20637
rect 26601 20634 26667 20637
rect 23657 20632 26667 20634
rect 23657 20576 23662 20632
rect 23718 20576 26606 20632
rect 26662 20576 26667 20632
rect 23657 20574 26667 20576
rect 23657 20571 23723 20574
rect 26601 20571 26667 20574
rect 11789 20498 11855 20501
rect 32305 20498 32371 20501
rect 11789 20496 32371 20498
rect 11789 20440 11794 20496
rect 11850 20440 32310 20496
rect 32366 20440 32371 20496
rect 11789 20438 32371 20440
rect 11789 20435 11855 20438
rect 32305 20435 32371 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 11973 20362 12039 20365
rect 13905 20362 13971 20365
rect 11973 20360 13971 20362
rect 11973 20304 11978 20360
rect 12034 20304 13910 20360
rect 13966 20304 13971 20360
rect 11973 20302 13971 20304
rect 11973 20299 12039 20302
rect 13905 20299 13971 20302
rect 17217 20362 17283 20365
rect 31845 20362 31911 20365
rect 17217 20360 31911 20362
rect 17217 20304 17222 20360
rect 17278 20304 31850 20360
rect 31906 20304 31911 20360
rect 17217 20302 31911 20304
rect 17217 20299 17283 20302
rect 31845 20299 31911 20302
rect 13537 20226 13603 20229
rect 18505 20226 18571 20229
rect 13537 20224 18571 20226
rect 13537 20168 13542 20224
rect 13598 20168 18510 20224
rect 18566 20168 18571 20224
rect 13537 20166 18571 20168
rect 13537 20163 13603 20166
rect 18505 20163 18571 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 5625 20090 5691 20093
rect 6545 20090 6611 20093
rect 16573 20090 16639 20093
rect 19793 20090 19859 20093
rect 5625 20088 12450 20090
rect 5625 20032 5630 20088
rect 5686 20032 6550 20088
rect 6606 20032 12450 20088
rect 5625 20030 12450 20032
rect 5625 20027 5691 20030
rect 6545 20027 6611 20030
rect 0 19954 800 19984
rect 2773 19954 2839 19957
rect 0 19952 2839 19954
rect 0 19896 2778 19952
rect 2834 19896 2839 19952
rect 0 19894 2839 19896
rect 0 19864 800 19894
rect 2773 19891 2839 19894
rect 4429 19954 4495 19957
rect 11421 19954 11487 19957
rect 4429 19952 11487 19954
rect 4429 19896 4434 19952
rect 4490 19896 11426 19952
rect 11482 19896 11487 19952
rect 4429 19894 11487 19896
rect 12390 19954 12450 20030
rect 16573 20088 19859 20090
rect 16573 20032 16578 20088
rect 16634 20032 19798 20088
rect 19854 20032 19859 20088
rect 16573 20030 19859 20032
rect 16573 20027 16639 20030
rect 19793 20027 19859 20030
rect 28625 19954 28691 19957
rect 12390 19952 28691 19954
rect 12390 19896 28630 19952
rect 28686 19896 28691 19952
rect 12390 19894 28691 19896
rect 4429 19891 4495 19894
rect 11421 19891 11487 19894
rect 28625 19891 28691 19894
rect 1761 19818 1827 19821
rect 9305 19818 9371 19821
rect 1761 19816 9371 19818
rect 1761 19760 1766 19816
rect 1822 19760 9310 19816
rect 9366 19760 9371 19816
rect 1761 19758 9371 19760
rect 1761 19755 1827 19758
rect 9305 19755 9371 19758
rect 12985 19818 13051 19821
rect 29177 19818 29243 19821
rect 12985 19816 29243 19818
rect 12985 19760 12990 19816
rect 13046 19760 29182 19816
rect 29238 19760 29243 19816
rect 12985 19758 29243 19760
rect 12985 19755 13051 19758
rect 29177 19755 29243 19758
rect 2773 19682 2839 19685
rect 3325 19682 3391 19685
rect 2773 19680 3391 19682
rect 2773 19624 2778 19680
rect 2834 19624 3330 19680
rect 3386 19624 3391 19680
rect 2773 19622 3391 19624
rect 2773 19619 2839 19622
rect 3325 19619 3391 19622
rect 16021 19682 16087 19685
rect 17677 19682 17743 19685
rect 16021 19680 17743 19682
rect 16021 19624 16026 19680
rect 16082 19624 17682 19680
rect 17738 19624 17743 19680
rect 16021 19622 17743 19624
rect 16021 19619 16087 19622
rect 17677 19619 17743 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2957 19546 3023 19549
rect 0 19544 3023 19546
rect 0 19488 2962 19544
rect 3018 19488 3023 19544
rect 0 19486 3023 19488
rect 0 19456 800 19486
rect 2957 19483 3023 19486
rect 17401 19546 17467 19549
rect 17677 19546 17743 19549
rect 17401 19544 17743 19546
rect 17401 19488 17406 19544
rect 17462 19488 17682 19544
rect 17738 19488 17743 19544
rect 17401 19486 17743 19488
rect 17401 19483 17467 19486
rect 17677 19483 17743 19486
rect 18505 19546 18571 19549
rect 21357 19546 21423 19549
rect 18505 19544 21423 19546
rect 18505 19488 18510 19544
rect 18566 19488 21362 19544
rect 21418 19488 21423 19544
rect 18505 19486 21423 19488
rect 18505 19483 18571 19486
rect 21357 19483 21423 19486
rect 1485 19410 1551 19413
rect 7465 19410 7531 19413
rect 1485 19408 7531 19410
rect 1485 19352 1490 19408
rect 1546 19352 7470 19408
rect 7526 19352 7531 19408
rect 1485 19350 7531 19352
rect 1485 19347 1551 19350
rect 7465 19347 7531 19350
rect 9213 19410 9279 19413
rect 9622 19410 9628 19412
rect 9213 19408 9628 19410
rect 9213 19352 9218 19408
rect 9274 19352 9628 19408
rect 9213 19350 9628 19352
rect 9213 19347 9279 19350
rect 9622 19348 9628 19350
rect 9692 19348 9698 19412
rect 11421 19410 11487 19413
rect 30649 19410 30715 19413
rect 11421 19408 30715 19410
rect 11421 19352 11426 19408
rect 11482 19352 30654 19408
rect 30710 19352 30715 19408
rect 11421 19350 30715 19352
rect 11421 19347 11487 19350
rect 30649 19347 30715 19350
rect 6545 19274 6611 19277
rect 7005 19274 7071 19277
rect 6545 19272 7071 19274
rect 6545 19216 6550 19272
rect 6606 19216 7010 19272
rect 7066 19216 7071 19272
rect 6545 19214 7071 19216
rect 6545 19211 6611 19214
rect 7005 19211 7071 19214
rect 10133 19274 10199 19277
rect 11237 19274 11303 19277
rect 10133 19272 11303 19274
rect 10133 19216 10138 19272
rect 10194 19216 11242 19272
rect 11298 19216 11303 19272
rect 10133 19214 11303 19216
rect 10133 19211 10199 19214
rect 11237 19211 11303 19214
rect 12065 19274 12131 19277
rect 15009 19274 15075 19277
rect 17217 19274 17283 19277
rect 12065 19272 17283 19274
rect 12065 19216 12070 19272
rect 12126 19216 15014 19272
rect 15070 19216 17222 19272
rect 17278 19216 17283 19272
rect 12065 19214 17283 19216
rect 12065 19211 12131 19214
rect 15009 19211 15075 19214
rect 17217 19211 17283 19214
rect 17493 19274 17559 19277
rect 27429 19274 27495 19277
rect 17493 19272 27495 19274
rect 17493 19216 17498 19272
rect 17554 19216 27434 19272
rect 27490 19216 27495 19272
rect 17493 19214 27495 19216
rect 17493 19211 17559 19214
rect 27429 19211 27495 19214
rect 0 19138 800 19168
rect 2681 19138 2747 19141
rect 0 19136 2747 19138
rect 0 19080 2686 19136
rect 2742 19080 2747 19136
rect 0 19078 2747 19080
rect 0 19048 800 19078
rect 2681 19075 2747 19078
rect 3325 19138 3391 19141
rect 12709 19138 12775 19141
rect 3325 19136 12775 19138
rect 3325 19080 3330 19136
rect 3386 19080 12714 19136
rect 12770 19080 12775 19136
rect 3325 19078 12775 19080
rect 3325 19075 3391 19078
rect 12709 19075 12775 19078
rect 16297 19138 16363 19141
rect 16849 19138 16915 19141
rect 17677 19138 17743 19141
rect 16297 19136 17743 19138
rect 16297 19080 16302 19136
rect 16358 19080 16854 19136
rect 16910 19080 17682 19136
rect 17738 19080 17743 19136
rect 16297 19078 17743 19080
rect 16297 19075 16363 19078
rect 16849 19075 16915 19078
rect 17677 19075 17743 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 31753 19002 31819 19005
rect 31342 19000 31819 19002
rect 31342 18944 31758 19000
rect 31814 18944 31819 19000
rect 31342 18942 31819 18944
rect 4521 18866 4587 18869
rect 14457 18866 14523 18869
rect 4521 18864 14523 18866
rect 4521 18808 4526 18864
rect 4582 18808 14462 18864
rect 14518 18808 14523 18864
rect 4521 18806 14523 18808
rect 4521 18803 4587 18806
rect 14457 18803 14523 18806
rect 18505 18866 18571 18869
rect 31201 18866 31267 18869
rect 18505 18864 31267 18866
rect 18505 18808 18510 18864
rect 18566 18808 31206 18864
rect 31262 18808 31267 18864
rect 18505 18806 31267 18808
rect 18505 18803 18571 18806
rect 31201 18803 31267 18806
rect 0 18730 800 18760
rect 2865 18730 2931 18733
rect 0 18728 2931 18730
rect 0 18672 2870 18728
rect 2926 18672 2931 18728
rect 0 18670 2931 18672
rect 0 18640 800 18670
rect 2865 18667 2931 18670
rect 6085 18730 6151 18733
rect 8569 18730 8635 18733
rect 9121 18732 9187 18733
rect 6085 18728 8635 18730
rect 6085 18672 6090 18728
rect 6146 18672 8574 18728
rect 8630 18672 8635 18728
rect 6085 18670 8635 18672
rect 6085 18667 6151 18670
rect 8569 18667 8635 18670
rect 9070 18668 9076 18732
rect 9140 18730 9187 18732
rect 15837 18730 15903 18733
rect 23381 18730 23447 18733
rect 31342 18730 31402 18942
rect 31753 18939 31819 18942
rect 45369 18730 45435 18733
rect 9140 18728 9232 18730
rect 9182 18672 9232 18728
rect 9140 18670 9232 18672
rect 15837 18728 23447 18730
rect 15837 18672 15842 18728
rect 15898 18672 23386 18728
rect 23442 18672 23447 18728
rect 15837 18670 23447 18672
rect 9140 18668 9187 18670
rect 9121 18667 9187 18668
rect 15837 18667 15903 18670
rect 23381 18667 23447 18670
rect 24902 18670 31402 18730
rect 31710 18728 45435 18730
rect 31710 18672 45374 18728
rect 45430 18672 45435 18728
rect 31710 18670 45435 18672
rect 4705 18594 4771 18597
rect 6177 18594 6243 18597
rect 4705 18592 6243 18594
rect 4705 18536 4710 18592
rect 4766 18536 6182 18592
rect 6238 18536 6243 18592
rect 4705 18534 6243 18536
rect 4705 18531 4771 18534
rect 6177 18531 6243 18534
rect 18689 18594 18755 18597
rect 24209 18594 24275 18597
rect 24902 18594 24962 18670
rect 18689 18592 24962 18594
rect 18689 18536 18694 18592
rect 18750 18536 24214 18592
rect 24270 18536 24962 18592
rect 18689 18534 24962 18536
rect 18689 18531 18755 18534
rect 24209 18531 24275 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 14825 18458 14891 18461
rect 17769 18458 17835 18461
rect 14825 18456 17835 18458
rect 14825 18400 14830 18456
rect 14886 18400 17774 18456
rect 17830 18400 17835 18456
rect 14825 18398 17835 18400
rect 14825 18395 14891 18398
rect 17769 18395 17835 18398
rect 21449 18458 21515 18461
rect 23749 18458 23815 18461
rect 21449 18456 23815 18458
rect 21449 18400 21454 18456
rect 21510 18400 23754 18456
rect 23810 18400 23815 18456
rect 21449 18398 23815 18400
rect 21449 18395 21515 18398
rect 23749 18395 23815 18398
rect 24945 18458 25011 18461
rect 24945 18456 25330 18458
rect 24945 18400 24950 18456
rect 25006 18400 25330 18456
rect 24945 18398 25330 18400
rect 24945 18395 25011 18398
rect 0 18322 800 18352
rect 2773 18322 2839 18325
rect 0 18320 2839 18322
rect 0 18264 2778 18320
rect 2834 18264 2839 18320
rect 0 18262 2839 18264
rect 0 18232 800 18262
rect 2773 18259 2839 18262
rect 7557 18322 7623 18325
rect 9673 18322 9739 18325
rect 7557 18320 9739 18322
rect 7557 18264 7562 18320
rect 7618 18264 9678 18320
rect 9734 18264 9739 18320
rect 7557 18262 9739 18264
rect 7557 18259 7623 18262
rect 9673 18259 9739 18262
rect 15009 18322 15075 18325
rect 25129 18322 25195 18325
rect 15009 18320 25195 18322
rect 15009 18264 15014 18320
rect 15070 18264 25134 18320
rect 25190 18264 25195 18320
rect 15009 18262 25195 18264
rect 25270 18322 25330 18398
rect 31710 18322 31770 18670
rect 45369 18667 45435 18670
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 25270 18262 31770 18322
rect 15009 18259 15075 18262
rect 25129 18259 25195 18262
rect 2773 18186 2839 18189
rect 3325 18186 3391 18189
rect 2773 18184 3391 18186
rect 2773 18128 2778 18184
rect 2834 18128 3330 18184
rect 3386 18128 3391 18184
rect 2773 18126 3391 18128
rect 2773 18123 2839 18126
rect 3325 18123 3391 18126
rect 12157 18186 12223 18189
rect 32673 18186 32739 18189
rect 12157 18184 32739 18186
rect 12157 18128 12162 18184
rect 12218 18128 32678 18184
rect 32734 18128 32739 18184
rect 12157 18126 32739 18128
rect 12157 18123 12223 18126
rect 32673 18123 32739 18126
rect 5257 18052 5323 18053
rect 5206 18050 5212 18052
rect 5166 17990 5212 18050
rect 5276 18048 5323 18052
rect 5318 17992 5323 18048
rect 5206 17988 5212 17990
rect 5276 17988 5323 17992
rect 5257 17987 5323 17988
rect 5625 18050 5691 18053
rect 5942 18050 5948 18052
rect 5625 18048 5948 18050
rect 5625 17992 5630 18048
rect 5686 17992 5948 18048
rect 5625 17990 5948 17992
rect 5625 17987 5691 17990
rect 5942 17988 5948 17990
rect 6012 17988 6018 18052
rect 6085 18050 6151 18053
rect 9489 18050 9555 18053
rect 6085 18048 9555 18050
rect 6085 17992 6090 18048
rect 6146 17992 9494 18048
rect 9550 17992 9555 18048
rect 6085 17990 9555 17992
rect 6085 17987 6151 17990
rect 9489 17987 9555 17990
rect 15377 18050 15443 18053
rect 16481 18050 16547 18053
rect 18965 18050 19031 18053
rect 15377 18048 19031 18050
rect 15377 17992 15382 18048
rect 15438 17992 16486 18048
rect 16542 17992 18970 18048
rect 19026 17992 19031 18048
rect 15377 17990 19031 17992
rect 15377 17987 15443 17990
rect 16481 17987 16547 17990
rect 18965 17987 19031 17990
rect 23381 18050 23447 18053
rect 30649 18050 30715 18053
rect 23381 18048 30715 18050
rect 23381 17992 23386 18048
rect 23442 17992 30654 18048
rect 30710 17992 30715 18048
rect 23381 17990 30715 17992
rect 23381 17987 23447 17990
rect 30649 17987 30715 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 3417 17914 3483 17917
rect 7189 17914 7255 17917
rect 11646 17914 11652 17916
rect 3417 17912 11652 17914
rect 3417 17856 3422 17912
rect 3478 17856 7194 17912
rect 7250 17856 11652 17912
rect 3417 17854 11652 17856
rect 3417 17851 3483 17854
rect 7189 17851 7255 17854
rect 11646 17852 11652 17854
rect 11716 17852 11722 17916
rect 14181 17914 14247 17917
rect 20069 17914 20135 17917
rect 14181 17912 20135 17914
rect 14181 17856 14186 17912
rect 14242 17856 20074 17912
rect 20130 17856 20135 17912
rect 14181 17854 20135 17856
rect 14181 17851 14247 17854
rect 20069 17851 20135 17854
rect 7465 17778 7531 17781
rect 7598 17778 7604 17780
rect 7465 17776 7604 17778
rect 7465 17720 7470 17776
rect 7526 17720 7604 17776
rect 7465 17718 7604 17720
rect 7465 17715 7531 17718
rect 7598 17716 7604 17718
rect 7668 17716 7674 17780
rect 10869 17778 10935 17781
rect 13261 17778 13327 17781
rect 10869 17776 13327 17778
rect 10869 17720 10874 17776
rect 10930 17720 13266 17776
rect 13322 17720 13327 17776
rect 10869 17718 13327 17720
rect 10869 17715 10935 17718
rect 13261 17715 13327 17718
rect 17125 17778 17191 17781
rect 24301 17778 24367 17781
rect 17125 17776 24367 17778
rect 17125 17720 17130 17776
rect 17186 17720 24306 17776
rect 24362 17720 24367 17776
rect 17125 17718 24367 17720
rect 17125 17715 17191 17718
rect 24301 17715 24367 17718
rect 4797 17642 4863 17645
rect 11697 17642 11763 17645
rect 16941 17642 17007 17645
rect 20989 17642 21055 17645
rect 4797 17640 9506 17642
rect 4797 17584 4802 17640
rect 4858 17584 9506 17640
rect 4797 17582 9506 17584
rect 4797 17579 4863 17582
rect 0 17506 800 17536
rect 2037 17506 2103 17509
rect 0 17504 2103 17506
rect 0 17448 2042 17504
rect 2098 17448 2103 17504
rect 0 17446 2103 17448
rect 0 17416 800 17446
rect 2037 17443 2103 17446
rect 4245 17506 4311 17509
rect 7465 17506 7531 17509
rect 4245 17504 7531 17506
rect 4245 17448 4250 17504
rect 4306 17448 7470 17504
rect 7526 17448 7531 17504
rect 4245 17446 7531 17448
rect 4245 17443 4311 17446
rect 7465 17443 7531 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 9446 17373 9506 17582
rect 11697 17640 17007 17642
rect 11697 17584 11702 17640
rect 11758 17584 16946 17640
rect 17002 17584 17007 17640
rect 11697 17582 17007 17584
rect 11697 17579 11763 17582
rect 16941 17579 17007 17582
rect 17772 17640 21055 17642
rect 17772 17584 20994 17640
rect 21050 17584 21055 17640
rect 17772 17582 21055 17584
rect 10777 17506 10843 17509
rect 17772 17506 17832 17582
rect 20989 17579 21055 17582
rect 25681 17642 25747 17645
rect 44633 17642 44699 17645
rect 25681 17640 44699 17642
rect 25681 17584 25686 17640
rect 25742 17584 44638 17640
rect 44694 17584 44699 17640
rect 25681 17582 44699 17584
rect 25681 17579 25747 17582
rect 44633 17579 44699 17582
rect 10777 17504 17832 17506
rect 10777 17448 10782 17504
rect 10838 17448 17832 17504
rect 10777 17446 17832 17448
rect 19793 17506 19859 17509
rect 23657 17506 23723 17509
rect 19793 17504 23723 17506
rect 19793 17448 19798 17504
rect 19854 17448 23662 17504
rect 23718 17448 23723 17504
rect 19793 17446 23723 17448
rect 10777 17443 10843 17446
rect 19793 17443 19859 17446
rect 23657 17443 23723 17446
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 9305 17372 9371 17373
rect 9254 17370 9260 17372
rect 9214 17310 9260 17370
rect 9324 17368 9371 17372
rect 9366 17312 9371 17368
rect 9254 17308 9260 17310
rect 9324 17308 9371 17312
rect 9446 17368 9555 17373
rect 9446 17312 9494 17368
rect 9550 17312 9555 17368
rect 9446 17310 9555 17312
rect 9305 17307 9371 17308
rect 9489 17307 9555 17310
rect 10409 17370 10475 17373
rect 16757 17370 16823 17373
rect 10409 17368 16823 17370
rect 10409 17312 10414 17368
rect 10470 17312 16762 17368
rect 16818 17312 16823 17368
rect 10409 17310 16823 17312
rect 10409 17307 10475 17310
rect 16757 17307 16823 17310
rect 8109 17234 8175 17237
rect 18505 17234 18571 17237
rect 8109 17232 18571 17234
rect 8109 17176 8114 17232
rect 8170 17176 18510 17232
rect 18566 17176 18571 17232
rect 8109 17174 18571 17176
rect 8109 17171 8175 17174
rect 18505 17171 18571 17174
rect 21817 17234 21883 17237
rect 23841 17234 23907 17237
rect 21817 17232 23907 17234
rect 21817 17176 21822 17232
rect 21878 17176 23846 17232
rect 23902 17176 23907 17232
rect 21817 17174 23907 17176
rect 21817 17171 21883 17174
rect 23841 17171 23907 17174
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 5073 17098 5139 17101
rect 8201 17098 8267 17101
rect 18597 17098 18663 17101
rect 21909 17098 21975 17101
rect 28533 17098 28599 17101
rect 5073 17096 16866 17098
rect 5073 17040 5078 17096
rect 5134 17040 8206 17096
rect 8262 17040 16866 17096
rect 5073 17038 16866 17040
rect 5073 17035 5139 17038
rect 8201 17035 8267 17038
rect 4705 16962 4771 16965
rect 12801 16962 12867 16965
rect 4705 16960 12867 16962
rect 4705 16904 4710 16960
rect 4766 16904 12806 16960
rect 12862 16904 12867 16960
rect 4705 16902 12867 16904
rect 4705 16899 4771 16902
rect 12801 16899 12867 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 3693 16826 3759 16829
rect 9070 16826 9076 16828
rect 3693 16824 9076 16826
rect 3693 16768 3698 16824
rect 3754 16768 9076 16824
rect 3693 16766 9076 16768
rect 3693 16763 3759 16766
rect 9070 16764 9076 16766
rect 9140 16826 9146 16828
rect 9213 16826 9279 16829
rect 11697 16828 11763 16829
rect 9140 16824 9279 16826
rect 9140 16768 9218 16824
rect 9274 16768 9279 16824
rect 9140 16766 9279 16768
rect 9140 16764 9146 16766
rect 9213 16763 9279 16766
rect 11646 16764 11652 16828
rect 11716 16826 11763 16828
rect 16806 16826 16866 17038
rect 18597 17096 21975 17098
rect 18597 17040 18602 17096
rect 18658 17040 21914 17096
rect 21970 17040 21975 17096
rect 18597 17038 21975 17040
rect 18597 17035 18663 17038
rect 21909 17035 21975 17038
rect 22050 17096 28599 17098
rect 22050 17040 28538 17096
rect 28594 17040 28599 17096
rect 22050 17038 28599 17040
rect 16941 16962 17007 16965
rect 20345 16962 20411 16965
rect 16941 16960 20411 16962
rect 16941 16904 16946 16960
rect 17002 16904 20350 16960
rect 20406 16904 20411 16960
rect 16941 16902 20411 16904
rect 16941 16899 17007 16902
rect 20345 16899 20411 16902
rect 18781 16826 18847 16829
rect 21909 16826 21975 16829
rect 11716 16824 11808 16826
rect 11758 16768 11808 16824
rect 11716 16766 11808 16768
rect 16806 16824 21975 16826
rect 16806 16768 18786 16824
rect 18842 16768 21914 16824
rect 21970 16768 21975 16824
rect 16806 16766 21975 16768
rect 11716 16764 11763 16766
rect 11697 16763 11763 16764
rect 18781 16763 18847 16766
rect 21909 16763 21975 16766
rect 0 16690 800 16720
rect 1117 16690 1183 16693
rect 0 16688 1183 16690
rect 0 16632 1122 16688
rect 1178 16632 1183 16688
rect 0 16630 1183 16632
rect 0 16600 800 16630
rect 1117 16627 1183 16630
rect 1485 16690 1551 16693
rect 3417 16690 3483 16693
rect 8201 16690 8267 16693
rect 14181 16690 14247 16693
rect 1485 16688 14247 16690
rect 1485 16632 1490 16688
rect 1546 16632 3422 16688
rect 3478 16632 8206 16688
rect 8262 16632 14186 16688
rect 14242 16632 14247 16688
rect 1485 16630 14247 16632
rect 1485 16627 1551 16630
rect 3417 16627 3483 16630
rect 8201 16627 8267 16630
rect 14181 16627 14247 16630
rect 14549 16690 14615 16693
rect 22050 16690 22110 17038
rect 28533 17035 28599 17038
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 22502 16764 22508 16828
rect 22572 16826 22578 16828
rect 22645 16826 22711 16829
rect 22572 16824 22711 16826
rect 22572 16768 22650 16824
rect 22706 16768 22711 16824
rect 22572 16766 22711 16768
rect 22572 16764 22578 16766
rect 22645 16763 22711 16766
rect 23841 16690 23907 16693
rect 14549 16688 22110 16690
rect 14549 16632 14554 16688
rect 14610 16632 22110 16688
rect 14549 16630 22110 16632
rect 22188 16688 23907 16690
rect 22188 16632 23846 16688
rect 23902 16632 23907 16688
rect 22188 16630 23907 16632
rect 14549 16627 14615 16630
rect 2773 16554 2839 16557
rect 6453 16554 6519 16557
rect 8201 16554 8267 16557
rect 2773 16552 8267 16554
rect 2773 16496 2778 16552
rect 2834 16496 6458 16552
rect 6514 16496 8206 16552
rect 8262 16496 8267 16552
rect 2773 16494 8267 16496
rect 2773 16491 2839 16494
rect 6453 16491 6519 16494
rect 8201 16491 8267 16494
rect 9673 16554 9739 16557
rect 19333 16554 19399 16557
rect 9673 16552 19399 16554
rect 9673 16496 9678 16552
rect 9734 16496 19338 16552
rect 19394 16496 19399 16552
rect 9673 16494 19399 16496
rect 9673 16491 9739 16494
rect 19333 16491 19399 16494
rect 13169 16418 13235 16421
rect 16573 16418 16639 16421
rect 13169 16416 16639 16418
rect 13169 16360 13174 16416
rect 13230 16360 16578 16416
rect 16634 16360 16639 16416
rect 13169 16358 16639 16360
rect 13169 16355 13235 16358
rect 16573 16355 16639 16358
rect 21909 16418 21975 16421
rect 22188 16418 22248 16630
rect 23841 16627 23907 16630
rect 28257 16690 28323 16693
rect 31017 16690 31083 16693
rect 28257 16688 31083 16690
rect 28257 16632 28262 16688
rect 28318 16632 31022 16688
rect 31078 16632 31083 16688
rect 28257 16630 31083 16632
rect 28257 16627 28323 16630
rect 31017 16627 31083 16630
rect 21909 16416 22248 16418
rect 21909 16360 21914 16416
rect 21970 16360 22248 16416
rect 21909 16358 22248 16360
rect 21909 16355 21975 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1209 16282 1275 16285
rect 0 16280 1275 16282
rect 0 16224 1214 16280
rect 1270 16224 1275 16280
rect 0 16222 1275 16224
rect 0 16192 800 16222
rect 1209 16219 1275 16222
rect 3785 16282 3851 16285
rect 3785 16280 7850 16282
rect 3785 16224 3790 16280
rect 3846 16224 7850 16280
rect 3785 16222 7850 16224
rect 3785 16219 3851 16222
rect 7281 16146 7347 16149
rect 7557 16146 7623 16149
rect 7281 16144 7623 16146
rect 7281 16088 7286 16144
rect 7342 16088 7562 16144
rect 7618 16088 7623 16144
rect 7281 16086 7623 16088
rect 7790 16146 7850 16222
rect 9622 16220 9628 16284
rect 9692 16282 9698 16284
rect 10593 16282 10659 16285
rect 17125 16284 17191 16285
rect 17125 16282 17172 16284
rect 9692 16280 10659 16282
rect 9692 16224 10598 16280
rect 10654 16224 10659 16280
rect 9692 16222 10659 16224
rect 17080 16280 17172 16282
rect 17080 16224 17130 16280
rect 17080 16222 17172 16224
rect 9692 16220 9698 16222
rect 10593 16219 10659 16222
rect 17125 16220 17172 16222
rect 17236 16220 17242 16284
rect 17125 16219 17191 16220
rect 9489 16146 9555 16149
rect 7790 16144 9555 16146
rect 7790 16088 9494 16144
rect 9550 16088 9555 16144
rect 7790 16086 9555 16088
rect 7281 16083 7347 16086
rect 7557 16083 7623 16086
rect 9489 16083 9555 16086
rect 9622 16084 9628 16148
rect 9692 16146 9698 16148
rect 10542 16146 10548 16148
rect 9692 16086 10548 16146
rect 9692 16084 9698 16086
rect 10542 16084 10548 16086
rect 10612 16146 10618 16148
rect 19885 16146 19951 16149
rect 10612 16144 19951 16146
rect 10612 16088 19890 16144
rect 19946 16088 19951 16144
rect 10612 16086 19951 16088
rect 10612 16084 10618 16086
rect 19885 16083 19951 16086
rect 7557 16010 7623 16013
rect 8109 16010 8175 16013
rect 7557 16008 8175 16010
rect 7557 15952 7562 16008
rect 7618 15952 8114 16008
rect 8170 15952 8175 16008
rect 7557 15950 8175 15952
rect 7557 15947 7623 15950
rect 8109 15947 8175 15950
rect 10961 16010 11027 16013
rect 29545 16010 29611 16013
rect 10961 16008 29611 16010
rect 10961 15952 10966 16008
rect 11022 15952 29550 16008
rect 29606 15952 29611 16008
rect 10961 15950 29611 15952
rect 10961 15947 11027 15950
rect 29545 15947 29611 15950
rect 0 15874 800 15904
rect 1117 15874 1183 15877
rect 0 15872 1183 15874
rect 0 15816 1122 15872
rect 1178 15816 1183 15872
rect 0 15814 1183 15816
rect 0 15784 800 15814
rect 1117 15811 1183 15814
rect 3918 15812 3924 15876
rect 3988 15874 3994 15876
rect 11329 15874 11395 15877
rect 3988 15872 11395 15874
rect 3988 15816 11334 15872
rect 11390 15816 11395 15872
rect 3988 15814 11395 15816
rect 3988 15812 3994 15814
rect 11329 15811 11395 15814
rect 13905 15874 13971 15877
rect 21265 15874 21331 15877
rect 13905 15872 21331 15874
rect 13905 15816 13910 15872
rect 13966 15816 21270 15872
rect 21326 15816 21331 15872
rect 13905 15814 21331 15816
rect 13905 15811 13971 15814
rect 21265 15811 21331 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 7649 15738 7715 15741
rect 12617 15738 12683 15741
rect 7649 15736 12683 15738
rect 7649 15680 7654 15736
rect 7710 15680 12622 15736
rect 12678 15680 12683 15736
rect 7649 15678 12683 15680
rect 7649 15675 7715 15678
rect 12617 15675 12683 15678
rect 13721 15738 13787 15741
rect 20897 15738 20963 15741
rect 13721 15736 20963 15738
rect 13721 15680 13726 15736
rect 13782 15680 20902 15736
rect 20958 15680 20963 15736
rect 13721 15678 20963 15680
rect 13721 15675 13787 15678
rect 20897 15675 20963 15678
rect 12065 15602 12131 15605
rect 29913 15602 29979 15605
rect 12065 15600 29979 15602
rect 12065 15544 12070 15600
rect 12126 15544 29918 15600
rect 29974 15544 29979 15600
rect 12065 15542 29979 15544
rect 12065 15539 12131 15542
rect 29913 15539 29979 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 4061 15466 4127 15469
rect 7097 15466 7163 15469
rect 4061 15464 7163 15466
rect 4061 15408 4066 15464
rect 4122 15408 7102 15464
rect 7158 15408 7163 15464
rect 4061 15406 7163 15408
rect 4061 15403 4127 15406
rect 7097 15403 7163 15406
rect 7373 15466 7439 15469
rect 9213 15466 9279 15469
rect 31937 15466 32003 15469
rect 7373 15464 32003 15466
rect 7373 15408 7378 15464
rect 7434 15408 9218 15464
rect 9274 15408 31942 15464
rect 31998 15408 32003 15464
rect 7373 15406 32003 15408
rect 7373 15403 7439 15406
rect 9213 15403 9279 15406
rect 31937 15403 32003 15406
rect 10961 15330 11027 15333
rect 15469 15330 15535 15333
rect 10961 15328 15535 15330
rect 10961 15272 10966 15328
rect 11022 15272 15474 15328
rect 15530 15272 15535 15328
rect 10961 15270 15535 15272
rect 10961 15267 11027 15270
rect 15469 15267 15535 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 8334 15132 8340 15196
rect 8404 15194 8410 15196
rect 11145 15194 11211 15197
rect 8404 15192 11211 15194
rect 8404 15136 11150 15192
rect 11206 15136 11211 15192
rect 8404 15134 11211 15136
rect 8404 15132 8410 15134
rect 11145 15131 11211 15134
rect 11881 15194 11947 15197
rect 16757 15194 16823 15197
rect 11881 15192 16823 15194
rect 11881 15136 11886 15192
rect 11942 15136 16762 15192
rect 16818 15136 16823 15192
rect 11881 15134 16823 15136
rect 11881 15131 11947 15134
rect 16757 15131 16823 15134
rect 18597 15194 18663 15197
rect 20345 15194 20411 15197
rect 25589 15194 25655 15197
rect 18597 15192 25655 15194
rect 18597 15136 18602 15192
rect 18658 15136 20350 15192
rect 20406 15136 25594 15192
rect 25650 15136 25655 15192
rect 18597 15134 25655 15136
rect 18597 15131 18663 15134
rect 20345 15131 20411 15134
rect 25589 15131 25655 15134
rect 0 15058 800 15088
rect 1117 15058 1183 15061
rect 0 15056 1183 15058
rect 0 15000 1122 15056
rect 1178 15000 1183 15056
rect 0 14998 1183 15000
rect 0 14968 800 14998
rect 1117 14995 1183 14998
rect 9254 14996 9260 15060
rect 9324 15058 9330 15060
rect 9397 15058 9463 15061
rect 9324 15056 9463 15058
rect 9324 15000 9402 15056
rect 9458 15000 9463 15056
rect 9324 14998 9463 15000
rect 9324 14996 9330 14998
rect 9397 14995 9463 14998
rect 9673 15058 9739 15061
rect 10961 15058 11027 15061
rect 9673 15056 11027 15058
rect 9673 15000 9678 15056
rect 9734 15000 10966 15056
rect 11022 15000 11027 15056
rect 9673 14998 11027 15000
rect 9673 14995 9739 14998
rect 10961 14995 11027 14998
rect 11973 15058 12039 15061
rect 33317 15058 33383 15061
rect 11973 15056 33383 15058
rect 11973 15000 11978 15056
rect 12034 15000 33322 15056
rect 33378 15000 33383 15056
rect 11973 14998 33383 15000
rect 11973 14995 12039 14998
rect 33317 14995 33383 14998
rect 7833 14922 7899 14925
rect 10961 14922 11027 14925
rect 7833 14920 11027 14922
rect 7833 14864 7838 14920
rect 7894 14864 10966 14920
rect 11022 14864 11027 14920
rect 7833 14862 11027 14864
rect 7833 14859 7899 14862
rect 10961 14859 11027 14862
rect 12065 14922 12131 14925
rect 13537 14922 13603 14925
rect 12065 14920 13603 14922
rect 12065 14864 12070 14920
rect 12126 14864 13542 14920
rect 13598 14864 13603 14920
rect 12065 14862 13603 14864
rect 12065 14859 12131 14862
rect 13537 14859 13603 14862
rect 17125 14922 17191 14925
rect 19333 14922 19399 14925
rect 17125 14920 19399 14922
rect 17125 14864 17130 14920
rect 17186 14864 19338 14920
rect 19394 14864 19399 14920
rect 17125 14862 19399 14864
rect 17125 14859 17191 14862
rect 19333 14859 19399 14862
rect 20161 14922 20227 14925
rect 25129 14922 25195 14925
rect 20161 14920 25195 14922
rect 20161 14864 20166 14920
rect 20222 14864 25134 14920
rect 25190 14864 25195 14920
rect 20161 14862 25195 14864
rect 20161 14859 20227 14862
rect 25129 14859 25195 14862
rect 6637 14786 6703 14789
rect 9489 14786 9555 14789
rect 6637 14784 9555 14786
rect 6637 14728 6642 14784
rect 6698 14728 9494 14784
rect 9550 14728 9555 14784
rect 6637 14726 9555 14728
rect 6637 14723 6703 14726
rect 9489 14723 9555 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 5441 14650 5507 14653
rect 11053 14650 11119 14653
rect 5441 14648 11119 14650
rect 5441 14592 5446 14648
rect 5502 14592 11058 14648
rect 11114 14592 11119 14648
rect 5441 14590 11119 14592
rect 5441 14587 5507 14590
rect 11053 14587 11119 14590
rect 5165 14514 5231 14517
rect 8569 14514 8635 14517
rect 5165 14512 8635 14514
rect 5165 14456 5170 14512
rect 5226 14456 8574 14512
rect 8630 14456 8635 14512
rect 5165 14454 8635 14456
rect 5165 14451 5231 14454
rect 8569 14451 8635 14454
rect 11053 14514 11119 14517
rect 15653 14514 15719 14517
rect 11053 14512 15719 14514
rect 11053 14456 11058 14512
rect 11114 14456 15658 14512
rect 15714 14456 15719 14512
rect 11053 14454 15719 14456
rect 11053 14451 11119 14454
rect 15653 14451 15719 14454
rect 7649 14380 7715 14381
rect 7598 14378 7604 14380
rect 7558 14318 7604 14378
rect 7668 14376 7715 14380
rect 7710 14320 7715 14376
rect 7598 14316 7604 14318
rect 7668 14316 7715 14320
rect 7649 14315 7715 14316
rect 9765 14378 9831 14381
rect 10501 14378 10567 14381
rect 10961 14378 11027 14381
rect 9765 14376 11027 14378
rect 9765 14320 9770 14376
rect 9826 14320 10506 14376
rect 10562 14320 10966 14376
rect 11022 14320 11027 14376
rect 9765 14318 11027 14320
rect 9765 14315 9831 14318
rect 10501 14315 10567 14318
rect 10961 14315 11027 14318
rect 15653 14378 15719 14381
rect 21357 14378 21423 14381
rect 15653 14376 21423 14378
rect 15653 14320 15658 14376
rect 15714 14320 21362 14376
rect 21418 14320 21423 14376
rect 15653 14318 21423 14320
rect 15653 14315 15719 14318
rect 21357 14315 21423 14318
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 4521 14106 4587 14109
rect 5717 14106 5783 14109
rect 4521 14104 5783 14106
rect 4521 14048 4526 14104
rect 4582 14048 5722 14104
rect 5778 14048 5783 14104
rect 4521 14046 5783 14048
rect 4521 14043 4587 14046
rect 5717 14043 5783 14046
rect 1853 13972 1919 13973
rect 1853 13970 1900 13972
rect 1812 13968 1900 13970
rect 1964 13970 1970 13972
rect 19517 13970 19583 13973
rect 1964 13968 19583 13970
rect 1812 13912 1858 13968
rect 1964 13912 19522 13968
rect 19578 13912 19583 13968
rect 1812 13910 1900 13912
rect 1853 13908 1900 13910
rect 1964 13910 19583 13912
rect 1964 13908 1970 13910
rect 1853 13907 1919 13908
rect 19517 13907 19583 13910
rect 22369 13970 22435 13973
rect 22502 13970 22508 13972
rect 22369 13968 22508 13970
rect 22369 13912 22374 13968
rect 22430 13912 22508 13968
rect 22369 13910 22508 13912
rect 22369 13907 22435 13910
rect 22502 13908 22508 13910
rect 22572 13908 22578 13972
rect 22645 13970 22711 13973
rect 23841 13970 23907 13973
rect 22645 13968 23907 13970
rect 22645 13912 22650 13968
rect 22706 13912 23846 13968
rect 23902 13912 23907 13968
rect 22645 13910 23907 13912
rect 22645 13907 22711 13910
rect 23841 13907 23907 13910
rect 0 13834 800 13864
rect 2037 13834 2103 13837
rect 0 13832 2103 13834
rect 0 13776 2042 13832
rect 2098 13776 2103 13832
rect 0 13774 2103 13776
rect 0 13744 800 13774
rect 2037 13771 2103 13774
rect 9765 13834 9831 13837
rect 10041 13834 10107 13837
rect 10777 13834 10843 13837
rect 9765 13832 9874 13834
rect 9765 13776 9770 13832
rect 9826 13776 9874 13832
rect 9765 13771 9874 13776
rect 10041 13832 10843 13834
rect 10041 13776 10046 13832
rect 10102 13776 10782 13832
rect 10838 13776 10843 13832
rect 10041 13774 10843 13776
rect 10041 13771 10107 13774
rect 10777 13771 10843 13774
rect 3325 13698 3391 13701
rect 4521 13698 4587 13701
rect 3325 13696 4587 13698
rect 3325 13640 3330 13696
rect 3386 13640 4526 13696
rect 4582 13640 4587 13696
rect 3325 13638 4587 13640
rect 3325 13635 3391 13638
rect 4521 13635 4587 13638
rect 6545 13698 6611 13701
rect 9814 13698 9874 13771
rect 11329 13698 11395 13701
rect 6545 13696 11395 13698
rect 6545 13640 6550 13696
rect 6606 13640 11334 13696
rect 11390 13640 11395 13696
rect 6545 13638 11395 13640
rect 6545 13635 6611 13638
rect 11329 13635 11395 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 0 13426 800 13456
rect 1209 13426 1275 13429
rect 0 13424 1275 13426
rect 0 13368 1214 13424
rect 1270 13368 1275 13424
rect 0 13366 1275 13368
rect 0 13336 800 13366
rect 1209 13363 1275 13366
rect 1945 13426 2011 13429
rect 19425 13426 19491 13429
rect 1945 13424 19491 13426
rect 1945 13368 1950 13424
rect 2006 13368 19430 13424
rect 19486 13368 19491 13424
rect 1945 13366 19491 13368
rect 1945 13363 2011 13366
rect 19425 13363 19491 13366
rect 3877 13290 3943 13293
rect 5942 13290 5948 13292
rect 3877 13288 5948 13290
rect 3877 13232 3882 13288
rect 3938 13232 5948 13288
rect 3877 13230 5948 13232
rect 3877 13227 3943 13230
rect 5942 13228 5948 13230
rect 6012 13290 6018 13292
rect 6494 13290 6500 13292
rect 6012 13230 6500 13290
rect 6012 13228 6018 13230
rect 6494 13228 6500 13230
rect 6564 13228 6570 13292
rect 9397 13290 9463 13293
rect 26141 13290 26207 13293
rect 9397 13288 26207 13290
rect 9397 13232 9402 13288
rect 9458 13232 26146 13288
rect 26202 13232 26207 13288
rect 9397 13230 26207 13232
rect 9397 13227 9463 13230
rect 26141 13227 26207 13230
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 3877 13018 3943 13021
rect 10685 13018 10751 13021
rect 0 13016 3943 13018
rect 0 12960 3882 13016
rect 3938 12960 3943 13016
rect 0 12958 3943 12960
rect 0 12928 800 12958
rect 3877 12955 3943 12958
rect 9998 13016 10751 13018
rect 9998 12960 10690 13016
rect 10746 12960 10751 13016
rect 9998 12958 10751 12960
rect 7465 12882 7531 12885
rect 8753 12882 8819 12885
rect 7465 12880 8819 12882
rect 7465 12824 7470 12880
rect 7526 12824 8758 12880
rect 8814 12824 8819 12880
rect 7465 12822 8819 12824
rect 7465 12819 7531 12822
rect 8753 12819 8819 12822
rect 4061 12746 4127 12749
rect 2730 12744 4127 12746
rect 2730 12688 4066 12744
rect 4122 12688 4127 12744
rect 2730 12686 4127 12688
rect 0 12610 800 12640
rect 2730 12610 2790 12686
rect 4061 12683 4127 12686
rect 9998 12613 10058 12958
rect 10685 12955 10751 12958
rect 10685 12882 10751 12885
rect 22277 12882 22343 12885
rect 10685 12880 22343 12882
rect 10685 12824 10690 12880
rect 10746 12824 22282 12880
rect 22338 12824 22343 12880
rect 10685 12822 22343 12824
rect 10685 12819 10751 12822
rect 22277 12819 22343 12822
rect 13169 12746 13235 12749
rect 16573 12746 16639 12749
rect 13169 12744 16639 12746
rect 13169 12688 13174 12744
rect 13230 12688 16578 12744
rect 16634 12688 16639 12744
rect 13169 12686 16639 12688
rect 13169 12683 13235 12686
rect 16573 12683 16639 12686
rect 0 12550 2790 12610
rect 4153 12610 4219 12613
rect 4429 12610 4495 12613
rect 4153 12608 4495 12610
rect 4153 12552 4158 12608
rect 4214 12552 4434 12608
rect 4490 12552 4495 12608
rect 4153 12550 4495 12552
rect 0 12520 800 12550
rect 4153 12547 4219 12550
rect 4429 12547 4495 12550
rect 9949 12608 10058 12613
rect 9949 12552 9954 12608
rect 10010 12552 10058 12608
rect 9949 12550 10058 12552
rect 9949 12547 10015 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 4153 12338 4219 12341
rect 4286 12338 4292 12340
rect 4153 12336 4292 12338
rect 4153 12280 4158 12336
rect 4214 12280 4292 12336
rect 4153 12278 4292 12280
rect 4153 12275 4219 12278
rect 4286 12276 4292 12278
rect 4356 12276 4362 12340
rect 6729 12338 6795 12341
rect 15193 12338 15259 12341
rect 20253 12338 20319 12341
rect 6729 12336 12450 12338
rect 6729 12280 6734 12336
rect 6790 12280 12450 12336
rect 6729 12278 12450 12280
rect 6729 12275 6795 12278
rect 0 12202 800 12232
rect 933 12202 999 12205
rect 0 12200 999 12202
rect 0 12144 938 12200
rect 994 12144 999 12200
rect 0 12142 999 12144
rect 0 12112 800 12142
rect 933 12139 999 12142
rect 3509 12202 3575 12205
rect 9622 12202 9628 12204
rect 3509 12200 9628 12202
rect 3509 12144 3514 12200
rect 3570 12144 9628 12200
rect 3509 12142 9628 12144
rect 3509 12139 3575 12142
rect 9622 12140 9628 12142
rect 9692 12140 9698 12204
rect 12390 12202 12450 12278
rect 15193 12336 20319 12338
rect 15193 12280 15198 12336
rect 15254 12280 20258 12336
rect 20314 12280 20319 12336
rect 15193 12278 20319 12280
rect 15193 12275 15259 12278
rect 20253 12275 20319 12278
rect 27705 12202 27771 12205
rect 12390 12200 27771 12202
rect 12390 12144 27710 12200
rect 27766 12144 27771 12200
rect 12390 12142 27771 12144
rect 27705 12139 27771 12142
rect 13261 12066 13327 12069
rect 16205 12066 16271 12069
rect 13261 12064 16271 12066
rect 13261 12008 13266 12064
rect 13322 12008 16210 12064
rect 16266 12008 16271 12064
rect 13261 12006 16271 12008
rect 13261 12003 13327 12006
rect 16205 12003 16271 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 1761 11930 1827 11933
rect 1894 11930 1900 11932
rect 1761 11928 1900 11930
rect 1761 11872 1766 11928
rect 1822 11872 1900 11928
rect 1761 11870 1900 11872
rect 1761 11867 1827 11870
rect 1894 11868 1900 11870
rect 1964 11868 1970 11932
rect 13169 11930 13235 11933
rect 14365 11930 14431 11933
rect 13169 11928 14431 11930
rect 13169 11872 13174 11928
rect 13230 11872 14370 11928
rect 14426 11872 14431 11928
rect 13169 11870 14431 11872
rect 13169 11867 13235 11870
rect 14365 11867 14431 11870
rect 0 11794 800 11824
rect 6453 11794 6519 11797
rect 9305 11794 9371 11797
rect 0 11734 1594 11794
rect 0 11704 800 11734
rect 1534 11658 1594 11734
rect 6453 11792 9371 11794
rect 6453 11736 6458 11792
rect 6514 11736 9310 11792
rect 9366 11736 9371 11792
rect 6453 11734 9371 11736
rect 6453 11731 6519 11734
rect 9305 11731 9371 11734
rect 14273 11794 14339 11797
rect 17401 11794 17467 11797
rect 14273 11792 17467 11794
rect 14273 11736 14278 11792
rect 14334 11736 17406 11792
rect 17462 11736 17467 11792
rect 14273 11734 17467 11736
rect 14273 11731 14339 11734
rect 17401 11731 17467 11734
rect 1669 11658 1735 11661
rect 1534 11656 1735 11658
rect 1534 11600 1674 11656
rect 1730 11600 1735 11656
rect 1534 11598 1735 11600
rect 1669 11595 1735 11598
rect 3509 11658 3575 11661
rect 3734 11658 3740 11660
rect 3509 11656 3740 11658
rect 3509 11600 3514 11656
rect 3570 11600 3740 11656
rect 3509 11598 3740 11600
rect 3509 11595 3575 11598
rect 3734 11596 3740 11598
rect 3804 11658 3810 11660
rect 11145 11658 11211 11661
rect 3804 11656 11211 11658
rect 3804 11600 11150 11656
rect 11206 11600 11211 11656
rect 3804 11598 11211 11600
rect 3804 11596 3810 11598
rect 11145 11595 11211 11598
rect 3785 11522 3851 11525
rect 3785 11520 12450 11522
rect 3785 11464 3790 11520
rect 3846 11464 12450 11520
rect 3785 11462 12450 11464
rect 3785 11459 3851 11462
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 7281 11386 7347 11389
rect 7414 11386 7420 11388
rect 0 11326 2790 11386
rect 0 11296 800 11326
rect 2730 11250 2790 11326
rect 7281 11384 7420 11386
rect 7281 11328 7286 11384
rect 7342 11328 7420 11384
rect 7281 11326 7420 11328
rect 7281 11323 7347 11326
rect 7414 11324 7420 11326
rect 7484 11324 7490 11388
rect 3693 11250 3759 11253
rect 2730 11248 3759 11250
rect 2730 11192 3698 11248
rect 3754 11192 3759 11248
rect 2730 11190 3759 11192
rect 3693 11187 3759 11190
rect 6177 11250 6243 11253
rect 7230 11250 7236 11252
rect 6177 11248 7236 11250
rect 6177 11192 6182 11248
rect 6238 11192 7236 11248
rect 6177 11190 7236 11192
rect 6177 11187 6243 11190
rect 7230 11188 7236 11190
rect 7300 11188 7306 11252
rect 12390 11250 12450 11462
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 20621 11250 20687 11253
rect 12390 11248 20687 11250
rect 12390 11192 20626 11248
rect 20682 11192 20687 11248
rect 12390 11190 20687 11192
rect 20621 11187 20687 11190
rect 2589 11114 2655 11117
rect 3366 11114 3372 11116
rect 2589 11112 3372 11114
rect 2589 11056 2594 11112
rect 2650 11056 3372 11112
rect 2589 11054 3372 11056
rect 2589 11051 2655 11054
rect 3366 11052 3372 11054
rect 3436 11114 3442 11116
rect 3785 11114 3851 11117
rect 3436 11112 3851 11114
rect 3436 11056 3790 11112
rect 3846 11056 3851 11112
rect 3436 11054 3851 11056
rect 3436 11052 3442 11054
rect 3785 11051 3851 11054
rect 3918 11052 3924 11116
rect 3988 11114 3994 11116
rect 5441 11114 5507 11117
rect 3988 11112 5507 11114
rect 3988 11056 5446 11112
rect 5502 11056 5507 11112
rect 3988 11054 5507 11056
rect 3988 11052 3994 11054
rect 5441 11051 5507 11054
rect 5901 11114 5967 11117
rect 6310 11114 6316 11116
rect 5901 11112 6316 11114
rect 5901 11056 5906 11112
rect 5962 11056 6316 11112
rect 5901 11054 6316 11056
rect 5901 11051 5967 11054
rect 6310 11052 6316 11054
rect 6380 11052 6386 11116
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 5349 10980 5415 10981
rect 5349 10976 5396 10980
rect 5460 10978 5466 10980
rect 5349 10920 5354 10976
rect 5349 10916 5396 10920
rect 5460 10918 5506 10978
rect 5460 10916 5466 10918
rect 5349 10915 5415 10916
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 5206 10780 5212 10844
rect 5276 10842 5282 10844
rect 5625 10842 5691 10845
rect 5276 10840 5691 10842
rect 5276 10784 5630 10840
rect 5686 10784 5691 10840
rect 5276 10782 5691 10784
rect 5276 10780 5282 10782
rect 5625 10779 5691 10782
rect 7005 10706 7071 10709
rect 22134 10706 22140 10708
rect 7005 10704 22140 10706
rect 7005 10648 7010 10704
rect 7066 10648 22140 10704
rect 7005 10646 22140 10648
rect 7005 10643 7071 10646
rect 22134 10644 22140 10646
rect 22204 10644 22210 10708
rect 0 10570 800 10600
rect 2773 10570 2839 10573
rect 0 10568 2839 10570
rect 0 10512 2778 10568
rect 2834 10512 2839 10568
rect 0 10510 2839 10512
rect 0 10480 800 10510
rect 2773 10507 2839 10510
rect 4337 10434 4403 10437
rect 11513 10434 11579 10437
rect 11881 10434 11947 10437
rect 4337 10432 11947 10434
rect 4337 10376 4342 10432
rect 4398 10376 11518 10432
rect 11574 10376 11886 10432
rect 11942 10376 11947 10432
rect 4337 10374 11947 10376
rect 4337 10371 4403 10374
rect 11513 10371 11579 10374
rect 11881 10371 11947 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 13721 10298 13787 10301
rect 22686 10298 22692 10300
rect 13721 10296 22692 10298
rect 13721 10240 13726 10296
rect 13782 10240 22692 10296
rect 13721 10238 22692 10240
rect 13721 10235 13787 10238
rect 22686 10236 22692 10238
rect 22756 10236 22762 10300
rect 0 10162 800 10192
rect 2865 10162 2931 10165
rect 0 10160 2931 10162
rect 0 10104 2870 10160
rect 2926 10104 2931 10160
rect 0 10102 2931 10104
rect 0 10072 800 10102
rect 2865 10099 2931 10102
rect 6913 10162 6979 10165
rect 13854 10162 13860 10164
rect 6913 10160 13860 10162
rect 6913 10104 6918 10160
rect 6974 10104 13860 10160
rect 6913 10102 13860 10104
rect 6913 10099 6979 10102
rect 13854 10100 13860 10102
rect 13924 10100 13930 10164
rect 3417 10026 3483 10029
rect 4061 10026 4127 10029
rect 14641 10026 14707 10029
rect 3417 10024 14707 10026
rect 3417 9968 3422 10024
rect 3478 9968 4066 10024
rect 4122 9968 14646 10024
rect 14702 9968 14707 10024
rect 3417 9966 14707 9968
rect 3417 9963 3483 9966
rect 4061 9963 4127 9966
rect 14641 9963 14707 9966
rect 5625 9890 5691 9893
rect 5758 9890 5764 9892
rect 5625 9888 5764 9890
rect 5625 9832 5630 9888
rect 5686 9832 5764 9888
rect 5625 9830 5764 9832
rect 5625 9827 5691 9830
rect 5758 9828 5764 9830
rect 5828 9828 5834 9892
rect 11513 9890 11579 9893
rect 15653 9890 15719 9893
rect 11513 9888 15719 9890
rect 11513 9832 11518 9888
rect 11574 9832 15658 9888
rect 15714 9832 15719 9888
rect 11513 9830 15719 9832
rect 11513 9827 11579 9830
rect 15653 9827 15719 9830
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1577 9754 1643 9757
rect 0 9752 1643 9754
rect 0 9696 1582 9752
rect 1638 9696 1643 9752
rect 0 9694 1643 9696
rect 0 9664 800 9694
rect 1577 9691 1643 9694
rect 3233 9618 3299 9621
rect 5533 9620 5599 9621
rect 3366 9618 3372 9620
rect 3233 9616 3372 9618
rect 3233 9560 3238 9616
rect 3294 9560 3372 9616
rect 3233 9558 3372 9560
rect 3233 9555 3299 9558
rect 3366 9556 3372 9558
rect 3436 9556 3442 9620
rect 5533 9616 5580 9620
rect 5644 9618 5650 9620
rect 5533 9560 5538 9616
rect 5533 9556 5580 9560
rect 5644 9558 5690 9618
rect 5644 9556 5650 9558
rect 5533 9555 5599 9556
rect 2262 9420 2268 9484
rect 2332 9482 2338 9484
rect 3601 9482 3667 9485
rect 2332 9480 3667 9482
rect 2332 9424 3606 9480
rect 3662 9424 3667 9480
rect 2332 9422 3667 9424
rect 2332 9420 2338 9422
rect 3601 9419 3667 9422
rect 3785 9482 3851 9485
rect 13721 9482 13787 9485
rect 3785 9480 13787 9482
rect 3785 9424 3790 9480
rect 3846 9424 13726 9480
rect 13782 9424 13787 9480
rect 3785 9422 13787 9424
rect 3785 9419 3851 9422
rect 13721 9419 13787 9422
rect 0 9346 800 9376
rect 2773 9346 2839 9349
rect 0 9344 2839 9346
rect 0 9288 2778 9344
rect 2834 9288 2839 9344
rect 0 9286 2839 9288
rect 0 9256 800 9286
rect 2773 9283 2839 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 7189 9210 7255 9213
rect 8334 9210 8340 9212
rect 7189 9208 8340 9210
rect 7189 9152 7194 9208
rect 7250 9152 8340 9208
rect 7189 9150 8340 9152
rect 7189 9147 7255 9150
rect 8334 9148 8340 9150
rect 8404 9148 8410 9212
rect 7741 9074 7807 9077
rect 24117 9074 24183 9077
rect 7741 9072 24183 9074
rect 7741 9016 7746 9072
rect 7802 9016 24122 9072
rect 24178 9016 24183 9072
rect 7741 9014 24183 9016
rect 7741 9011 7807 9014
rect 24117 9011 24183 9014
rect 0 8938 800 8968
rect 1761 8938 1827 8941
rect 0 8936 1827 8938
rect 0 8880 1766 8936
rect 1822 8880 1827 8936
rect 0 8878 1827 8880
rect 0 8848 800 8878
rect 1761 8875 1827 8878
rect 6637 8938 6703 8941
rect 9806 8938 9812 8940
rect 6637 8936 9812 8938
rect 6637 8880 6642 8936
rect 6698 8880 9812 8936
rect 6637 8878 9812 8880
rect 6637 8875 6703 8878
rect 9806 8876 9812 8878
rect 9876 8876 9882 8940
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 6453 8668 6519 8669
rect 6453 8666 6500 8668
rect 6408 8664 6500 8666
rect 6408 8608 6458 8664
rect 6408 8606 6500 8608
rect 6453 8604 6500 8606
rect 6564 8604 6570 8668
rect 6453 8603 6519 8604
rect 0 8530 800 8560
rect 2865 8530 2931 8533
rect 0 8528 2931 8530
rect 0 8472 2870 8528
rect 2926 8472 2931 8528
rect 0 8470 2931 8472
rect 0 8440 800 8470
rect 2865 8467 2931 8470
rect 9857 8394 9923 8397
rect 32857 8394 32923 8397
rect 9857 8392 32923 8394
rect 9857 8336 9862 8392
rect 9918 8336 32862 8392
rect 32918 8336 32923 8392
rect 9857 8334 32923 8336
rect 9857 8331 9923 8334
rect 32857 8331 32923 8334
rect 9305 8258 9371 8261
rect 9438 8258 9444 8260
rect 9305 8256 9444 8258
rect 9305 8200 9310 8256
rect 9366 8200 9444 8256
rect 9305 8198 9444 8200
rect 9305 8195 9371 8198
rect 9438 8196 9444 8198
rect 9508 8196 9514 8260
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 2773 8122 2839 8125
rect 0 8120 2839 8122
rect 0 8064 2778 8120
rect 2834 8064 2839 8120
rect 0 8062 2839 8064
rect 0 8032 800 8062
rect 2773 8059 2839 8062
rect 3325 7850 3391 7853
rect 3877 7850 3943 7853
rect 3325 7848 3943 7850
rect 3325 7792 3330 7848
rect 3386 7792 3882 7848
rect 3938 7792 3943 7848
rect 3325 7790 3943 7792
rect 3325 7787 3391 7790
rect 3877 7787 3943 7790
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 0 7306 800 7336
rect 2865 7306 2931 7309
rect 0 7304 2931 7306
rect 0 7248 2870 7304
rect 2926 7248 2931 7304
rect 0 7246 2931 7248
rect 0 7216 800 7246
rect 2865 7243 2931 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 3325 6898 3391 6901
rect 0 6896 3391 6898
rect 0 6840 3330 6896
rect 3386 6840 3391 6896
rect 0 6838 3391 6840
rect 0 6808 800 6838
rect 3325 6835 3391 6838
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 0 4450 800 4480
rect 1761 4450 1827 4453
rect 0 4448 1827 4450
rect 0 4392 1766 4448
rect 1822 4392 1827 4448
rect 0 4390 1827 4392
rect 0 4360 800 4390
rect 1761 4387 1827 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4042 800 4072
rect 1301 4042 1367 4045
rect 0 4040 1367 4042
rect 0 3984 1306 4040
rect 1362 3984 1367 4040
rect 0 3982 1367 3984
rect 0 3952 800 3982
rect 1301 3979 1367 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1209 3634 1275 3637
rect 0 3632 1275 3634
rect 0 3576 1214 3632
rect 1270 3576 1275 3632
rect 0 3574 1275 3576
rect 0 3544 800 3574
rect 1209 3571 1275 3574
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 0 2410 800 2440
rect 1209 2410 1275 2413
rect 0 2408 1275 2410
rect 0 2352 1214 2408
rect 1270 2352 1275 2408
rect 0 2350 1275 2352
rect 0 2320 800 2350
rect 1209 2347 1275 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1301 2002 1367 2005
rect 0 2000 1367 2002
rect 0 1944 1306 2000
rect 1362 1944 1367 2000
rect 0 1942 1367 1944
rect 0 1912 800 1942
rect 1301 1939 1367 1942
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
<< via3 >>
rect 11652 24924 11716 24988
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 9812 23700 9876 23764
rect 2268 23428 2332 23492
rect 4292 23428 4356 23492
rect 22140 23488 22204 23492
rect 22140 23432 22190 23488
rect 22190 23432 22204 23488
rect 22140 23428 22204 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 5580 23156 5644 23220
rect 7420 23020 7484 23084
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 5396 22612 5460 22676
rect 7236 22672 7300 22676
rect 7236 22616 7250 22672
rect 7250 22616 7300 22672
rect 7236 22612 7300 22616
rect 17172 22476 17236 22540
rect 3924 22340 3988 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 17172 22204 17236 22268
rect 10548 21796 10612 21860
rect 22692 21796 22756 21860
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 5764 21388 5828 21452
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 3740 20708 3804 20772
rect 6316 20708 6380 20772
rect 9444 20768 9508 20772
rect 9444 20712 9458 20768
rect 9458 20712 9508 20768
rect 9444 20708 9508 20712
rect 13860 20768 13924 20772
rect 13860 20712 13910 20768
rect 13910 20712 13924 20768
rect 13860 20708 13924 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 9628 19348 9692 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 9076 18728 9140 18732
rect 9076 18672 9126 18728
rect 9126 18672 9140 18728
rect 9076 18668 9140 18672
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 5212 18048 5276 18052
rect 5212 17992 5262 18048
rect 5262 17992 5276 18048
rect 5212 17988 5276 17992
rect 5948 17988 6012 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 11652 17852 11716 17916
rect 7604 17716 7668 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 9260 17368 9324 17372
rect 9260 17312 9310 17368
rect 9310 17312 9324 17368
rect 9260 17308 9324 17312
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 9076 16764 9140 16828
rect 11652 16824 11716 16828
rect 11652 16768 11702 16824
rect 11702 16768 11716 16824
rect 11652 16764 11716 16768
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 22508 16764 22572 16828
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 9628 16220 9692 16284
rect 17172 16280 17236 16284
rect 17172 16224 17186 16280
rect 17186 16224 17236 16280
rect 17172 16220 17236 16224
rect 9628 16084 9692 16148
rect 10548 16084 10612 16148
rect 3924 15812 3988 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 8340 15132 8404 15196
rect 9260 14996 9324 15060
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7604 14376 7668 14380
rect 7604 14320 7654 14376
rect 7654 14320 7668 14376
rect 7604 14316 7668 14320
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 1900 13968 1964 13972
rect 1900 13912 1914 13968
rect 1914 13912 1964 13968
rect 1900 13908 1964 13912
rect 22508 13908 22572 13972
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 5948 13228 6012 13292
rect 6500 13228 6564 13292
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 4292 12276 4356 12340
rect 9628 12140 9692 12204
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 1900 11868 1964 11932
rect 3740 11596 3804 11660
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 7420 11324 7484 11388
rect 7236 11188 7300 11252
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 3372 11052 3436 11116
rect 3924 11052 3988 11116
rect 6316 11052 6380 11116
rect 5396 10976 5460 10980
rect 5396 10920 5410 10976
rect 5410 10920 5460 10976
rect 5396 10916 5460 10920
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 5212 10780 5276 10844
rect 22140 10644 22204 10708
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 22692 10236 22756 10300
rect 13860 10100 13924 10164
rect 5764 9828 5828 9892
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 3372 9556 3436 9620
rect 5580 9616 5644 9620
rect 5580 9560 5594 9616
rect 5594 9560 5644 9616
rect 5580 9556 5644 9560
rect 2268 9420 2332 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 8340 9148 8404 9212
rect 9812 8876 9876 8940
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 6500 8664 6564 8668
rect 6500 8608 6514 8664
rect 6514 8608 6564 8664
rect 6500 8604 6564 8608
rect 9444 8196 9508 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 11651 24988 11717 24989
rect 11651 24924 11652 24988
rect 11716 24924 11717 24988
rect 11651 24923 11717 24924
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2267 23492 2333 23493
rect 2267 23428 2268 23492
rect 2332 23428 2333 23492
rect 2267 23427 2333 23428
rect 1899 13972 1965 13973
rect 1899 13908 1900 13972
rect 1964 13908 1965 13972
rect 1899 13907 1965 13908
rect 1902 11933 1962 13907
rect 1899 11932 1965 11933
rect 1899 11868 1900 11932
rect 1964 11868 1965 11932
rect 1899 11867 1965 11868
rect 2270 9485 2330 23427
rect 2944 23424 3264 24448
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 4291 23492 4357 23493
rect 4291 23428 4292 23492
rect 4356 23428 4357 23492
rect 4291 23427 4357 23428
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 3923 22404 3989 22405
rect 3923 22340 3924 22404
rect 3988 22340 3989 22404
rect 3923 22339 3989 22340
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 3739 20772 3805 20773
rect 3739 20708 3740 20772
rect 3804 20708 3805 20772
rect 3739 20707 3805 20708
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 3742 11661 3802 20707
rect 3926 15877 3986 22339
rect 3923 15876 3989 15877
rect 3923 15812 3924 15876
rect 3988 15812 3989 15876
rect 3923 15811 3989 15812
rect 3739 11660 3805 11661
rect 3739 11596 3740 11660
rect 3804 11596 3805 11660
rect 3739 11595 3805 11596
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 3926 11117 3986 15811
rect 4294 12341 4354 23427
rect 5579 23220 5645 23221
rect 5579 23156 5580 23220
rect 5644 23156 5645 23220
rect 5579 23155 5645 23156
rect 5395 22676 5461 22677
rect 5395 22612 5396 22676
rect 5460 22612 5461 22676
rect 5395 22611 5461 22612
rect 5211 18052 5277 18053
rect 5211 17988 5212 18052
rect 5276 17988 5277 18052
rect 5211 17987 5277 17988
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 3371 11116 3437 11117
rect 3371 11052 3372 11116
rect 3436 11052 3437 11116
rect 3371 11051 3437 11052
rect 3923 11116 3989 11117
rect 3923 11052 3924 11116
rect 3988 11052 3989 11116
rect 3923 11051 3989 11052
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2267 9484 2333 9485
rect 2267 9420 2268 9484
rect 2332 9420 2333 9484
rect 2267 9419 2333 9420
rect 2944 9280 3264 10304
rect 3374 9621 3434 11051
rect 5214 10845 5274 17987
rect 5398 10981 5458 22611
rect 5395 10980 5461 10981
rect 5395 10916 5396 10980
rect 5460 10916 5461 10980
rect 5395 10915 5461 10916
rect 5211 10844 5277 10845
rect 5211 10780 5212 10844
rect 5276 10780 5277 10844
rect 5211 10779 5277 10780
rect 5582 9621 5642 23155
rect 7419 23084 7485 23085
rect 7419 23020 7420 23084
rect 7484 23020 7485 23084
rect 7419 23019 7485 23020
rect 7235 22676 7301 22677
rect 7235 22612 7236 22676
rect 7300 22612 7301 22676
rect 7235 22611 7301 22612
rect 5763 21452 5829 21453
rect 5763 21388 5764 21452
rect 5828 21388 5829 21452
rect 5763 21387 5829 21388
rect 5766 9893 5826 21387
rect 6315 20772 6381 20773
rect 6315 20708 6316 20772
rect 6380 20708 6381 20772
rect 6315 20707 6381 20708
rect 5947 18052 6013 18053
rect 5947 17988 5948 18052
rect 6012 17988 6013 18052
rect 5947 17987 6013 17988
rect 5950 13293 6010 17987
rect 5947 13292 6013 13293
rect 5947 13228 5948 13292
rect 6012 13228 6013 13292
rect 5947 13227 6013 13228
rect 6318 11117 6378 20707
rect 6499 13292 6565 13293
rect 6499 13228 6500 13292
rect 6564 13228 6565 13292
rect 6499 13227 6565 13228
rect 6315 11116 6381 11117
rect 6315 11052 6316 11116
rect 6380 11052 6381 11116
rect 6315 11051 6381 11052
rect 5763 9892 5829 9893
rect 5763 9828 5764 9892
rect 5828 9828 5829 9892
rect 5763 9827 5829 9828
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 5579 9620 5645 9621
rect 5579 9556 5580 9620
rect 5644 9556 5645 9620
rect 5579 9555 5645 9556
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 6502 8669 6562 13227
rect 7238 11253 7298 22611
rect 7422 11389 7482 23019
rect 7944 22880 8264 23904
rect 9811 23764 9877 23765
rect 9811 23700 9812 23764
rect 9876 23700 9877 23764
rect 9811 23699 9877 23700
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 9443 20772 9509 20773
rect 9443 20708 9444 20772
rect 9508 20708 9509 20772
rect 9443 20707 9509 20708
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 9075 18732 9141 18733
rect 9075 18668 9076 18732
rect 9140 18668 9141 18732
rect 9075 18667 9141 18668
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7603 17780 7669 17781
rect 7603 17716 7604 17780
rect 7668 17716 7669 17780
rect 7603 17715 7669 17716
rect 7606 14381 7666 17715
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 9078 16829 9138 18667
rect 9259 17372 9325 17373
rect 9259 17308 9260 17372
rect 9324 17308 9325 17372
rect 9259 17307 9325 17308
rect 9075 16828 9141 16829
rect 9075 16764 9076 16828
rect 9140 16764 9141 16828
rect 9075 16763 9141 16764
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7603 14380 7669 14381
rect 7603 14316 7604 14380
rect 7668 14316 7669 14380
rect 7603 14315 7669 14316
rect 7944 14176 8264 15200
rect 8339 15196 8405 15197
rect 8339 15132 8340 15196
rect 8404 15132 8405 15196
rect 8339 15131 8405 15132
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7419 11388 7485 11389
rect 7419 11324 7420 11388
rect 7484 11324 7485 11388
rect 7419 11323 7485 11324
rect 7235 11252 7301 11253
rect 7235 11188 7236 11252
rect 7300 11188 7301 11252
rect 7235 11187 7301 11188
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 8342 9213 8402 15131
rect 9262 15061 9322 17307
rect 9259 15060 9325 15061
rect 9259 14996 9260 15060
rect 9324 14996 9325 15060
rect 9259 14995 9325 14996
rect 8339 9212 8405 9213
rect 8339 9148 8340 9212
rect 8404 9148 8405 9212
rect 8339 9147 8405 9148
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 6499 8668 6565 8669
rect 6499 8604 6500 8668
rect 6564 8604 6565 8668
rect 6499 8603 6565 8604
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 7648 8264 8672
rect 9446 8261 9506 20707
rect 9627 19412 9693 19413
rect 9627 19348 9628 19412
rect 9692 19348 9693 19412
rect 9627 19347 9693 19348
rect 9630 16285 9690 19347
rect 9627 16284 9693 16285
rect 9627 16220 9628 16284
rect 9692 16220 9693 16284
rect 9627 16219 9693 16220
rect 9627 16148 9693 16149
rect 9627 16084 9628 16148
rect 9692 16084 9693 16148
rect 9627 16083 9693 16084
rect 9630 12205 9690 16083
rect 9627 12204 9693 12205
rect 9627 12140 9628 12204
rect 9692 12140 9693 12204
rect 9627 12139 9693 12140
rect 9814 8941 9874 23699
rect 10547 21860 10613 21861
rect 10547 21796 10548 21860
rect 10612 21796 10613 21860
rect 10547 21795 10613 21796
rect 10550 16149 10610 21795
rect 11654 17917 11714 24923
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22139 23492 22205 23493
rect 22139 23428 22140 23492
rect 22204 23428 22205 23492
rect 22139 23427 22205 23428
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17171 22540 17237 22541
rect 17171 22476 17172 22540
rect 17236 22476 17237 22540
rect 17171 22475 17237 22476
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 17174 22269 17234 22475
rect 17171 22268 17237 22269
rect 17171 22204 17172 22268
rect 17236 22204 17237 22268
rect 17171 22203 17237 22204
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 13859 20772 13925 20773
rect 13859 20708 13860 20772
rect 13924 20708 13925 20772
rect 13859 20707 13925 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 11651 17916 11717 17917
rect 11651 17852 11652 17916
rect 11716 17852 11717 17916
rect 11651 17851 11717 17852
rect 11654 16829 11714 17851
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 11651 16828 11717 16829
rect 11651 16764 11652 16828
rect 11716 16764 11717 16828
rect 11651 16763 11717 16764
rect 10547 16148 10613 16149
rect 10547 16084 10548 16148
rect 10612 16084 10613 16148
rect 10547 16083 10613 16084
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 13862 10165 13922 20707
rect 17174 16285 17234 22203
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17171 16284 17237 16285
rect 17171 16220 17172 16284
rect 17236 16220 17237 16284
rect 17171 16219 17237 16220
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 13859 10164 13925 10165
rect 13859 10100 13860 10164
rect 13924 10100 13925 10164
rect 13859 10099 13925 10100
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 9811 8940 9877 8941
rect 9811 8876 9812 8940
rect 9876 8876 9877 8940
rect 9811 8875 9877 8876
rect 9443 8260 9509 8261
rect 9443 8196 9444 8260
rect 9508 8196 9509 8260
rect 9443 8195 9509 8196
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 9824 18264 10848
rect 22142 10709 22202 23427
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22691 21860 22757 21861
rect 22691 21796 22692 21860
rect 22756 21796 22757 21860
rect 22691 21795 22757 21796
rect 22507 16828 22573 16829
rect 22507 16764 22508 16828
rect 22572 16764 22573 16828
rect 22507 16763 22573 16764
rect 22510 13973 22570 16763
rect 22507 13972 22573 13973
rect 22507 13908 22508 13972
rect 22572 13908 22573 13972
rect 22507 13907 22573 13908
rect 22139 10708 22205 10709
rect 22139 10644 22140 10708
rect 22204 10644 22205 10708
rect 22139 10643 22205 10644
rect 22694 10301 22754 21795
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22691 10300 22757 10301
rect 22691 10236 22692 10300
rect 22756 10236 22757 10300
rect 22691 10235 22757 10236
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1676037725
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 10672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 4140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 3404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 6072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 4232 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _132_
timestamp 1676037725
transform 1 0 8372 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1676037725
transform 1 0 2208 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _134_
timestamp 1676037725
transform 1 0 5888 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _135_
timestamp 1676037725
transform 1 0 3404 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 33764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 32292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 31280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 34592 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 33028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _147_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _149_
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1676037725
transform 1 0 18584 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _151_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1676037725
transform 1 0 33580 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1676037725
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 4876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1676037725
transform 1 0 3864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1676037725
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1676037725
transform 1 0 1656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1676037725
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1676037725
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1676037725
transform 1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1676037725
transform 1 0 3128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1676037725
transform 1 0 33672 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 32200 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 35052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1676037725
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform 1 0 22448 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform 1 0 31556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform 1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 11132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 9016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 3036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 5152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 9016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 6440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 13800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
timestamp 1676037725
transform 1 0 22816 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1676037725
transform 1 0 28520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 28336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
timestamp 1676037725
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 14996 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold4_A
timestamp 1676037725
transform 1 0 48484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold6_A
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 4140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 34868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 36984 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 33396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 33580 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 35328 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 36616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 34684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 37904 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 36984 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 31832 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 38548 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 36800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 37260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 38180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 38916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 39836 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 40296 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 41768 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 32752 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 33396 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 25944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 47748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 43516 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 44988 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 48668 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 48024 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1676037725
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1676037725
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1676037725
transform 1 0 7728 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1676037725
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1676037725
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1676037725
transform 1 0 10856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 1676037725
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output142_A
timestamp 1676037725
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 21896 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 27876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 30912 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30820 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 31740 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 30728 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 31556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 32844 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 21620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20056 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 4140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 27600 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14168 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 36800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_19.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 33028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 32016 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_49.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 31464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 30912 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 30544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 26128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l2_in_1__S
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22724 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 27416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 3864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 30176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 32936 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 31096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 19872 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 1472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 32844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 33028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22448 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4140 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5336 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 5428 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 7360 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9568 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4232 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 6808 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 4048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10580 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14260 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9384 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10856 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 6716 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28612 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8740 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 26956 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 25760 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 22908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22172 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 14720 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 8464 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 13616 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 19504 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 19596 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 24932 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1676037725
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1676037725
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1676037725
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1676037725
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1676037725
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1676037725
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_395
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_407
timestamp 1676037725
transform 1 0 38548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_67
timestamp 1676037725
transform 1 0 7268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1676037725
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_142
timestamp 1676037725
transform 1 0 14168 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1676037725
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp 1676037725
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1676037725
transform 1 0 19504 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1676037725
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_31
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_43
timestamp 1676037725
transform 1 0 5060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_67
timestamp 1676037725
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1676037725
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_120
timestamp 1676037725
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1676037725
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_28
timestamp 1676037725
transform 1 0 3680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_40
timestamp 1676037725
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1676037725
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1676037725
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1676037725
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1676037725
transform 1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1676037725
transform 1 0 24840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1676037725
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1676037725
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1676037725
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1676037725
transform 1 0 15548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp 1676037725
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1676037725
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_238
timestamp 1676037725
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1676037725
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1676037725
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1676037725
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1676037725
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1676037725
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1676037725
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_199
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_211
timestamp 1676037725
transform 1 0 20516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_225
timestamp 1676037725
transform 1 0 21804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_237
timestamp 1676037725
transform 1 0 22908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1676037725
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1676037725
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1676037725
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 1676037725
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 1676037725
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1676037725
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp 1676037725
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_238
timestamp 1676037725
transform 1 0 23000 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_250
timestamp 1676037725
transform 1 0 24104 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_262
timestamp 1676037725
transform 1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1676037725
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1676037725
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1676037725
transform 1 0 3128 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_35
timestamp 1676037725
transform 1 0 4324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_59
timestamp 1676037725
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_71
timestamp 1676037725
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_106
timestamp 1676037725
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_243
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1676037725
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1676037725
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1676037725
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1676037725
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1676037725
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_120
timestamp 1676037725
transform 1 0 12144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_127
timestamp 1676037725
transform 1 0 12788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_133
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_144
timestamp 1676037725
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_8
timestamp 1676037725
transform 1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1676037725
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1676037725
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_40
timestamp 1676037725
transform 1 0 4784 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_52
timestamp 1676037725
transform 1 0 5888 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1676037725
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_68
timestamp 1676037725
transform 1 0 7360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1676037725
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1676037725
transform 1 0 9384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_101
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_120
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_128
timestamp 1676037725
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_145
timestamp 1676037725
transform 1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_161
timestamp 1676037725
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_173
timestamp 1676037725
transform 1 0 17020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1676037725
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_22
timestamp 1676037725
transform 1 0 3128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_28
timestamp 1676037725
transform 1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1676037725
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1676037725
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_45
timestamp 1676037725
transform 1 0 5244 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1676037725
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1676037725
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1676037725
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1676037725
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1676037725
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_129
timestamp 1676037725
transform 1 0 12972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1676037725
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1676037725
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_34
timestamp 1676037725
transform 1 0 4232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_42
timestamp 1676037725
transform 1 0 4968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1676037725
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1676037725
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1676037725
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1676037725
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1676037725
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1676037725
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1676037725
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1676037725
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_19
timestamp 1676037725
transform 1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_24
timestamp 1676037725
transform 1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1676037725
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_44
timestamp 1676037725
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_60
timestamp 1676037725
transform 1 0 6624 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1676037725
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1676037725
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1676037725
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_294
timestamp 1676037725
transform 1 0 28152 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_300
timestamp 1676037725
transform 1 0 28704 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_312
timestamp 1676037725
transform 1 0 29808 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_324
timestamp 1676037725
transform 1 0 30912 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1676037725
transform 1 0 4048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1676037725
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_48
timestamp 1676037725
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_54
timestamp 1676037725
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1676037725
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1676037725
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1676037725
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1676037725
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1676037725
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_143
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_219
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_225
timestamp 1676037725
transform 1 0 21804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_237
timestamp 1676037725
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1676037725
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1676037725
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1676037725
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_42
timestamp 1676037725
transform 1 0 4968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1676037725
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1676037725
transform 1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_116
timestamp 1676037725
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1676037725
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_229
timestamp 1676037725
transform 1 0 22172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_241
timestamp 1676037725
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_253
timestamp 1676037725
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_265
timestamp 1676037725
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1676037725
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_8
timestamp 1676037725
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1676037725
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1676037725
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1676037725
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1676037725
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1676037725
transform 1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1676037725
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_143
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_172
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1676037725
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_235
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_239
timestamp 1676037725
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_334
timestamp 1676037725
transform 1 0 31832 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1676037725
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_28
timestamp 1676037725
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1676037725
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1676037725
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1676037725
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1676037725
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1676037725
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_228
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_251
timestamp 1676037725
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_255
timestamp 1676037725
transform 1 0 24564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_267
timestamp 1676037725
transform 1 0 25668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1676037725
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_34
timestamp 1676037725
transform 1 0 4232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_42
timestamp 1676037725
transform 1 0 4968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1676037725
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_143
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1676037725
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_191
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1676037725
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_255
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_267
timestamp 1676037725
transform 1 0 25668 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_279
timestamp 1676037725
transform 1 0 26772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_291
timestamp 1676037725
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1676037725
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1676037725
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1676037725
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1676037725
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1676037725
transform 1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1676037725
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1676037725
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1676037725
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_60
timestamp 1676037725
transform 1 0 6624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1676037725
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1676037725
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_120
timestamp 1676037725
transform 1 0 12144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_133
timestamp 1676037725
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_174
timestamp 1676037725
transform 1 0 17112 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1676037725
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_231
timestamp 1676037725
transform 1 0 22356 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1676037725
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_31
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_201
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_229
timestamp 1676037725
transform 1 0 22172 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_234
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_266
timestamp 1676037725
transform 1 0 25576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_278
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1676037725
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1676037725
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1676037725
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_28
timestamp 1676037725
transform 1 0 3680 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1676037725
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1676037725
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1676037725
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_171
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1676037725
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_227
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1676037725
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1676037725
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1676037725
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1676037725
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1676037725
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1676037725
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1676037725
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_72
timestamp 1676037725
transform 1 0 7728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1676037725
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_191
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1676037725
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_210
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_220
timestamp 1676037725
transform 1 0 21344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1676037725
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1676037725
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_277
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_283
timestamp 1676037725
transform 1 0 27140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_295
timestamp 1676037725
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1676037725
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1676037725
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1676037725
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1676037725
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1676037725
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1676037725
transform 1 0 3404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1676037725
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_63
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1676037725
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1676037725
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1676037725
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_171
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_211
timestamp 1676037725
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1676037725
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_257
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_283
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_295
timestamp 1676037725
transform 1 0 28244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_307
timestamp 1676037725
transform 1 0 29348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_319
timestamp 1676037725
transform 1 0 30452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 1676037725
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1676037725
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1676037725
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1676037725
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1676037725
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1676037725
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1676037725
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1676037725
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1676037725
transform 1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_202
timestamp 1676037725
transform 1 0 19688 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1676037725
transform 1 0 20056 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1676037725
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_234
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_237
timestamp 1676037725
transform 1 0 22908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_255
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1676037725
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1676037725
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_63
timestamp 1676037725
transform 1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1676037725
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1676037725
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1676037725
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_250
timestamp 1676037725
transform 1 0 24104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_256
timestamp 1676037725
transform 1 0 24656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_283
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1676037725
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_290
timestamp 1676037725
transform 1 0 27784 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_302
timestamp 1676037725
transform 1 0 28888 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_314
timestamp 1676037725
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1676037725
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1676037725
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1676037725
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1676037725
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1676037725
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_91
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_95
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1676037725
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1676037725
transform 1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1676037725
transform 1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1676037725
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1676037725
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1676037725
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1676037725
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1676037725
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1676037725
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1676037725
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1676037725
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1676037725
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1676037725
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_133
timestamp 1676037725
transform 1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1676037725
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1676037725
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_240
timestamp 1676037725
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_250
timestamp 1676037725
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_276
timestamp 1676037725
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1676037725
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_310
timestamp 1676037725
transform 1 0 29624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_314
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_326
timestamp 1676037725
transform 1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1676037725
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1676037725
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1676037725
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1676037725
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1676037725
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1676037725
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1676037725
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1676037725
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_158
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_255
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1676037725
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1676037725
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1676037725
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1676037725
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1676037725
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1676037725
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1676037725
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1676037725
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_79
timestamp 1676037725
transform 1 0 8372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1676037725
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1676037725
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_127
timestamp 1676037725
transform 1 0 12788 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1676037725
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1676037725
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_230
timestamp 1676037725
transform 1 0 22264 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_234
timestamp 1676037725
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1676037725
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1676037725
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_286
timestamp 1676037725
transform 1 0 27416 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_326
timestamp 1676037725
transform 1 0 31096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1676037725
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1676037725
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1676037725
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1676037725
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_99
timestamp 1676037725
transform 1 0 10212 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp 1676037725
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1676037725
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1676037725
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_216
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1676037725
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_262
timestamp 1676037725
transform 1 0 25208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1676037725
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_324
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_336
timestamp 1676037725
transform 1 0 32016 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_348
timestamp 1676037725
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1676037725
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1676037725
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1676037725
transform 1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_135
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_142
timestamp 1676037725
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_178
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1676037725
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1676037725
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1676037725
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_274
timestamp 1676037725
transform 1 0 26312 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_283
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_288
timestamp 1676037725
transform 1 0 27600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_315
timestamp 1676037725
transform 1 0 30084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_322
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1676037725
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1676037725
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1676037725
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_35
timestamp 1676037725
transform 1 0 4324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1676037725
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1676037725
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1676037725
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_166
timestamp 1676037725
transform 1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1676037725
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1676037725
transform 1 0 23184 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_293
timestamp 1676037725
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_314
timestamp 1676037725
transform 1 0 29992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_331
timestamp 1676037725
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_343
timestamp 1676037725
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1676037725
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1676037725
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_80
timestamp 1676037725
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_123
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_182
timestamp 1676037725
transform 1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_245
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_250
timestamp 1676037725
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1676037725
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1676037725
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1676037725
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_339
timestamp 1676037725
transform 1 0 32292 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_351
timestamp 1676037725
transform 1 0 33396 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_363
timestamp 1676037725
transform 1 0 34500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_375
timestamp 1676037725
transform 1 0 35604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_387
timestamp 1676037725
transform 1 0 36708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_45
timestamp 1676037725
transform 1 0 5244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_108
timestamp 1676037725
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_114
timestamp 1676037725
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_144
timestamp 1676037725
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1676037725
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1676037725
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1676037725
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_226
timestamp 1676037725
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_269
timestamp 1676037725
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1676037725
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1676037725
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_337
timestamp 1676037725
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_344
timestamp 1676037725
transform 1 0 32752 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_348
timestamp 1676037725
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1676037725
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1676037725
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_61
timestamp 1676037725
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_67
timestamp 1676037725
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_91
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_104
timestamp 1676037725
transform 1 0 10672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_129
timestamp 1676037725
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1676037725
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1676037725
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_211
timestamp 1676037725
transform 1 0 20516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_275
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_330
timestamp 1676037725
transform 1 0 31464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_343
timestamp 1676037725
transform 1 0 32660 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_355
timestamp 1676037725
transform 1 0 33764 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_367
timestamp 1676037725
transform 1 0 34868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_379
timestamp 1676037725
transform 1 0 35972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1676037725
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_507
timestamp 1676037725
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1676037725
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_57
timestamp 1676037725
transform 1 0 6348 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_78
timestamp 1676037725
transform 1 0 8280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1676037725
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_147
timestamp 1676037725
transform 1 0 14628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1676037725
transform 1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1676037725
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1676037725
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_229
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_232
timestamp 1676037725
transform 1 0 22448 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1676037725
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1676037725
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_302
timestamp 1676037725
transform 1 0 28888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_313
timestamp 1676037725
transform 1 0 29900 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_324
timestamp 1676037725
transform 1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_332
timestamp 1676037725
transform 1 0 31648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_340
timestamp 1676037725
transform 1 0 32384 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_352
timestamp 1676037725
transform 1 0 33488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_519
timestamp 1676037725
transform 1 0 48852 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1676037725
transform 1 0 14260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_230
timestamp 1676037725
transform 1 0 22264 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1676037725
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1676037725
transform 1 0 26128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1676037725
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1676037725
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_343
timestamp 1676037725
transform 1 0 32660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_351
timestamp 1676037725
transform 1 0 33396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_363
timestamp 1676037725
transform 1 0 34500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_371
timestamp 1676037725
transform 1 0 35236 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1676037725
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_397
timestamp 1676037725
transform 1 0 37628 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_419
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_423
timestamp 1676037725
transform 1 0 40020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_435
timestamp 1676037725
transform 1 0 41124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_513
timestamp 1676037725
transform 1 0 48300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_519
timestamp 1676037725
transform 1 0 48852 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_87
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_152
timestamp 1676037725
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1676037725
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_281
timestamp 1676037725
transform 1 0 26956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_304
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_331
timestamp 1676037725
transform 1 0 31556 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_337
timestamp 1676037725
transform 1 0 32108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_343
timestamp 1676037725
transform 1 0 32660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_351
timestamp 1676037725
transform 1 0 33396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_359
timestamp 1676037725
transform 1 0 34132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_370
timestamp 1676037725
transform 1 0 35144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_384
timestamp 1676037725
transform 1 0 36432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_392
timestamp 1676037725
transform 1 0 37168 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_395
timestamp 1676037725
transform 1 0 37444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_407
timestamp 1676037725
transform 1 0 38548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_455
timestamp 1676037725
transform 1 0 42964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_463
timestamp 1676037725
transform 1 0 43700 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_473
timestamp 1676037725
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_509
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_512
timestamp 1676037725
transform 1 0 48208 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_517
timestamp 1676037725
transform 1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_8
timestamp 1676037725
transform 1 0 1840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_115
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1676037725
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1676037725
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1676037725
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 1676037725
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_318
timestamp 1676037725
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_326
timestamp 1676037725
transform 1 0 31096 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_331
timestamp 1676037725
transform 1 0 31556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_342
timestamp 1676037725
transform 1 0 32568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_353
timestamp 1676037725
transform 1 0 33580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_360
timestamp 1676037725
transform 1 0 34224 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_368
timestamp 1676037725
transform 1 0 34960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_376
timestamp 1676037725
transform 1 0 35696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_383
timestamp 1676037725
transform 1 0 36340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1676037725
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_395
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_401
timestamp 1676037725
transform 1 0 37996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_409
timestamp 1676037725
transform 1 0 38732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_413
timestamp 1676037725
transform 1 0 39100 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_423
timestamp 1676037725
transform 1 0 40020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_428
timestamp 1676037725
transform 1 0 40480 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_433
timestamp 1676037725
transform 1 0 40940 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_444
timestamp 1676037725
transform 1 0 41952 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_459
timestamp 1676037725
transform 1 0 43332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_467
timestamp 1676037725
transform 1 0 44068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_475
timestamp 1676037725
transform 1 0 44804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_479
timestamp 1676037725
transform 1 0 45172 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_487
timestamp 1676037725
transform 1 0 45908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_495
timestamp 1676037725
transform 1 0 46644 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1676037725
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_511
timestamp 1676037725
transform 1 0 48116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1676037725
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_299
timestamp 1676037725
transform 1 0 28612 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_325
timestamp 1676037725
transform 1 0 31004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_331
timestamp 1676037725
transform 1 0 31556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1676037725
transform 1 0 31924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_346
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1676037725
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_371
timestamp 1676037725
transform 1 0 35236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_379
timestamp 1676037725
transform 1 0 35972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_386
timestamp 1676037725
transform 1 0 36616 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_398
timestamp 1676037725
transform 1 0 37720 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_402
timestamp 1676037725
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_409
timestamp 1676037725
transform 1 0 38732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1676037725
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_437
timestamp 1676037725
transform 1 0 41308 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_446
timestamp 1676037725
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_454
timestamp 1676037725
transform 1 0 42872 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_466
timestamp 1676037725
transform 1 0 43976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1676037725
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1676037725
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_515
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_524
timestamp 1676037725
transform 1 0 49312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold2
timestamp 1676037725
transform 1 0 41124 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform 1 0 41400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1676037725
transform 1 0 48576 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1676037725
transform 1 0 43884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 48392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 35512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 36064 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 36340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 37720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 38364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 40664 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 41308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 28336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 36064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 42596 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1676037725
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 49036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 43700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 44436 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 49036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 48300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 3956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 6532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 3404 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 11960 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 7912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 12144 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21160 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18676 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20056 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25852 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27232 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28244 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37812 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24840 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14628 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4600 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11500 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__194
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11224 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18492 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6808 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__195
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__196
timestamp 1676037725
transform 1 0 36156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__197
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28336 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__198
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27232 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30084 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 26404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__188
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__189
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__169
timestamp 1676037725
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15824 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__175
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11316 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__176
timestamp 1676037725
transform 1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__177
timestamp 1676037725
transform 1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__178
timestamp 1676037725
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 30452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4140 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 6716 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 32936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 4692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32568 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__187
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40866 26200 40922 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 41510 26200 41566 27000 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 test_enable
port 142 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 22856 51000 22976 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 24760 51000 24880 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 17526 6188 17526 6188 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 12466 6188 12466 6188 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 14812 5746 14812 5746 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 14858 7956 14858 7956 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 21298 17680 21298 17680 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 9752 10166 9752 10166 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 21482 16456 21482 16456 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 10304 7922 10304 7922 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 8280 9010 8280 9010 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 5704 12138 5704 12138 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal2 10166 17748 10166 17748 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 6670 12750 6670 12750 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 5842 13804 5842 13804 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 8694 12750 8694 12750 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 6164 16014 6164 16014 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 12650 15861 12650 15861 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 8096 13158 8096 13158 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal2 9982 17408 9982 17408 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel via2 13294 17765 13294 17765 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 8142 20910 8142 20910 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 8050 14314 8050 14314 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8786 9146 8786 9146 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 14306 7412 14306 7412 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 8234 14416 8234 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9338 15096 9338 15096 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10258 14960 10258 14960 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11546 14042 11546 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8142 11186 8142 11186 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8740 11118 8740 11118 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8970 8058 8970 8058 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 8234 9214 8234 9214 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10718 9622 10718 9622 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4416 14042 4416 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4876 11866 4876 11866 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 10810 7344 10810 7344 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 2668 18972 2668 18972 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6762 15470 6762 15470 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7636 15402 7636 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8970 12954 8970 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 5750 14025 5750 14025 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6026 14042 6026 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 6302 11798 6302 11798 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 5474 12614 5474 12614 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 4922 11730 4922 11730 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 5612 15538 5612 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9982 11118 9982 11118 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 10902 7412 10902 7412 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 4784 15402 4784 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6348 13906 6348 13906 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7314 14416 7314 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10074 14790 10074 14790 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 8602 14229 8602 14229 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6946 14008 6946 14008 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9384 12410 9384 12410 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 13386 15912 13386 15912 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8878 14042 8878 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 8786 17578 8786 17578 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10626 18139 10626 18139 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel via3 5267 18020 5267 18020 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 7958 17646 7958 17646 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6302 17306 6302 17306 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7544 15674 7544 15674 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9936 14450 9936 14450 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7544 22610 7544 22610 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6762 17034 6762 17034 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 9430 14807 9430 14807 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11362 17646 11362 17646 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 6256 19482 6256 19482 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 17434 4284 17434 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal2 17710 4114 17710 4114 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 20562 4012 20562 4012 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 26795 4794 26795 4794 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 19964 5882 19964 5882 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 15686 5134 15686 5134 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 18124 3026 18124 3026 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 25047 5338 25047 5338 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25806 7514 25806 7514 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 16468 5678 16468 5678 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 17066 4284 17066 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 25990 4760 25990 4760 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 15456 7854 15456 7854 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 15226 6052 15226 6052 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 23828 5746 23828 5746 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 1426 1894 1426 1894 0 ccff_head
rlabel metal2 48622 25238 48622 25238 0 ccff_head_1
rlabel metal2 49174 21233 49174 21233 0 ccff_tail
rlabel metal2 2254 24252 2254 24252 0 ccff_tail_0
rlabel metal3 1786 1564 1786 1564 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6222 1472 6222 0 chanx_left_in[11]
rlabel metal3 1004 6460 1004 6460 0 chanx_left_in[12]
rlabel metal1 3220 7378 3220 7378 0 chanx_left_in[13]
rlabel metal1 2990 6290 2990 6290 0 chanx_left_in[14]
rlabel metal3 1004 7684 1004 7684 0 chanx_left_in[15]
rlabel via1 2622 6749 2622 6749 0 chanx_left_in[16]
rlabel metal1 2990 7854 2990 7854 0 chanx_left_in[17]
rlabel metal2 1794 7837 1794 7837 0 chanx_left_in[18]
rlabel metal2 2714 7769 2714 7769 0 chanx_left_in[19]
rlabel metal1 3082 2380 3082 2380 0 chanx_left_in[1]
rlabel metal2 1610 9367 1610 9367 0 chanx_left_in[20]
rlabel metal1 2990 8942 2990 8942 0 chanx_left_in[21]
rlabel metal2 2622 8721 2622 8721 0 chanx_left_in[22]
rlabel metal1 1472 8398 1472 8398 0 chanx_left_in[23]
rlabel metal3 1717 11356 1717 11356 0 chanx_left_in[24]
rlabel metal1 1656 10098 1656 10098 0 chanx_left_in[25]
rlabel metal1 1564 12206 1564 12206 0 chanx_left_in[26]
rlabel metal1 1794 7446 1794 7446 0 chanx_left_in[27]
rlabel metal1 1794 7820 1794 7820 0 chanx_left_in[28]
rlabel metal1 1426 12750 1426 12750 0 chanx_left_in[29]
rlabel metal1 2530 2482 2530 2482 0 chanx_left_in[2]
rlabel metal1 1472 2958 1472 2958 0 chanx_left_in[3]
rlabel metal1 1472 3502 1472 3502 0 chanx_left_in[4]
rlabel metal1 2162 4114 2162 4114 0 chanx_left_in[5]
rlabel metal3 1004 4012 1004 4012 0 chanx_left_in[6]
rlabel metal2 1794 4267 1794 4267 0 chanx_left_in[7]
rlabel metal1 1472 4658 1472 4658 0 chanx_left_in[8]
rlabel metal1 1472 5202 1472 5202 0 chanx_left_in[9]
rlabel metal3 1372 13804 1372 13804 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal2 2806 18819 2806 18819 0 chanx_left_out[11]
rlabel metal2 2898 19227 2898 19227 0 chanx_left_out[12]
rlabel metal3 1694 19108 1694 19108 0 chanx_left_out[13]
rlabel metal2 2990 19720 2990 19720 0 chanx_left_out[14]
rlabel metal2 2806 20689 2806 20689 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal3 1717 21148 1717 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal2 4278 22015 4278 22015 0 chanx_left_out[20]
rlabel metal3 1487 22372 1487 22372 0 chanx_left_out[21]
rlabel metal3 2154 22780 2154 22780 0 chanx_left_out[22]
rlabel metal3 1096 23188 1096 23188 0 chanx_left_out[23]
rlabel metal1 9108 20978 9108 20978 0 chanx_left_out[24]
rlabel metal1 4876 17238 4876 17238 0 chanx_left_out[25]
rlabel via2 2806 24395 2806 24395 0 chanx_left_out[26]
rlabel metal2 7222 20135 7222 20135 0 chanx_left_out[27]
rlabel metal1 9246 19414 9246 19414 0 chanx_left_out[28]
rlabel metal1 4140 20502 4140 20502 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 912 15028 912 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 912 15844 912 15844 0 chanx_left_out[5]
rlabel metal3 958 16252 958 16252 0 chanx_left_out[6]
rlabel metal3 912 16660 912 16660 0 chanx_left_out[7]
rlabel metal3 820 17068 820 17068 0 chanx_left_out[8]
rlabel metal3 1372 17476 1372 17476 0 chanx_left_out[9]
rlabel metal1 6118 8398 6118 8398 0 chany_top_in[0]
rlabel metal1 35098 23120 35098 23120 0 chany_top_in[10]
rlabel metal1 29532 24242 29532 24242 0 chany_top_in[11]
rlabel metal2 30268 21828 30268 21828 0 chany_top_in[12]
rlabel metal1 32614 21590 32614 21590 0 chany_top_in[13]
rlabel metal1 34362 22406 34362 22406 0 chany_top_in[14]
rlabel metal1 33488 22066 33488 22066 0 chany_top_in[15]
rlabel metal1 35282 23018 35282 23018 0 chany_top_in[16]
rlabel metal2 33350 24412 33350 24412 0 chany_top_in[17]
rlabel metal2 34086 25245 34086 25245 0 chany_top_in[18]
rlabel metal1 34776 24174 34776 24174 0 chany_top_in[19]
rlabel metal1 28842 21964 28842 21964 0 chany_top_in[1]
rlabel metal1 35466 24106 35466 24106 0 chany_top_in[20]
rlabel metal1 36248 24174 36248 24174 0 chany_top_in[21]
rlabel metal1 36662 23698 36662 23698 0 chany_top_in[22]
rlabel metal1 37490 24174 37490 24174 0 chany_top_in[23]
rlabel metal1 37812 23698 37812 23698 0 chany_top_in[24]
rlabel metal2 38502 25245 38502 25245 0 chany_top_in[25]
rlabel metal2 39238 25245 39238 25245 0 chany_top_in[26]
rlabel metal1 39836 24242 39836 24242 0 chany_top_in[27]
rlabel metal2 40342 25075 40342 25075 0 chany_top_in[28]
rlabel metal1 41676 23698 41676 23698 0 chany_top_in[29]
rlabel metal2 6670 8755 6670 8755 0 chany_top_in[2]
rlabel metal2 17986 23239 17986 23239 0 chany_top_in[3]
rlabel metal2 14490 23749 14490 23749 0 chany_top_in[4]
rlabel metal2 17802 22899 17802 22899 0 chany_top_in[5]
rlabel metal2 29210 24480 29210 24480 0 chany_top_in[6]
rlabel metal1 28428 24174 28428 24174 0 chany_top_in[7]
rlabel metal1 32591 23698 32591 23698 0 chany_top_in[8]
rlabel metal1 32338 21386 32338 21386 0 chany_top_in[9]
rlabel metal1 3634 21454 3634 21454 0 chany_top_out[0]
rlabel metal1 8740 24242 8740 24242 0 chany_top_out[10]
rlabel metal1 9568 23766 9568 23766 0 chany_top_out[11]
rlabel metal2 10718 24497 10718 24497 0 chany_top_out[12]
rlabel metal2 11270 24184 11270 24184 0 chany_top_out[13]
rlabel metal2 12604 21556 12604 21556 0 chany_top_out[14]
rlabel metal2 12558 25034 12558 25034 0 chany_top_out[15]
rlabel metal2 13301 26316 13301 26316 0 chany_top_out[16]
rlabel metal2 13846 25204 13846 25204 0 chany_top_out[17]
rlabel metal1 13570 24276 13570 24276 0 chany_top_out[18]
rlabel metal1 15410 22134 15410 22134 0 chany_top_out[19]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[1]
rlabel metal1 15042 23766 15042 23766 0 chany_top_out[20]
rlabel metal2 16146 24497 16146 24497 0 chany_top_out[21]
rlabel metal2 17211 26316 17211 26316 0 chany_top_out[22]
rlabel metal1 16514 22984 16514 22984 0 chany_top_out[23]
rlabel metal1 17250 23766 17250 23766 0 chany_top_out[24]
rlabel metal1 16468 24242 16468 24242 0 chany_top_out[25]
rlabel metal2 17894 23392 17894 23392 0 chany_top_out[26]
rlabel metal1 20792 22202 20792 22202 0 chany_top_out[27]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[28]
rlabel metal2 22034 25279 22034 25279 0 chany_top_out[29]
rlabel metal1 4048 23766 4048 23766 0 chany_top_out[2]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[3]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[4]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[5]
rlabel metal1 7176 22066 7176 22066 0 chany_top_out[6]
rlabel metal1 6348 24242 6348 24242 0 chany_top_out[7]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[8]
rlabel metal2 8694 24422 8694 24422 0 chany_top_out[9]
rlabel metal1 22448 15538 22448 15538 0 clknet_0_prog_clk
rlabel metal1 8004 9486 8004 9486 0 clknet_4_0_0_prog_clk
rlabel metal1 26174 13226 26174 13226 0 clknet_4_10_0_prog_clk
rlabel metal2 22034 16320 22034 16320 0 clknet_4_11_0_prog_clk
rlabel metal1 19734 19244 19734 19244 0 clknet_4_12_0_prog_clk
rlabel metal1 19734 20502 19734 20502 0 clknet_4_13_0_prog_clk
rlabel metal1 25852 19822 25852 19822 0 clknet_4_14_0_prog_clk
rlabel metal1 21758 22474 21758 22474 0 clknet_4_15_0_prog_clk
rlabel metal1 8372 12614 8372 12614 0 clknet_4_1_0_prog_clk
rlabel metal1 11500 9486 11500 9486 0 clknet_4_2_0_prog_clk
rlabel metal2 14306 13090 14306 13090 0 clknet_4_3_0_prog_clk
rlabel metal1 4554 17646 4554 17646 0 clknet_4_4_0_prog_clk
rlabel metal1 9660 17714 9660 17714 0 clknet_4_5_0_prog_clk
rlabel metal2 14582 19890 14582 19890 0 clknet_4_6_0_prog_clk
rlabel metal2 13754 20196 13754 20196 0 clknet_4_7_0_prog_clk
rlabel metal2 16882 7616 16882 7616 0 clknet_4_8_0_prog_clk
rlabel metal1 19964 12750 19964 12750 0 clknet_4_9_0_prog_clk
rlabel metal2 4094 1622 4094 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 1622 6762 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 9430 1622 9430 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12098 1622 12098 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 25576 2414 25576 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal2 28382 1581 28382 1581 0 gfpga_pad_io_soc_in[1]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[2]
rlabel metal1 33580 2414 33580 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal2 14766 1622 14766 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 17434 1622 17434 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 20102 959 20102 959 0 gfpga_pad_io_soc_out[2]
rlabel metal2 22770 1622 22770 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 36110 1588 36110 1588 0 isol_n
rlabel metal1 6578 2992 6578 2992 0 net1
rlabel metal2 12558 16966 12558 16966 0 net10
rlabel metal1 3726 17170 3726 17170 0 net100
rlabel metal1 4094 16490 4094 16490 0 net101
rlabel metal2 19826 20995 19826 20995 0 net102
rlabel metal1 8648 19346 8648 19346 0 net103
rlabel metal2 3542 15606 3542 15606 0 net104
rlabel metal1 2277 14382 2277 14382 0 net105
rlabel metal1 1794 15028 1794 15028 0 net106
rlabel metal2 3450 14756 3450 14756 0 net107
rlabel metal1 1840 16082 1840 16082 0 net108
rlabel metal1 4002 16592 4002 16592 0 net109
rlabel metal1 11684 16626 11684 16626 0 net11
rlabel metal1 2668 17170 2668 17170 0 net110
rlabel metal1 1794 17680 1794 17680 0 net111
rlabel metal1 1794 18292 1794 18292 0 net112
rlabel metal2 2254 15538 2254 15538 0 net113
rlabel metal2 8372 18428 8372 18428 0 net114
rlabel metal1 4922 11322 4922 11322 0 net115
rlabel metal2 33626 24650 33626 24650 0 net116
rlabel metal2 35006 24616 35006 24616 0 net117
rlabel metal2 33994 24514 33994 24514 0 net118
rlabel via2 17158 16235 17158 16235 0 net119
rlabel metal1 1610 6664 1610 6664 0 net12
rlabel metal2 32522 24276 32522 24276 0 net120
rlabel metal1 27876 22066 27876 22066 0 net121
rlabel metal2 13754 25160 13754 25160 0 net122
rlabel metal2 15226 21420 15226 21420 0 net123
rlabel metal1 2346 24174 2346 24174 0 net124
rlabel metal2 13294 23647 13294 23647 0 net125
rlabel metal1 15962 22610 15962 22610 0 net126
rlabel metal2 14122 21658 14122 21658 0 net127
rlabel metal1 16100 23086 16100 23086 0 net128
rlabel metal1 16698 21590 16698 21590 0 net129
rlabel metal2 2254 7582 2254 7582 0 net13
rlabel metal2 15502 20604 15502 20604 0 net130
rlabel metal3 17388 21828 17388 21828 0 net131
rlabel metal2 20378 22039 20378 22039 0 net132
rlabel metal1 19044 20026 19044 20026 0 net133
rlabel metal1 21896 24174 21896 24174 0 net134
rlabel metal2 3450 17204 3450 17204 0 net135
rlabel metal1 14306 22168 14306 22168 0 net136
rlabel metal2 21206 24293 21206 24293 0 net137
rlabel metal1 1748 10506 1748 10506 0 net138
rlabel metal1 7268 21998 7268 21998 0 net139
rlabel metal1 3910 2550 3910 2550 0 net14
rlabel metal2 1748 23596 1748 23596 0 net140
rlabel metal3 6739 11220 6739 11220 0 net141
rlabel metal2 7038 16252 7038 16252 0 net142
rlabel metal1 4968 2414 4968 2414 0 net143
rlabel metal1 7682 2414 7682 2414 0 net144
rlabel metal1 9706 2414 9706 2414 0 net145
rlabel metal1 12420 2414 12420 2414 0 net146
rlabel metal2 15042 3162 15042 3162 0 net147
rlabel metal1 17204 2822 17204 2822 0 net148
rlabel metal1 19136 2822 19136 2822 0 net149
rlabel metal1 4646 20842 4646 20842 0 net15
rlabel metal1 22356 2414 22356 2414 0 net150
rlabel metal1 21850 21522 21850 21522 0 net151
rlabel metal1 22954 20570 22954 20570 0 net152
rlabel metal1 18469 18258 18469 18258 0 net153
rlabel metal1 23828 21930 23828 21930 0 net154
rlabel metal1 23092 22678 23092 22678 0 net155
rlabel metal1 24610 23834 24610 23834 0 net156
rlabel metal2 25990 21692 25990 21692 0 net157
rlabel metal1 26358 19482 26358 19482 0 net158
rlabel metal1 28658 18394 28658 18394 0 net159
rlabel metal1 5888 16218 5888 16218 0 net16
rlabel metal2 15134 18972 15134 18972 0 net160
rlabel metal1 20010 17578 20010 17578 0 net161
rlabel metal1 24150 18802 24150 18802 0 net162
rlabel metal1 12673 20570 12673 20570 0 net163
rlabel metal1 19596 16218 19596 16218 0 net164
rlabel metal1 14122 8806 14122 8806 0 net165
rlabel metal1 14168 8466 14168 8466 0 net166
rlabel metal1 10580 6834 10580 6834 0 net167
rlabel metal2 11914 8194 11914 8194 0 net168
rlabel metal2 13570 12002 13570 12002 0 net169
rlabel metal2 2254 8160 2254 8160 0 net17
rlabel metal1 13432 7514 13432 7514 0 net170
rlabel metal1 17020 16626 17020 16626 0 net171
rlabel metal2 15410 16677 15410 16677 0 net172
rlabel metal1 15180 15470 15180 15470 0 net173
rlabel metal1 9568 11866 9568 11866 0 net174
rlabel metal2 9430 10030 9430 10030 0 net175
rlabel metal2 8142 15725 8142 15725 0 net176
rlabel metal2 12282 15334 12282 15334 0 net177
rlabel metal3 17802 17544 17802 17544 0 net178
rlabel metal2 19918 15861 19918 15861 0 net179
rlabel metal2 1518 16610 1518 16610 0 net18
rlabel metal1 5290 16966 5290 16966 0 net180
rlabel metal1 12512 8466 12512 8466 0 net181
rlabel metal3 6417 20740 6417 20740 0 net182
rlabel metal3 15870 21692 15870 21692 0 net183
rlabel metal2 9706 19805 9706 19805 0 net184
rlabel metal1 10534 18258 10534 18258 0 net185
rlabel metal1 13110 11798 13110 11798 0 net186
rlabel metal1 10350 15538 10350 15538 0 net187
rlabel metal1 14030 12206 14030 12206 0 net188
rlabel metal1 16284 8602 16284 8602 0 net189
rlabel metal1 13110 16626 13110 16626 0 net19
rlabel metal1 7452 10778 7452 10778 0 net190
rlabel metal1 5750 12886 5750 12886 0 net191
rlabel metal2 16514 14756 16514 14756 0 net192
rlabel metal2 13202 13192 13202 13192 0 net193
rlabel metal1 27922 16558 27922 16558 0 net194
rlabel metal2 32338 24548 32338 24548 0 net195
rlabel via2 15962 21573 15962 21573 0 net196
rlabel metal1 14674 20774 14674 20774 0 net197
rlabel metal1 17158 18802 17158 18802 0 net198
rlabel metal2 43286 24004 43286 24004 0 net199
rlabel metal1 44735 23086 44735 23086 0 net2
rlabel metal1 14812 18598 14812 18598 0 net20
rlabel metal1 1656 24038 1656 24038 0 net200
rlabel metal1 42366 23698 42366 23698 0 net201
rlabel metal1 48668 23086 48668 23086 0 net202
rlabel metal2 44574 22848 44574 22848 0 net203
rlabel metal1 3864 3026 3864 3026 0 net204
rlabel metal1 8142 2958 8142 2958 0 net205
rlabel metal1 6992 16626 6992 16626 0 net21
rlabel metal2 1610 10217 1610 10217 0 net22
rlabel metal1 2162 9486 2162 9486 0 net23
rlabel metal1 20148 16150 20148 16150 0 net24
rlabel metal1 4209 2278 4209 2278 0 net25
rlabel metal2 2438 6426 2438 6426 0 net26
rlabel metal1 1978 3570 1978 3570 0 net27
rlabel metal2 14214 8126 14214 8126 0 net28
rlabel metal1 6762 3910 6762 3910 0 net29
rlabel metal2 13478 5576 13478 5576 0 net3
rlabel metal2 1610 3808 1610 3808 0 net30
rlabel metal1 10626 15402 10626 15402 0 net31
rlabel metal1 9016 14246 9016 14246 0 net32
rlabel via2 13938 20757 13938 20757 0 net33
rlabel via2 14398 23035 14398 23035 0 net34
rlabel metal2 21942 24208 21942 24208 0 net35
rlabel metal2 9890 16524 9890 16524 0 net36
rlabel metal1 28336 20570 28336 20570 0 net37
rlabel metal2 35098 23086 35098 23086 0 net38
rlabel metal1 27462 22542 27462 22542 0 net39
rlabel metal1 6256 13838 6256 13838 0 net4
rlabel metal2 31050 23222 31050 23222 0 net40
rlabel metal2 13616 20774 13616 20774 0 net41
rlabel metal1 15870 18054 15870 18054 0 net42
rlabel metal2 35098 24089 35098 24089 0 net43
rlabel metal1 17480 20978 17480 20978 0 net44
rlabel metal2 35926 24633 35926 24633 0 net45
rlabel metal1 30866 21930 30866 21930 0 net46
rlabel metal2 36754 22576 36754 22576 0 net47
rlabel metal1 37214 24310 37214 24310 0 net48
rlabel metal1 32982 17646 32982 17646 0 net49
rlabel metal1 13800 12818 13800 12818 0 net5
rlabel metal1 18584 15878 18584 15878 0 net50
rlabel metal2 21574 24905 21574 24905 0 net51
rlabel metal1 19780 19754 19780 19754 0 net52
rlabel metal1 40710 23596 40710 23596 0 net53
rlabel metal1 38180 23562 38180 23562 0 net54
rlabel metal2 13570 24123 13570 24123 0 net55
rlabel metal1 13156 20026 13156 20026 0 net56
rlabel metal2 14306 24582 14306 24582 0 net57
rlabel metal1 25760 24106 25760 24106 0 net58
rlabel metal1 26036 23086 26036 23086 0 net59
rlabel metal1 3588 6902 3588 6902 0 net6
rlabel metal1 26772 23018 26772 23018 0 net60
rlabel metal2 25806 23290 25806 23290 0 net61
rlabel metal1 14536 21930 14536 21930 0 net62
rlabel metal1 25116 5610 25116 5610 0 net63
rlabel metal1 28014 2618 28014 2618 0 net64
rlabel metal1 29808 2618 29808 2618 0 net65
rlabel metal2 33534 3842 33534 3842 0 net66
rlabel metal1 33994 2482 33994 2482 0 net67
rlabel metal2 42642 23562 42642 23562 0 net68
rlabel metal2 45402 21369 45402 21369 0 net69
rlabel metal1 5658 7242 5658 7242 0 net7
rlabel metal1 45540 24072 45540 24072 0 net70
rlabel metal1 35880 18734 35880 18734 0 net71
rlabel metal2 31786 19465 31786 19465 0 net72
rlabel metal2 47058 20502 47058 20502 0 net73
rlabel metal2 21482 15555 21482 15555 0 net74
rlabel metal2 41446 20808 41446 20808 0 net75
rlabel metal2 44666 20553 44666 20553 0 net76
rlabel metal2 49266 20944 49266 20944 0 net77
rlabel metal2 47242 19992 47242 19992 0 net78
rlabel metal2 48346 19822 48346 19822 0 net79
rlabel metal1 3634 6426 3634 6426 0 net8
rlabel metal1 35880 18904 35880 18904 0 net80
rlabel metal1 47794 21318 47794 21318 0 net81
rlabel metal1 7130 20774 7130 20774 0 net82
rlabel metal1 1886 13294 1886 13294 0 net83
rlabel metal2 14490 18989 14490 18989 0 net84
rlabel metal1 1978 19346 1978 19346 0 net85
rlabel metal2 4462 19873 4462 19873 0 net86
rlabel metal2 1794 21964 1794 21964 0 net87
rlabel metal1 1840 20910 1840 20910 0 net88
rlabel metal1 1794 21590 1794 21590 0 net89
rlabel metal2 13386 14790 13386 14790 0 net9
rlabel metal1 3818 20434 3818 20434 0 net90
rlabel metal1 2898 21998 2898 21998 0 net91
rlabel metal2 3450 22916 3450 22916 0 net92
rlabel metal1 12696 22066 12696 22066 0 net93
rlabel metal1 1840 13906 1840 13906 0 net94
rlabel metal1 3358 21930 3358 21930 0 net95
rlabel metal2 3634 16150 3634 16150 0 net96
rlabel metal2 6118 21148 6118 21148 0 net97
rlabel viali 6670 19333 6670 19333 0 net98
rlabel metal1 9614 20876 9614 20876 0 net99
rlabel metal2 38778 2098 38778 2098 0 prog_clk
rlabel metal1 41492 24174 41492 24174 0 prog_reset
rlabel metal1 18722 16966 18722 16966 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal1 25760 19890 25760 19890 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal1 28750 16626 28750 16626 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal2 16652 21420 16652 21420 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal2 17434 23324 17434 23324 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal2 17158 23902 17158 23902 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 18492 22542 18492 22542 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel metal1 19044 23766 19044 23766 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 15088 20978 15088 20978 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel metal1 20930 22746 20930 22746 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel metal1 18032 22202 18032 22202 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal2 23782 23358 23782 23358 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 23920 21454 23920 21454 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal1 23828 21590 23828 21590 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal1 26818 18802 26818 18802 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal1 26680 20366 26680 20366 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 18308 19890 18308 19890 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 19918 19278 19918 19278 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 27094 21114 27094 21114 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal1 27738 19958 27738 19958 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel metal2 26634 23392 26634 23392 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal1 27462 22202 27462 22202 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal2 29026 23715 29026 23715 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal1 28842 23494 28842 23494 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal2 30130 21930 30130 21930 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel metal1 31096 22134 31096 22134 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 26956 19414 26956 19414 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal2 30222 20842 30222 20842 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel metal1 28612 18054 28612 18054 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal1 29348 19142 29348 19142 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal1 19688 19890 19688 19890 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel metal2 19734 21148 19734 21148 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 28842 17408 28842 17408 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal2 20654 19822 20654 19822 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal1 21804 19890 21804 19890 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 19090 20332 19090 20332 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal1 25070 15062 25070 15062 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal1 37122 22542 37122 22542 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 20654 16082 20654 16082 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 20654 13804 20654 13804 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal1 17250 9962 17250 9962 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal1 20010 11832 20010 11832 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 21436 12750 21436 12750 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal2 16330 9724 16330 9724 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal1 20470 14450 20470 14450 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 15548 10098 15548 10098 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel metal2 14766 9010 14766 9010 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 16606 12495 16606 12495 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal2 15042 9996 15042 9996 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 17473 13702 17473 13702 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal1 15630 13498 15630 13498 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 21206 9690 21206 9690 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 25162 14416 25162 14416 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 13984 7922 13984 7922 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 18124 15334 18124 15334 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal2 17342 14722 17342 14722 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal2 16330 14620 16330 14620 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal1 14904 14926 14904 14926 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 15042 13158 15042 13158 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal1 15502 13362 15502 13362 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 12558 11628 12558 11628 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal2 12098 11900 12098 11900 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 13432 9418 13432 9418 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal2 12006 9860 12006 9860 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12834 13974 12834 13974 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal1 12328 13226 12328 13226 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 12650 17238 12650 17238 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal1 13662 14586 13662 14586 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 10994 19822 10994 19822 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal2 13754 18564 13754 18564 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal2 10902 20060 10902 20060 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal2 11178 19516 11178 19516 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 4830 18666 4830 18666 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal1 8004 16014 8004 16014 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal1 19688 13226 19688 13226 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal1 23322 13838 23322 13838 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 18538 12750 18538 12750 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 7130 21590 7130 21590 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel metal1 7406 18598 7406 18598 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 10304 22950 10304 22950 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel metal1 9430 21624 9430 21624 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal2 13386 20672 13386 20672 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel metal1 14168 22066 14168 22066 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 15180 19890 15180 19890 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal1 14536 20366 14536 20366 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 16790 17714 16790 17714 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal1 16376 19686 16376 19686 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16376 17238 16376 17238 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 21942 14824 21942 14824 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal1 21390 17068 21390 17068 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 20424 15402 20424 15402 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 23874 14518 23874 14518 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 20378 10268 20378 10268 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel metal2 3726 13158 3726 13158 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 30774 19720 30774 19720 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27278 16422 27278 16422 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18170 18360 18170 18360 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 4324 12886 4324 12886 0 sb_8__0_.mux_left_track_11.out
rlabel metal2 12374 24242 12374 24242 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4186 12257 4186 12257 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 18538 18020 18538 18020 0 sb_8__0_.mux_left_track_13.out
rlabel metal1 16192 21658 16192 21658 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 15594 21403 15594 21403 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6440 21998 6440 21998 0 sb_8__0_.mux_left_track_15.out
rlabel metal1 15180 20774 15180 20774 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17342 20961 17342 20961 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3864 12886 3864 12886 0 sb_8__0_.mux_left_track_17.out
rlabel metal2 19734 20791 19734 20791 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14674 15674 14674 15674 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19412 15334 19412 15334 0 sb_8__0_.mux_left_track_19.out
rlabel metal2 22494 21284 22494 21284 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19642 18564 19642 18564 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9890 14314 9890 14314 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 26404 20298 26404 20298 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22310 14416 22310 14416 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 31970 18105 31970 18105 0 sb_8__0_.mux_left_track_3.out
rlabel metal2 17710 20332 17710 20332 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 31878 20587 31878 20587 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12098 17272 12098 17272 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 27278 21420 27278 21420 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17158 17459 17158 17459 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 2231 23460 2231 23460 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 24242 21998 24242 21998 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13754 9860 13754 9860 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 9775 15164 9775 15164 0 sb_8__0_.mux_left_track_35.out
rlabel metal1 30544 22746 30544 22746 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24104 17204 24104 17204 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 21298 15861 21298 15861 0 sb_8__0_.mux_left_track_45.out
rlabel metal1 29578 21862 29578 21862 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22218 16048 22218 16048 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9246 16048 9246 16048 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 26450 20774 26450 20774 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13754 15589 13754 15589 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6302 14994 6302 14994 0 sb_8__0_.mux_left_track_49.out
rlabel metal2 30222 19516 30222 19516 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21574 15640 21574 15640 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16882 21862 16882 21862 0 sb_8__0_.mux_left_track_5.out
rlabel metal1 17250 20570 17250 20570 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16192 16252 16192 16252 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14030 14926 14030 14926 0 sb_8__0_.mux_left_track_51.out
rlabel metal1 21206 17782 21206 17782 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16376 16082 16376 16082 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6992 16422 6992 16422 0 sb_8__0_.mux_left_track_7.out
rlabel metal1 22586 19414 22586 19414 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 19482 22862 19482 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14858 18666 14858 18666 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11546 17714 11546 17714 0 sb_8__0_.mux_left_track_9.out
rlabel metal2 18538 20383 18538 20383 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13570 12954 13570 12954 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16054 17850 16054 17850 0 sb_8__0_.mux_top_track_0.out
rlabel metal2 27094 17408 27094 17408 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27738 16490 27738 16490 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26634 16456 26634 16456 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22862 17646 22862 17646 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23598 18938 23598 18938 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18906 16082 18906 16082 0 sb_8__0_.mux_top_track_10.out
rlabel metal2 22126 13175 22126 13175 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21114 13498 21114 13498 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20102 12614 20102 12614 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15134 9078 15134 9078 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17388 11526 17388 11526 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel via2 14582 16677 14582 16677 0 sb_8__0_.mux_top_track_12.out
rlabel metal1 16100 10574 16100 10574 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14858 8602 14858 8602 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15318 13838 15318 13838 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12696 13124 12696 13124 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 15088 10778 15088 10778 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14766 10608 14766 10608 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15962 14620 15962 14620 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 10994 15963 10994 15963 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 17710 11594 17710 11594 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12673 12818 12673 12818 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11822 14518 11822 14518 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21850 16014 21850 16014 0 sb_8__0_.mux_top_track_18.out
rlabel metal2 17894 16762 17894 16762 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13202 13804 13202 13804 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17572 19788 17572 19788 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19090 19652 19090 19652 0 sb_8__0_.mux_top_track_2.out
rlabel metal1 24840 13974 24840 13974 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25392 14042 25392 14042 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22080 9622 22080 9622 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15134 8058 15134 8058 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19182 19346 19182 19346 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33718 21998 33718 21998 0 sb_8__0_.mux_top_track_20.out
rlabel metal1 15916 15674 15916 15674 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13110 15062 13110 15062 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34914 22746 34914 22746 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 14398 13804 14398 13804 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19044 14382 19044 14382 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 9430 13277 9430 13277 0 sb_8__0_.mux_top_track_24.out
rlabel metal2 13754 14144 13754 14144 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13662 14382 13662 14382 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32660 23018 32660 23018 0 sb_8__0_.mux_top_track_26.out
rlabel metal2 10626 11934 10626 11934 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 3887 20740 3887 20740 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33074 21862 33074 21862 0 sb_8__0_.mux_top_track_28.out
rlabel metal1 10442 10234 10442 10234 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11362 10098 11362 10098 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32982 23086 32982 23086 0 sb_8__0_.mux_top_track_30.out
rlabel metal2 12558 13872 12558 13872 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 12098 15589 12098 15589 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32568 21114 32568 21114 0 sb_8__0_.mux_top_track_32.out
rlabel metal1 12742 15130 12742 15130 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32706 19533 32706 19533 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33074 23630 33074 23630 0 sb_8__0_.mux_top_track_34.out
rlabel metal2 12558 18343 12558 18343 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 11454 19397 11454 19397 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2185 11254 2185 11254 0 sb_8__0_.mux_top_track_36.out
rlabel metal1 10764 18870 10764 18870 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 1794 10370 1794 10370 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4738 9554 4738 9554 0 sb_8__0_.mux_top_track_38.out
rlabel metal1 7360 16218 7360 16218 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 5405 10948 5405 10948 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19826 24174 19826 24174 0 sb_8__0_.mux_top_track_4.out
rlabel metal1 20194 12750 20194 12750 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19182 12954 19182 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17388 12954 17388 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15870 13906 15870 13906 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16192 14042 16192 14042 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5474 8602 5474 8602 0 sb_8__0_.mux_top_track_40.out
rlabel metal1 7912 17306 7912 17306 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 1288 16660 1288 16660 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9154 8194 9154 8194 0 sb_8__0_.mux_top_track_42.out
rlabel metal1 8326 21012 8326 21012 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 9453 20740 9453 20740 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32522 17340 32522 17340 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 16514 19482 16514 19482 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11730 19686 11730 19686 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32384 21522 32384 21522 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32890 15181 32890 15181 0 sb_8__0_.mux_top_track_46.out
rlabel metal1 18262 18870 18262 18870 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13386 19040 13386 19040 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32936 21318 32936 21318 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 2024 10574 2024 10574 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 18952 18054 18952 18054 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14214 17306 14214 17306 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15042 18343 15042 18343 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20056 14042 20056 14042 0 sb_8__0_.mux_top_track_50.out
rlabel metal1 20746 18088 20746 18088 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13110 16422 13110 16422 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19642 13872 19642 13872 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 19458 23205 19458 23205 0 sb_8__0_.mux_top_track_6.out
rlabel metal2 20746 16796 20746 16796 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 16558 22862 16558 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20884 15062 20884 15062 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19918 14994 19918 14994 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20148 14790 20148 14790 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19458 18564 19458 18564 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 23322 13396 23322 13396 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23276 13226 23276 13226 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21666 13668 21666 13668 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15594 8534 15594 8534 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20102 13804 20102 13804 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 44758 25340 44758 25340 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 45494 25296 45494 25296 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46368 24174 46368 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 46736 23698 46736 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47564 24174 47564 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal2 47886 25075 47886 25075 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal2 43746 25007 43746 25007 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 44344 23698 44344 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel via2 49082 21981 49082 21981 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 49082 23001 49082 23001 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 49174 22610 49174 22610 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 48346 24259 48346 24259 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 41446 2948 41446 2948 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 44114 2200 44114 2200 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 46782 2166 46782 2166 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 49450 2132 49450 2132 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
