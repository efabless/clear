VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bottom_left_tile
  CLASS BLOCK ;
  FOREIGN bottom_left_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 135.000 BY 135.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.720 10.640 41.320 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.720 10.640 91.320 122.640 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.720 10.640 16.320 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 10.640 66.320 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 10.640 116.320 122.640 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 1.400 135.000 2.000 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 64.640 135.000 65.240 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 85.040 135.000 85.640 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 87.080 135.000 87.680 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 89.120 135.000 89.720 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 91.160 135.000 91.760 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 93.200 135.000 93.800 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 95.240 135.000 95.840 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 97.280 135.000 97.880 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 99.320 135.000 99.920 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 101.360 135.000 101.960 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 103.400 135.000 104.000 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 66.680 135.000 67.280 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 105.440 135.000 106.040 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 107.480 135.000 108.080 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 109.520 135.000 110.120 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 111.560 135.000 112.160 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 113.600 135.000 114.200 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 115.640 135.000 116.240 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 117.680 135.000 118.280 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 119.720 135.000 120.320 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 121.760 135.000 122.360 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 123.800 135.000 124.400 ;
    END
  END chanx_right_in[29]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 68.720 135.000 69.320 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 70.760 135.000 71.360 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 72.800 135.000 73.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 74.840 135.000 75.440 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 76.880 135.000 77.480 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 78.920 135.000 79.520 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 80.960 135.000 81.560 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 83.000 135.000 83.600 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 3.440 135.000 4.040 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 23.840 135.000 24.440 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 25.880 135.000 26.480 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 27.920 135.000 28.520 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 29.960 135.000 30.560 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 32.000 135.000 32.600 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 34.040 135.000 34.640 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 36.080 135.000 36.680 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 38.120 135.000 38.720 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 40.160 135.000 40.760 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 42.200 135.000 42.800 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 5.480 135.000 6.080 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 44.240 135.000 44.840 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 46.280 135.000 46.880 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 48.320 135.000 48.920 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 50.360 135.000 50.960 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 52.400 135.000 53.000 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 54.440 135.000 55.040 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 56.480 135.000 57.080 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 58.520 135.000 59.120 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 60.560 135.000 61.160 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 62.600 135.000 63.200 ;
    END
  END chanx_right_out[29]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 7.520 135.000 8.120 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 9.560 135.000 10.160 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 11.600 135.000 12.200 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 13.640 135.000 14.240 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 15.680 135.000 16.280 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 17.720 135.000 18.320 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 19.760 135.000 20.360 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 21.800 135.000 22.400 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 131.000 63.850 135.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 131.000 82.250 135.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 131.000 84.090 135.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 131.000 85.930 135.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 131.000 87.770 135.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 131.000 89.610 135.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 131.000 91.450 135.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 131.000 93.290 135.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 131.000 95.130 135.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 131.000 96.970 135.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 131.000 98.810 135.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 131.000 65.690 135.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 131.000 100.650 135.000 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 131.000 102.490 135.000 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 131.000 104.330 135.000 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 131.000 106.170 135.000 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 131.000 108.010 135.000 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 131.000 109.850 135.000 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 131.000 111.690 135.000 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 131.000 113.530 135.000 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 131.000 115.370 135.000 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 131.000 117.210 135.000 ;
    END
  END chany_top_in[29]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 131.000 67.530 135.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 131.000 69.370 135.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 131.000 71.210 135.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 131.000 73.050 135.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 131.000 74.890 135.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 131.000 76.730 135.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 131.000 78.570 135.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 131.000 80.410 135.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 131.000 8.650 135.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 131.000 27.050 135.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 131.000 28.890 135.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 131.000 30.730 135.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 131.000 32.570 135.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 131.000 34.410 135.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 131.000 36.250 135.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 131.000 38.090 135.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 131.000 39.930 135.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 131.000 41.770 135.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 131.000 43.610 135.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 131.000 10.490 135.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 131.000 45.450 135.000 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 131.000 47.290 135.000 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 131.000 49.130 135.000 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 131.000 50.970 135.000 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 131.000 52.810 135.000 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 131.000 54.650 135.000 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 131.000 56.490 135.000 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 131.000 58.330 135.000 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 131.000 60.170 135.000 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 131.000 62.010 135.000 ;
    END
  END chany_top_out[29]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 131.000 12.330 135.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 131.000 14.170 135.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 131.000 16.010 135.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 131.000 17.850 135.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 131.000 19.690 135.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 131.000 21.530 135.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 131.000 23.370 135.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 131.000 25.210 135.000 ;
    END
  END chany_top_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END prog_clk
  PIN prog_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 131.000 122.730 135.000 ;
    END
  END prog_reset
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 131.000 124.570 135.000 ;
    END
  END reset
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 125.840 135.000 126.440 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 127.880 135.000 128.480 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 129.920 135.000 130.520 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 131.960 135.000 132.560 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
  PIN test_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 131.000 126.410 135.000 ;
    END
  END test_enable
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 129.260 122.485 ;
      LAYER met1 ;
        RECT 5.520 10.640 132.870 132.220 ;
      LAYER met2 ;
        RECT 7.000 130.720 8.090 132.445 ;
        RECT 8.930 130.720 9.930 132.445 ;
        RECT 10.770 130.720 11.770 132.445 ;
        RECT 12.610 130.720 13.610 132.445 ;
        RECT 14.450 130.720 15.450 132.445 ;
        RECT 16.290 130.720 17.290 132.445 ;
        RECT 18.130 130.720 19.130 132.445 ;
        RECT 19.970 130.720 20.970 132.445 ;
        RECT 21.810 130.720 22.810 132.445 ;
        RECT 23.650 130.720 24.650 132.445 ;
        RECT 25.490 130.720 26.490 132.445 ;
        RECT 27.330 130.720 28.330 132.445 ;
        RECT 29.170 130.720 30.170 132.445 ;
        RECT 31.010 130.720 32.010 132.445 ;
        RECT 32.850 130.720 33.850 132.445 ;
        RECT 34.690 130.720 35.690 132.445 ;
        RECT 36.530 130.720 37.530 132.445 ;
        RECT 38.370 130.720 39.370 132.445 ;
        RECT 40.210 130.720 41.210 132.445 ;
        RECT 42.050 130.720 43.050 132.445 ;
        RECT 43.890 130.720 44.890 132.445 ;
        RECT 45.730 130.720 46.730 132.445 ;
        RECT 47.570 130.720 48.570 132.445 ;
        RECT 49.410 130.720 50.410 132.445 ;
        RECT 51.250 130.720 52.250 132.445 ;
        RECT 53.090 130.720 54.090 132.445 ;
        RECT 54.930 130.720 55.930 132.445 ;
        RECT 56.770 130.720 57.770 132.445 ;
        RECT 58.610 130.720 59.610 132.445 ;
        RECT 60.450 130.720 61.450 132.445 ;
        RECT 62.290 130.720 63.290 132.445 ;
        RECT 64.130 130.720 65.130 132.445 ;
        RECT 65.970 130.720 66.970 132.445 ;
        RECT 67.810 130.720 68.810 132.445 ;
        RECT 69.650 130.720 70.650 132.445 ;
        RECT 71.490 130.720 72.490 132.445 ;
        RECT 73.330 130.720 74.330 132.445 ;
        RECT 75.170 130.720 76.170 132.445 ;
        RECT 77.010 130.720 78.010 132.445 ;
        RECT 78.850 130.720 79.850 132.445 ;
        RECT 80.690 130.720 81.690 132.445 ;
        RECT 82.530 130.720 83.530 132.445 ;
        RECT 84.370 130.720 85.370 132.445 ;
        RECT 86.210 130.720 87.210 132.445 ;
        RECT 88.050 130.720 89.050 132.445 ;
        RECT 89.890 130.720 90.890 132.445 ;
        RECT 91.730 130.720 92.730 132.445 ;
        RECT 93.570 130.720 94.570 132.445 ;
        RECT 95.410 130.720 96.410 132.445 ;
        RECT 97.250 130.720 98.250 132.445 ;
        RECT 99.090 130.720 100.090 132.445 ;
        RECT 100.930 130.720 101.930 132.445 ;
        RECT 102.770 130.720 103.770 132.445 ;
        RECT 104.610 130.720 105.610 132.445 ;
        RECT 106.450 130.720 107.450 132.445 ;
        RECT 108.290 130.720 109.290 132.445 ;
        RECT 110.130 130.720 111.130 132.445 ;
        RECT 111.970 130.720 112.970 132.445 ;
        RECT 113.810 130.720 114.810 132.445 ;
        RECT 115.650 130.720 116.650 132.445 ;
        RECT 117.490 130.720 122.170 132.445 ;
        RECT 123.010 130.720 124.010 132.445 ;
        RECT 124.850 130.720 125.850 132.445 ;
        RECT 126.690 130.720 132.840 132.445 ;
        RECT 7.000 4.280 132.840 130.720 ;
        RECT 7.000 1.515 33.390 4.280 ;
        RECT 34.230 1.515 100.550 4.280 ;
        RECT 101.390 1.515 132.840 4.280 ;
      LAYER met3 ;
        RECT 4.000 131.560 130.600 132.425 ;
        RECT 4.000 130.920 131.000 131.560 ;
        RECT 4.000 130.240 130.600 130.920 ;
        RECT 4.400 129.520 130.600 130.240 ;
        RECT 4.400 128.880 131.000 129.520 ;
        RECT 4.400 128.840 130.600 128.880 ;
        RECT 4.000 127.480 130.600 128.840 ;
        RECT 4.000 126.840 131.000 127.480 ;
        RECT 4.000 125.440 130.600 126.840 ;
        RECT 4.000 124.800 131.000 125.440 ;
        RECT 4.400 123.400 130.600 124.800 ;
        RECT 4.000 122.760 131.000 123.400 ;
        RECT 4.000 121.360 130.600 122.760 ;
        RECT 4.000 120.720 131.000 121.360 ;
        RECT 4.000 119.360 130.600 120.720 ;
        RECT 4.400 119.320 130.600 119.360 ;
        RECT 4.400 118.680 131.000 119.320 ;
        RECT 4.400 117.960 130.600 118.680 ;
        RECT 4.000 117.280 130.600 117.960 ;
        RECT 4.000 116.640 131.000 117.280 ;
        RECT 4.000 115.240 130.600 116.640 ;
        RECT 4.000 114.600 131.000 115.240 ;
        RECT 4.000 113.920 130.600 114.600 ;
        RECT 4.400 113.200 130.600 113.920 ;
        RECT 4.400 112.560 131.000 113.200 ;
        RECT 4.400 112.520 130.600 112.560 ;
        RECT 4.000 111.160 130.600 112.520 ;
        RECT 4.000 110.520 131.000 111.160 ;
        RECT 4.000 109.120 130.600 110.520 ;
        RECT 4.000 108.480 131.000 109.120 ;
        RECT 4.000 107.080 130.600 108.480 ;
        RECT 4.000 106.440 131.000 107.080 ;
        RECT 4.000 105.040 130.600 106.440 ;
        RECT 4.000 104.400 131.000 105.040 ;
        RECT 4.000 103.000 130.600 104.400 ;
        RECT 4.000 102.360 131.000 103.000 ;
        RECT 4.000 100.960 130.600 102.360 ;
        RECT 4.000 100.320 131.000 100.960 ;
        RECT 4.000 98.920 130.600 100.320 ;
        RECT 4.000 98.280 131.000 98.920 ;
        RECT 4.000 96.880 130.600 98.280 ;
        RECT 4.000 96.240 131.000 96.880 ;
        RECT 4.000 94.840 130.600 96.240 ;
        RECT 4.000 94.200 131.000 94.840 ;
        RECT 4.000 92.800 130.600 94.200 ;
        RECT 4.000 92.160 131.000 92.800 ;
        RECT 4.000 90.760 130.600 92.160 ;
        RECT 4.000 90.120 131.000 90.760 ;
        RECT 4.000 88.720 130.600 90.120 ;
        RECT 4.000 88.080 131.000 88.720 ;
        RECT 4.000 86.680 130.600 88.080 ;
        RECT 4.000 86.040 131.000 86.680 ;
        RECT 4.000 84.640 130.600 86.040 ;
        RECT 4.000 84.000 131.000 84.640 ;
        RECT 4.000 82.600 130.600 84.000 ;
        RECT 4.000 81.960 131.000 82.600 ;
        RECT 4.000 80.560 130.600 81.960 ;
        RECT 4.000 79.920 131.000 80.560 ;
        RECT 4.000 78.520 130.600 79.920 ;
        RECT 4.000 77.880 131.000 78.520 ;
        RECT 4.000 76.480 130.600 77.880 ;
        RECT 4.000 75.840 131.000 76.480 ;
        RECT 4.000 74.440 130.600 75.840 ;
        RECT 4.000 73.800 131.000 74.440 ;
        RECT 4.000 72.400 130.600 73.800 ;
        RECT 4.000 71.760 131.000 72.400 ;
        RECT 4.000 70.360 130.600 71.760 ;
        RECT 4.000 69.720 131.000 70.360 ;
        RECT 4.000 68.320 130.600 69.720 ;
        RECT 4.000 67.680 131.000 68.320 ;
        RECT 4.000 66.280 130.600 67.680 ;
        RECT 4.000 65.640 131.000 66.280 ;
        RECT 4.000 64.240 130.600 65.640 ;
        RECT 4.000 63.600 131.000 64.240 ;
        RECT 4.000 62.200 130.600 63.600 ;
        RECT 4.000 61.560 131.000 62.200 ;
        RECT 4.000 60.160 130.600 61.560 ;
        RECT 4.000 59.520 131.000 60.160 ;
        RECT 4.000 58.120 130.600 59.520 ;
        RECT 4.000 57.480 131.000 58.120 ;
        RECT 4.000 56.080 130.600 57.480 ;
        RECT 4.000 55.440 131.000 56.080 ;
        RECT 4.000 54.040 130.600 55.440 ;
        RECT 4.000 53.400 131.000 54.040 ;
        RECT 4.000 52.000 130.600 53.400 ;
        RECT 4.000 51.360 131.000 52.000 ;
        RECT 4.000 49.960 130.600 51.360 ;
        RECT 4.000 49.320 131.000 49.960 ;
        RECT 4.000 47.920 130.600 49.320 ;
        RECT 4.000 47.280 131.000 47.920 ;
        RECT 4.000 45.880 130.600 47.280 ;
        RECT 4.000 45.240 131.000 45.880 ;
        RECT 4.000 43.840 130.600 45.240 ;
        RECT 4.000 43.200 131.000 43.840 ;
        RECT 4.000 41.800 130.600 43.200 ;
        RECT 4.000 41.160 131.000 41.800 ;
        RECT 4.000 39.760 130.600 41.160 ;
        RECT 4.000 39.120 131.000 39.760 ;
        RECT 4.000 37.720 130.600 39.120 ;
        RECT 4.000 37.080 131.000 37.720 ;
        RECT 4.000 35.680 130.600 37.080 ;
        RECT 4.000 35.040 131.000 35.680 ;
        RECT 4.000 33.640 130.600 35.040 ;
        RECT 4.000 33.000 131.000 33.640 ;
        RECT 4.000 31.600 130.600 33.000 ;
        RECT 4.000 30.960 131.000 31.600 ;
        RECT 4.000 29.560 130.600 30.960 ;
        RECT 4.000 28.920 131.000 29.560 ;
        RECT 4.000 27.520 130.600 28.920 ;
        RECT 4.000 26.880 131.000 27.520 ;
        RECT 4.000 25.480 130.600 26.880 ;
        RECT 4.000 24.840 131.000 25.480 ;
        RECT 4.000 23.440 130.600 24.840 ;
        RECT 4.000 22.800 131.000 23.440 ;
        RECT 4.000 21.400 130.600 22.800 ;
        RECT 4.000 20.760 131.000 21.400 ;
        RECT 4.000 19.360 130.600 20.760 ;
        RECT 4.000 18.720 131.000 19.360 ;
        RECT 4.000 17.320 130.600 18.720 ;
        RECT 4.000 16.680 131.000 17.320 ;
        RECT 4.000 15.280 130.600 16.680 ;
        RECT 4.000 14.640 131.000 15.280 ;
        RECT 4.000 13.240 130.600 14.640 ;
        RECT 4.000 12.600 131.000 13.240 ;
        RECT 4.000 11.200 130.600 12.600 ;
        RECT 4.000 10.560 131.000 11.200 ;
        RECT 4.000 9.160 130.600 10.560 ;
        RECT 4.000 8.520 131.000 9.160 ;
        RECT 4.000 7.120 130.600 8.520 ;
        RECT 4.000 6.480 131.000 7.120 ;
        RECT 4.000 5.080 130.600 6.480 ;
        RECT 4.000 4.440 131.000 5.080 ;
        RECT 4.000 3.040 130.600 4.440 ;
        RECT 4.000 2.400 131.000 3.040 ;
        RECT 4.000 1.535 130.600 2.400 ;
      LAYER met4 ;
        RECT 11.335 123.040 123.905 131.745 ;
        RECT 11.335 41.655 14.320 123.040 ;
        RECT 16.720 41.655 39.320 123.040 ;
        RECT 41.720 41.655 64.320 123.040 ;
        RECT 66.720 41.655 89.320 123.040 ;
        RECT 91.720 41.655 114.320 123.040 ;
        RECT 116.720 41.655 123.905 123.040 ;
  END
END bottom_left_tile
END LIBRARY

