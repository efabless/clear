magic
tech sky130A
magscale 1 2
timestamp 1682557371
<< obsli1 >>
rect 1104 2159 25852 54417
<< obsm1 >>
rect 934 1844 26114 54448
<< metal2 >>
rect 1490 56200 1546 57000
rect 1858 56200 1914 57000
rect 2226 56200 2282 57000
rect 2594 56200 2650 57000
rect 2962 56200 3018 57000
rect 3330 56200 3386 57000
rect 3698 56200 3754 57000
rect 4066 56200 4122 57000
rect 4434 56200 4490 57000
rect 4802 56200 4858 57000
rect 5170 56200 5226 57000
rect 5538 56200 5594 57000
rect 5906 56200 5962 57000
rect 6274 56200 6330 57000
rect 6642 56200 6698 57000
rect 7010 56200 7066 57000
rect 7378 56200 7434 57000
rect 7746 56200 7802 57000
rect 8114 56200 8170 57000
rect 8482 56200 8538 57000
rect 8850 56200 8906 57000
rect 9218 56200 9274 57000
rect 9586 56200 9642 57000
rect 9954 56200 10010 57000
rect 10322 56200 10378 57000
rect 10690 56200 10746 57000
rect 11058 56200 11114 57000
rect 11426 56200 11482 57000
rect 11794 56200 11850 57000
rect 12162 56200 12218 57000
rect 12530 56200 12586 57000
rect 12898 56200 12954 57000
rect 13266 56200 13322 57000
rect 13634 56200 13690 57000
rect 14002 56200 14058 57000
rect 14370 56200 14426 57000
rect 14738 56200 14794 57000
rect 15106 56200 15162 57000
rect 15474 56200 15530 57000
rect 15842 56200 15898 57000
rect 16210 56200 16266 57000
rect 16578 56200 16634 57000
rect 16946 56200 17002 57000
rect 17314 56200 17370 57000
rect 17682 56200 17738 57000
rect 18050 56200 18106 57000
rect 18418 56200 18474 57000
rect 18786 56200 18842 57000
rect 19154 56200 19210 57000
rect 19522 56200 19578 57000
rect 19890 56200 19946 57000
rect 20258 56200 20314 57000
rect 20626 56200 20682 57000
rect 20994 56200 21050 57000
rect 21362 56200 21418 57000
rect 21730 56200 21786 57000
rect 22098 56200 22154 57000
rect 22466 56200 22522 57000
rect 22834 56200 22890 57000
rect 23202 56200 23258 57000
rect 23570 56200 23626 57000
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
<< obsm2 >>
rect 938 56144 1434 56273
rect 1602 56144 1802 56273
rect 1970 56144 2170 56273
rect 2338 56144 2538 56273
rect 2706 56144 2906 56273
rect 3074 56144 3274 56273
rect 3442 56144 3642 56273
rect 3810 56144 4010 56273
rect 4178 56144 4378 56273
rect 4546 56144 4746 56273
rect 4914 56144 5114 56273
rect 5282 56144 5482 56273
rect 5650 56144 5850 56273
rect 6018 56144 6218 56273
rect 6386 56144 6586 56273
rect 6754 56144 6954 56273
rect 7122 56144 7322 56273
rect 7490 56144 7690 56273
rect 7858 56144 8058 56273
rect 8226 56144 8426 56273
rect 8594 56144 8794 56273
rect 8962 56144 9162 56273
rect 9330 56144 9530 56273
rect 9698 56144 9898 56273
rect 10066 56144 10266 56273
rect 10434 56144 10634 56273
rect 10802 56144 11002 56273
rect 11170 56144 11370 56273
rect 11538 56144 11738 56273
rect 11906 56144 12106 56273
rect 12274 56144 12474 56273
rect 12642 56144 12842 56273
rect 13010 56144 13210 56273
rect 13378 56144 13578 56273
rect 13746 56144 13946 56273
rect 14114 56144 14314 56273
rect 14482 56144 14682 56273
rect 14850 56144 15050 56273
rect 15218 56144 15418 56273
rect 15586 56144 15786 56273
rect 15954 56144 16154 56273
rect 16322 56144 16522 56273
rect 16690 56144 16890 56273
rect 17058 56144 17258 56273
rect 17426 56144 17626 56273
rect 17794 56144 17994 56273
rect 18162 56144 18362 56273
rect 18530 56144 18730 56273
rect 18898 56144 19098 56273
rect 19266 56144 19466 56273
rect 19634 56144 19834 56273
rect 20002 56144 20202 56273
rect 20370 56144 20570 56273
rect 20738 56144 20938 56273
rect 21106 56144 21306 56273
rect 21474 56144 21674 56273
rect 21842 56144 22042 56273
rect 22210 56144 22410 56273
rect 22578 56144 22778 56273
rect 22946 56144 23146 56273
rect 23314 56144 23514 56273
rect 23682 56144 26108 56273
rect 938 856 26108 56144
rect 938 711 1618 856
rect 1786 711 1986 856
rect 2154 711 2354 856
rect 2522 711 2722 856
rect 2890 711 3090 856
rect 3258 711 3458 856
rect 3626 711 3826 856
rect 3994 711 4194 856
rect 4362 711 4562 856
rect 4730 711 4930 856
rect 5098 711 5298 856
rect 5466 711 5666 856
rect 5834 711 6034 856
rect 6202 711 6402 856
rect 6570 711 6770 856
rect 6938 711 7138 856
rect 7306 711 7506 856
rect 7674 711 7874 856
rect 8042 711 8242 856
rect 8410 711 8610 856
rect 8778 711 8978 856
rect 9146 711 9346 856
rect 9514 711 9714 856
rect 9882 711 10082 856
rect 10250 711 10450 856
rect 10618 711 10818 856
rect 10986 711 11186 856
rect 11354 711 11554 856
rect 11722 711 11922 856
rect 12090 711 12290 856
rect 12458 711 12658 856
rect 12826 711 13026 856
rect 13194 711 13394 856
rect 13562 711 13762 856
rect 13930 711 14130 856
rect 14298 711 14498 856
rect 14666 711 14866 856
rect 15034 711 15234 856
rect 15402 711 15602 856
rect 15770 711 15970 856
rect 16138 711 16338 856
rect 16506 711 16706 856
rect 16874 711 17074 856
rect 17242 711 17442 856
rect 17610 711 17810 856
rect 17978 711 18178 856
rect 18346 711 18546 856
rect 18714 711 18914 856
rect 19082 711 19282 856
rect 19450 711 19650 856
rect 19818 711 20018 856
rect 20186 711 20386 856
rect 20554 711 20754 856
rect 20922 711 21122 856
rect 21290 711 21490 856
rect 21658 711 21858 856
rect 22026 711 22226 856
rect 22394 711 22594 856
rect 22762 711 22962 856
rect 23130 711 23330 856
rect 23498 711 23698 856
rect 23866 711 24066 856
rect 24234 711 24434 856
rect 24602 711 24802 856
rect 24970 711 26108 856
<< metal3 >>
rect 26200 56176 27000 56296
rect 0 55360 800 55480
rect 26200 55360 27000 55480
rect 26200 54544 27000 54664
rect 26200 53728 27000 53848
rect 0 52912 800 53032
rect 26200 52912 27000 53032
rect 26200 52096 27000 52216
rect 26200 51280 27000 51400
rect 0 50464 800 50584
rect 26200 50464 27000 50584
rect 26200 49648 27000 49768
rect 26200 48832 27000 48952
rect 0 48016 800 48136
rect 26200 48016 27000 48136
rect 26200 47200 27000 47320
rect 26200 46384 27000 46504
rect 0 45568 800 45688
rect 26200 45568 27000 45688
rect 26200 44752 27000 44872
rect 26200 43936 27000 44056
rect 0 43120 800 43240
rect 26200 43120 27000 43240
rect 26200 42304 27000 42424
rect 26200 41488 27000 41608
rect 0 40672 800 40792
rect 26200 40672 27000 40792
rect 26200 39856 27000 39976
rect 26200 39040 27000 39160
rect 0 38224 800 38344
rect 26200 38224 27000 38344
rect 26200 37408 27000 37528
rect 26200 36592 27000 36712
rect 0 35776 800 35896
rect 26200 35776 27000 35896
rect 26200 34960 27000 35080
rect 26200 34144 27000 34264
rect 0 33328 800 33448
rect 26200 33328 27000 33448
rect 26200 32512 27000 32632
rect 26200 31696 27000 31816
rect 0 30880 800 31000
rect 26200 30880 27000 31000
rect 26200 30064 27000 30184
rect 26200 29248 27000 29368
rect 0 28432 800 28552
rect 26200 28432 27000 28552
rect 26200 27616 27000 27736
rect 26200 26800 27000 26920
rect 0 25984 800 26104
rect 26200 25984 27000 26104
rect 26200 25168 27000 25288
rect 26200 24352 27000 24472
rect 0 23536 800 23656
rect 26200 23536 27000 23656
rect 26200 22720 27000 22840
rect 26200 21904 27000 22024
rect 0 21088 800 21208
rect 26200 21088 27000 21208
rect 26200 20272 27000 20392
rect 26200 19456 27000 19576
rect 0 18640 800 18760
rect 26200 18640 27000 18760
rect 26200 17824 27000 17944
rect 26200 17008 27000 17128
rect 0 16192 800 16312
rect 26200 16192 27000 16312
rect 26200 15376 27000 15496
rect 26200 14560 27000 14680
rect 0 13744 800 13864
rect 26200 13744 27000 13864
rect 26200 12928 27000 13048
rect 26200 12112 27000 12232
rect 0 11296 800 11416
rect 26200 11296 27000 11416
rect 26200 10480 27000 10600
rect 26200 9664 27000 9784
rect 0 8848 800 8968
rect 26200 8848 27000 8968
rect 26200 8032 27000 8152
rect 26200 7216 27000 7336
rect 0 6400 800 6520
rect 26200 6400 27000 6520
rect 26200 5584 27000 5704
rect 26200 4768 27000 4888
rect 0 3952 800 4072
rect 26200 3952 27000 4072
rect 26200 3136 27000 3256
rect 26200 2320 27000 2440
rect 0 1504 800 1624
rect 26200 1504 27000 1624
rect 26200 688 27000 808
<< obsm3 >>
rect 800 56096 26120 56269
rect 800 55560 26200 56096
rect 880 55280 26120 55560
rect 800 54744 26200 55280
rect 800 54464 26120 54744
rect 800 53928 26200 54464
rect 800 53648 26120 53928
rect 800 53112 26200 53648
rect 880 52832 26120 53112
rect 800 52296 26200 52832
rect 800 52016 26120 52296
rect 800 51480 26200 52016
rect 800 51200 26120 51480
rect 800 50664 26200 51200
rect 880 50384 26120 50664
rect 800 49848 26200 50384
rect 800 49568 26120 49848
rect 800 49032 26200 49568
rect 800 48752 26120 49032
rect 800 48216 26200 48752
rect 880 47936 26120 48216
rect 800 47400 26200 47936
rect 800 47120 26120 47400
rect 800 46584 26200 47120
rect 800 46304 26120 46584
rect 800 45768 26200 46304
rect 880 45488 26120 45768
rect 800 44952 26200 45488
rect 800 44672 26120 44952
rect 800 44136 26200 44672
rect 800 43856 26120 44136
rect 800 43320 26200 43856
rect 880 43040 26120 43320
rect 800 42504 26200 43040
rect 800 42224 26120 42504
rect 800 41688 26200 42224
rect 800 41408 26120 41688
rect 800 40872 26200 41408
rect 880 40592 26120 40872
rect 800 40056 26200 40592
rect 800 39776 26120 40056
rect 800 39240 26200 39776
rect 800 38960 26120 39240
rect 800 38424 26200 38960
rect 880 38144 26120 38424
rect 800 37608 26200 38144
rect 800 37328 26120 37608
rect 800 36792 26200 37328
rect 800 36512 26120 36792
rect 800 35976 26200 36512
rect 880 35696 26120 35976
rect 800 35160 26200 35696
rect 800 34880 26120 35160
rect 800 34344 26200 34880
rect 800 34064 26120 34344
rect 800 33528 26200 34064
rect 880 33248 26120 33528
rect 800 32712 26200 33248
rect 800 32432 26120 32712
rect 800 31896 26200 32432
rect 800 31616 26120 31896
rect 800 31080 26200 31616
rect 880 30800 26120 31080
rect 800 30264 26200 30800
rect 800 29984 26120 30264
rect 800 29448 26200 29984
rect 800 29168 26120 29448
rect 800 28632 26200 29168
rect 880 28352 26120 28632
rect 800 27816 26200 28352
rect 800 27536 26120 27816
rect 800 27000 26200 27536
rect 800 26720 26120 27000
rect 800 26184 26200 26720
rect 880 25904 26120 26184
rect 800 25368 26200 25904
rect 800 25088 26120 25368
rect 800 24552 26200 25088
rect 800 24272 26120 24552
rect 800 23736 26200 24272
rect 880 23456 26120 23736
rect 800 22920 26200 23456
rect 800 22640 26120 22920
rect 800 22104 26200 22640
rect 800 21824 26120 22104
rect 800 21288 26200 21824
rect 880 21008 26120 21288
rect 800 20472 26200 21008
rect 800 20192 26120 20472
rect 800 19656 26200 20192
rect 800 19376 26120 19656
rect 800 18840 26200 19376
rect 880 18560 26120 18840
rect 800 18024 26200 18560
rect 800 17744 26120 18024
rect 800 17208 26200 17744
rect 800 16928 26120 17208
rect 800 16392 26200 16928
rect 880 16112 26120 16392
rect 800 15576 26200 16112
rect 800 15296 26120 15576
rect 800 14760 26200 15296
rect 800 14480 26120 14760
rect 800 13944 26200 14480
rect 880 13664 26120 13944
rect 800 13128 26200 13664
rect 800 12848 26120 13128
rect 800 12312 26200 12848
rect 800 12032 26120 12312
rect 800 11496 26200 12032
rect 880 11216 26120 11496
rect 800 10680 26200 11216
rect 800 10400 26120 10680
rect 800 9864 26200 10400
rect 800 9584 26120 9864
rect 800 9048 26200 9584
rect 880 8768 26120 9048
rect 800 8232 26200 8768
rect 800 7952 26120 8232
rect 800 7416 26200 7952
rect 800 7136 26120 7416
rect 800 6600 26200 7136
rect 880 6320 26120 6600
rect 800 5784 26200 6320
rect 800 5504 26120 5784
rect 800 4968 26200 5504
rect 800 4688 26120 4968
rect 800 4152 26200 4688
rect 880 3872 26120 4152
rect 800 3336 26200 3872
rect 800 3056 26120 3336
rect 800 2520 26200 3056
rect 800 2240 26120 2520
rect 800 1704 26200 2240
rect 880 1424 26120 1704
rect 800 888 26200 1424
rect 800 715 26120 888
<< metal4 >>
rect 2944 2128 3264 54448
rect 7944 2128 8264 54448
rect 12944 2128 13264 54448
rect 17944 2128 18264 54448
rect 22944 2128 23264 54448
<< obsm4 >>
rect 9075 2619 12864 53957
rect 13344 2619 17864 53957
rect 18344 2619 22864 53957
rect 23344 2619 24045 53957
<< labels >>
rlabel metal4 s 7944 2128 8264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 55360 800 55480 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 ccff_head_0
port 4 nsew signal input
rlabel metal3 s 26200 688 27000 808 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 1490 56200 1546 57000 6 ccff_tail_0
port 6 nsew signal output
rlabel metal3 s 26200 25984 27000 26104 6 chanx_right_in[0]
port 7 nsew signal input
rlabel metal3 s 26200 34144 27000 34264 6 chanx_right_in[10]
port 8 nsew signal input
rlabel metal3 s 26200 34960 27000 35080 6 chanx_right_in[11]
port 9 nsew signal input
rlabel metal3 s 26200 35776 27000 35896 6 chanx_right_in[12]
port 10 nsew signal input
rlabel metal3 s 26200 36592 27000 36712 6 chanx_right_in[13]
port 11 nsew signal input
rlabel metal3 s 26200 37408 27000 37528 6 chanx_right_in[14]
port 12 nsew signal input
rlabel metal3 s 26200 38224 27000 38344 6 chanx_right_in[15]
port 13 nsew signal input
rlabel metal3 s 26200 39040 27000 39160 6 chanx_right_in[16]
port 14 nsew signal input
rlabel metal3 s 26200 39856 27000 39976 6 chanx_right_in[17]
port 15 nsew signal input
rlabel metal3 s 26200 40672 27000 40792 6 chanx_right_in[18]
port 16 nsew signal input
rlabel metal3 s 26200 41488 27000 41608 6 chanx_right_in[19]
port 17 nsew signal input
rlabel metal3 s 26200 26800 27000 26920 6 chanx_right_in[1]
port 18 nsew signal input
rlabel metal3 s 26200 42304 27000 42424 6 chanx_right_in[20]
port 19 nsew signal input
rlabel metal3 s 26200 43120 27000 43240 6 chanx_right_in[21]
port 20 nsew signal input
rlabel metal3 s 26200 43936 27000 44056 6 chanx_right_in[22]
port 21 nsew signal input
rlabel metal3 s 26200 44752 27000 44872 6 chanx_right_in[23]
port 22 nsew signal input
rlabel metal3 s 26200 45568 27000 45688 6 chanx_right_in[24]
port 23 nsew signal input
rlabel metal3 s 26200 46384 27000 46504 6 chanx_right_in[25]
port 24 nsew signal input
rlabel metal3 s 26200 47200 27000 47320 6 chanx_right_in[26]
port 25 nsew signal input
rlabel metal3 s 26200 48016 27000 48136 6 chanx_right_in[27]
port 26 nsew signal input
rlabel metal3 s 26200 48832 27000 48952 6 chanx_right_in[28]
port 27 nsew signal input
rlabel metal3 s 26200 49648 27000 49768 6 chanx_right_in[29]
port 28 nsew signal input
rlabel metal3 s 26200 27616 27000 27736 6 chanx_right_in[2]
port 29 nsew signal input
rlabel metal3 s 26200 28432 27000 28552 6 chanx_right_in[3]
port 30 nsew signal input
rlabel metal3 s 26200 29248 27000 29368 6 chanx_right_in[4]
port 31 nsew signal input
rlabel metal3 s 26200 30064 27000 30184 6 chanx_right_in[5]
port 32 nsew signal input
rlabel metal3 s 26200 30880 27000 31000 6 chanx_right_in[6]
port 33 nsew signal input
rlabel metal3 s 26200 31696 27000 31816 6 chanx_right_in[7]
port 34 nsew signal input
rlabel metal3 s 26200 32512 27000 32632 6 chanx_right_in[8]
port 35 nsew signal input
rlabel metal3 s 26200 33328 27000 33448 6 chanx_right_in[9]
port 36 nsew signal input
rlabel metal3 s 26200 1504 27000 1624 6 chanx_right_out[0]
port 37 nsew signal output
rlabel metal3 s 26200 9664 27000 9784 6 chanx_right_out[10]
port 38 nsew signal output
rlabel metal3 s 26200 10480 27000 10600 6 chanx_right_out[11]
port 39 nsew signal output
rlabel metal3 s 26200 11296 27000 11416 6 chanx_right_out[12]
port 40 nsew signal output
rlabel metal3 s 26200 12112 27000 12232 6 chanx_right_out[13]
port 41 nsew signal output
rlabel metal3 s 26200 12928 27000 13048 6 chanx_right_out[14]
port 42 nsew signal output
rlabel metal3 s 26200 13744 27000 13864 6 chanx_right_out[15]
port 43 nsew signal output
rlabel metal3 s 26200 14560 27000 14680 6 chanx_right_out[16]
port 44 nsew signal output
rlabel metal3 s 26200 15376 27000 15496 6 chanx_right_out[17]
port 45 nsew signal output
rlabel metal3 s 26200 16192 27000 16312 6 chanx_right_out[18]
port 46 nsew signal output
rlabel metal3 s 26200 17008 27000 17128 6 chanx_right_out[19]
port 47 nsew signal output
rlabel metal3 s 26200 2320 27000 2440 6 chanx_right_out[1]
port 48 nsew signal output
rlabel metal3 s 26200 17824 27000 17944 6 chanx_right_out[20]
port 49 nsew signal output
rlabel metal3 s 26200 18640 27000 18760 6 chanx_right_out[21]
port 50 nsew signal output
rlabel metal3 s 26200 19456 27000 19576 6 chanx_right_out[22]
port 51 nsew signal output
rlabel metal3 s 26200 20272 27000 20392 6 chanx_right_out[23]
port 52 nsew signal output
rlabel metal3 s 26200 21088 27000 21208 6 chanx_right_out[24]
port 53 nsew signal output
rlabel metal3 s 26200 21904 27000 22024 6 chanx_right_out[25]
port 54 nsew signal output
rlabel metal3 s 26200 22720 27000 22840 6 chanx_right_out[26]
port 55 nsew signal output
rlabel metal3 s 26200 23536 27000 23656 6 chanx_right_out[27]
port 56 nsew signal output
rlabel metal3 s 26200 24352 27000 24472 6 chanx_right_out[28]
port 57 nsew signal output
rlabel metal3 s 26200 25168 27000 25288 6 chanx_right_out[29]
port 58 nsew signal output
rlabel metal3 s 26200 3136 27000 3256 6 chanx_right_out[2]
port 59 nsew signal output
rlabel metal3 s 26200 3952 27000 4072 6 chanx_right_out[3]
port 60 nsew signal output
rlabel metal3 s 26200 4768 27000 4888 6 chanx_right_out[4]
port 61 nsew signal output
rlabel metal3 s 26200 5584 27000 5704 6 chanx_right_out[5]
port 62 nsew signal output
rlabel metal3 s 26200 6400 27000 6520 6 chanx_right_out[6]
port 63 nsew signal output
rlabel metal3 s 26200 7216 27000 7336 6 chanx_right_out[7]
port 64 nsew signal output
rlabel metal3 s 26200 8032 27000 8152 6 chanx_right_out[8]
port 65 nsew signal output
rlabel metal3 s 26200 8848 27000 8968 6 chanx_right_out[9]
port 66 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 chany_bottom_in[0]
port 67 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[10]
port 68 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_in[11]
port 69 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 chany_bottom_in[12]
port 70 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[13]
port 71 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[14]
port 72 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[15]
port 73 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[16]
port 74 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 chany_bottom_in[17]
port 75 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[18]
port 76 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[19]
port 77 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 chany_bottom_in[1]
port 78 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[20]
port 79 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[21]
port 80 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[22]
port 81 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 chany_bottom_in[23]
port 82 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[24]
port 83 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[25]
port 84 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 chany_bottom_in[26]
port 85 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_in[27]
port 86 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 chany_bottom_in[28]
port 87 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[29]
port 88 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 chany_bottom_in[2]
port 89 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_in[3]
port 90 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_in[4]
port 91 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_in[5]
port 92 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[6]
port 93 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[7]
port 94 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 chany_bottom_in[8]
port 95 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[9]
port 96 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[0]
port 97 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[10]
port 98 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 chany_bottom_out[11]
port 99 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 chany_bottom_out[12]
port 100 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[13]
port 101 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 chany_bottom_out[14]
port 102 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[15]
port 103 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[16]
port 104 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[17]
port 105 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[18]
port 106 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 chany_bottom_out[19]
port 107 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[1]
port 108 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 chany_bottom_out[20]
port 109 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[21]
port 110 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[22]
port 111 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 chany_bottom_out[23]
port 112 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[24]
port 113 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 chany_bottom_out[25]
port 114 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 chany_bottom_out[26]
port 115 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 chany_bottom_out[27]
port 116 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 chany_bottom_out[28]
port 117 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 chany_bottom_out[29]
port 118 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_out[2]
port 119 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_out[3]
port 120 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 chany_bottom_out[4]
port 121 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[5]
port 122 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_out[6]
port 123 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 chany_bottom_out[7]
port 124 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[8]
port 125 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[9]
port 126 nsew signal output
rlabel metal2 s 12898 56200 12954 57000 6 chany_top_in_0[0]
port 127 nsew signal input
rlabel metal2 s 16578 56200 16634 57000 6 chany_top_in_0[10]
port 128 nsew signal input
rlabel metal2 s 16946 56200 17002 57000 6 chany_top_in_0[11]
port 129 nsew signal input
rlabel metal2 s 17314 56200 17370 57000 6 chany_top_in_0[12]
port 130 nsew signal input
rlabel metal2 s 17682 56200 17738 57000 6 chany_top_in_0[13]
port 131 nsew signal input
rlabel metal2 s 18050 56200 18106 57000 6 chany_top_in_0[14]
port 132 nsew signal input
rlabel metal2 s 18418 56200 18474 57000 6 chany_top_in_0[15]
port 133 nsew signal input
rlabel metal2 s 18786 56200 18842 57000 6 chany_top_in_0[16]
port 134 nsew signal input
rlabel metal2 s 19154 56200 19210 57000 6 chany_top_in_0[17]
port 135 nsew signal input
rlabel metal2 s 19522 56200 19578 57000 6 chany_top_in_0[18]
port 136 nsew signal input
rlabel metal2 s 19890 56200 19946 57000 6 chany_top_in_0[19]
port 137 nsew signal input
rlabel metal2 s 13266 56200 13322 57000 6 chany_top_in_0[1]
port 138 nsew signal input
rlabel metal2 s 20258 56200 20314 57000 6 chany_top_in_0[20]
port 139 nsew signal input
rlabel metal2 s 20626 56200 20682 57000 6 chany_top_in_0[21]
port 140 nsew signal input
rlabel metal2 s 20994 56200 21050 57000 6 chany_top_in_0[22]
port 141 nsew signal input
rlabel metal2 s 21362 56200 21418 57000 6 chany_top_in_0[23]
port 142 nsew signal input
rlabel metal2 s 21730 56200 21786 57000 6 chany_top_in_0[24]
port 143 nsew signal input
rlabel metal2 s 22098 56200 22154 57000 6 chany_top_in_0[25]
port 144 nsew signal input
rlabel metal2 s 22466 56200 22522 57000 6 chany_top_in_0[26]
port 145 nsew signal input
rlabel metal2 s 22834 56200 22890 57000 6 chany_top_in_0[27]
port 146 nsew signal input
rlabel metal2 s 23202 56200 23258 57000 6 chany_top_in_0[28]
port 147 nsew signal input
rlabel metal2 s 23570 56200 23626 57000 6 chany_top_in_0[29]
port 148 nsew signal input
rlabel metal2 s 13634 56200 13690 57000 6 chany_top_in_0[2]
port 149 nsew signal input
rlabel metal2 s 14002 56200 14058 57000 6 chany_top_in_0[3]
port 150 nsew signal input
rlabel metal2 s 14370 56200 14426 57000 6 chany_top_in_0[4]
port 151 nsew signal input
rlabel metal2 s 14738 56200 14794 57000 6 chany_top_in_0[5]
port 152 nsew signal input
rlabel metal2 s 15106 56200 15162 57000 6 chany_top_in_0[6]
port 153 nsew signal input
rlabel metal2 s 15474 56200 15530 57000 6 chany_top_in_0[7]
port 154 nsew signal input
rlabel metal2 s 15842 56200 15898 57000 6 chany_top_in_0[8]
port 155 nsew signal input
rlabel metal2 s 16210 56200 16266 57000 6 chany_top_in_0[9]
port 156 nsew signal input
rlabel metal2 s 1858 56200 1914 57000 6 chany_top_out_0[0]
port 157 nsew signal output
rlabel metal2 s 5538 56200 5594 57000 6 chany_top_out_0[10]
port 158 nsew signal output
rlabel metal2 s 5906 56200 5962 57000 6 chany_top_out_0[11]
port 159 nsew signal output
rlabel metal2 s 6274 56200 6330 57000 6 chany_top_out_0[12]
port 160 nsew signal output
rlabel metal2 s 6642 56200 6698 57000 6 chany_top_out_0[13]
port 161 nsew signal output
rlabel metal2 s 7010 56200 7066 57000 6 chany_top_out_0[14]
port 162 nsew signal output
rlabel metal2 s 7378 56200 7434 57000 6 chany_top_out_0[15]
port 163 nsew signal output
rlabel metal2 s 7746 56200 7802 57000 6 chany_top_out_0[16]
port 164 nsew signal output
rlabel metal2 s 8114 56200 8170 57000 6 chany_top_out_0[17]
port 165 nsew signal output
rlabel metal2 s 8482 56200 8538 57000 6 chany_top_out_0[18]
port 166 nsew signal output
rlabel metal2 s 8850 56200 8906 57000 6 chany_top_out_0[19]
port 167 nsew signal output
rlabel metal2 s 2226 56200 2282 57000 6 chany_top_out_0[1]
port 168 nsew signal output
rlabel metal2 s 9218 56200 9274 57000 6 chany_top_out_0[20]
port 169 nsew signal output
rlabel metal2 s 9586 56200 9642 57000 6 chany_top_out_0[21]
port 170 nsew signal output
rlabel metal2 s 9954 56200 10010 57000 6 chany_top_out_0[22]
port 171 nsew signal output
rlabel metal2 s 10322 56200 10378 57000 6 chany_top_out_0[23]
port 172 nsew signal output
rlabel metal2 s 10690 56200 10746 57000 6 chany_top_out_0[24]
port 173 nsew signal output
rlabel metal2 s 11058 56200 11114 57000 6 chany_top_out_0[25]
port 174 nsew signal output
rlabel metal2 s 11426 56200 11482 57000 6 chany_top_out_0[26]
port 175 nsew signal output
rlabel metal2 s 11794 56200 11850 57000 6 chany_top_out_0[27]
port 176 nsew signal output
rlabel metal2 s 12162 56200 12218 57000 6 chany_top_out_0[28]
port 177 nsew signal output
rlabel metal2 s 12530 56200 12586 57000 6 chany_top_out_0[29]
port 178 nsew signal output
rlabel metal2 s 2594 56200 2650 57000 6 chany_top_out_0[2]
port 179 nsew signal output
rlabel metal2 s 2962 56200 3018 57000 6 chany_top_out_0[3]
port 180 nsew signal output
rlabel metal2 s 3330 56200 3386 57000 6 chany_top_out_0[4]
port 181 nsew signal output
rlabel metal2 s 3698 56200 3754 57000 6 chany_top_out_0[5]
port 182 nsew signal output
rlabel metal2 s 4066 56200 4122 57000 6 chany_top_out_0[6]
port 183 nsew signal output
rlabel metal2 s 4434 56200 4490 57000 6 chany_top_out_0[7]
port 184 nsew signal output
rlabel metal2 s 4802 56200 4858 57000 6 chany_top_out_0[8]
port 185 nsew signal output
rlabel metal2 s 5170 56200 5226 57000 6 chany_top_out_0[9]
port 186 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 gfpga_pad_io_soc_dir[0]
port 187 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 gfpga_pad_io_soc_dir[1]
port 188 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 gfpga_pad_io_soc_dir[2]
port 189 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 gfpga_pad_io_soc_dir[3]
port 190 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 gfpga_pad_io_soc_in[0]
port 191 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 gfpga_pad_io_soc_in[1]
port 192 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 gfpga_pad_io_soc_in[2]
port 193 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 gfpga_pad_io_soc_in[3]
port 194 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 gfpga_pad_io_soc_out[0]
port 195 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 gfpga_pad_io_soc_out[1]
port 196 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 gfpga_pad_io_soc_out[2]
port 197 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 gfpga_pad_io_soc_out[3]
port 198 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 isol_n
port 199 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 prog_clk
port 200 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 prog_reset
port 201 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 reset
port 202 nsew signal input
rlabel metal3 s 26200 50464 27000 50584 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 203 nsew signal input
rlabel metal3 s 26200 51280 27000 51400 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 204 nsew signal input
rlabel metal3 s 26200 52096 27000 52216 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 205 nsew signal input
rlabel metal3 s 26200 52912 27000 53032 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 206 nsew signal input
rlabel metal3 s 26200 53728 27000 53848 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 207 nsew signal input
rlabel metal3 s 26200 54544 27000 54664 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 208 nsew signal input
rlabel metal3 s 26200 55360 27000 55480 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 209 nsew signal input
rlabel metal3 s 26200 56176 27000 56296 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 210 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 right_width_0_height_0_subtile_0__pin_inpad_0_
port 211 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 right_width_0_height_0_subtile_1__pin_inpad_0_
port 212 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 right_width_0_height_0_subtile_2__pin_inpad_0_
port 213 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 right_width_0_height_0_subtile_3__pin_inpad_0_
port 214 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 test_enable
port 215 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 216 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 217 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 218 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 219 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 27000 57000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3033730
string GDS_FILE /home/hosni/OpenFPGA/erc-fixes/clear/openlane/left_tile/runs/23_04_26_18_01/results/signoff/left_tile.magic.gds
string GDS_START 183514
<< end >>

