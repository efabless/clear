magic
tech sky130A
magscale 1 2
timestamp 1656242434
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 1104 1640 22802 20720
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20902 0 20958 800
<< obsm2 >>
rect 1490 22144 5666 22200
rect 5834 22144 17166 22200
rect 17334 22144 22796 22200
rect 1490 856 22796 22144
rect 1490 734 1986 856
rect 2154 734 2446 856
rect 2614 734 2906 856
rect 3074 734 3366 856
rect 3534 734 3826 856
rect 3994 734 4286 856
rect 4454 734 4746 856
rect 4914 734 5206 856
rect 5374 734 5666 856
rect 5834 734 6126 856
rect 6294 734 6586 856
rect 6754 734 7046 856
rect 7214 734 7506 856
rect 7674 734 7966 856
rect 8134 734 8426 856
rect 8594 734 8886 856
rect 9054 734 9346 856
rect 9514 734 9806 856
rect 9974 734 10266 856
rect 10434 734 10726 856
rect 10894 734 11186 856
rect 11354 734 11646 856
rect 11814 734 12106 856
rect 12274 734 12566 856
rect 12734 734 13026 856
rect 13194 734 13486 856
rect 13654 734 13946 856
rect 14114 734 14406 856
rect 14574 734 14866 856
rect 15034 734 15326 856
rect 15494 734 15786 856
rect 15954 734 16246 856
rect 16414 734 16706 856
rect 16874 734 17166 856
rect 17334 734 17626 856
rect 17794 734 18086 856
rect 18254 734 18546 856
rect 18714 734 19006 856
rect 19174 734 19466 856
rect 19634 734 19926 856
rect 20094 734 20386 856
rect 20554 734 20846 856
rect 21014 734 22796 856
<< metal3 >>
rect 22200 21360 23000 21480
rect 22200 20952 23000 21072
rect 22200 20544 23000 20664
rect 22200 20136 23000 20256
rect 22200 19728 23000 19848
rect 22200 19320 23000 19440
rect 22200 18912 23000 19032
rect 22200 18504 23000 18624
rect 22200 18096 23000 18216
rect 22200 17688 23000 17808
rect 22200 17280 23000 17400
rect 22200 16872 23000 16992
rect 22200 16464 23000 16584
rect 22200 16056 23000 16176
rect 22200 15648 23000 15768
rect 22200 15240 23000 15360
rect 22200 14832 23000 14952
rect 22200 14424 23000 14544
rect 22200 14016 23000 14136
rect 22200 13608 23000 13728
rect 22200 13200 23000 13320
rect 22200 12792 23000 12912
rect 22200 12384 23000 12504
rect 22200 11976 23000 12096
rect 0 11432 800 11552
rect 22200 11568 23000 11688
rect 22200 11160 23000 11280
rect 22200 10752 23000 10872
rect 22200 10344 23000 10464
rect 22200 9936 23000 10056
rect 22200 9528 23000 9648
rect 22200 9120 23000 9240
rect 22200 8712 23000 8832
rect 22200 8304 23000 8424
rect 22200 7896 23000 8016
rect 22200 7488 23000 7608
rect 22200 7080 23000 7200
rect 22200 6672 23000 6792
rect 22200 6264 23000 6384
rect 22200 5856 23000 5976
rect 22200 5448 23000 5568
rect 22200 5040 23000 5160
rect 22200 4632 23000 4752
rect 22200 4224 23000 4344
rect 22200 3816 23000 3936
rect 22200 3408 23000 3528
rect 22200 3000 23000 3120
rect 22200 2592 23000 2712
rect 22200 2184 23000 2304
rect 22200 1776 23000 1896
rect 22200 1368 23000 1488
<< obsm3 >>
rect 800 21280 22120 21453
rect 800 21152 22202 21280
rect 800 20872 22120 21152
rect 800 20744 22202 20872
rect 800 20464 22120 20744
rect 800 20336 22202 20464
rect 800 20056 22120 20336
rect 800 19928 22202 20056
rect 800 19648 22120 19928
rect 800 19520 22202 19648
rect 800 19240 22120 19520
rect 800 19112 22202 19240
rect 800 18832 22120 19112
rect 800 18704 22202 18832
rect 800 18424 22120 18704
rect 800 18296 22202 18424
rect 800 18016 22120 18296
rect 800 17888 22202 18016
rect 800 17608 22120 17888
rect 800 17480 22202 17608
rect 800 17200 22120 17480
rect 800 17072 22202 17200
rect 800 16792 22120 17072
rect 800 16664 22202 16792
rect 800 16384 22120 16664
rect 800 16256 22202 16384
rect 800 15976 22120 16256
rect 800 15848 22202 15976
rect 800 15568 22120 15848
rect 800 15440 22202 15568
rect 800 15160 22120 15440
rect 800 15032 22202 15160
rect 800 14752 22120 15032
rect 800 14624 22202 14752
rect 800 14344 22120 14624
rect 800 14216 22202 14344
rect 800 13936 22120 14216
rect 800 13808 22202 13936
rect 800 13528 22120 13808
rect 800 13400 22202 13528
rect 800 13120 22120 13400
rect 800 12992 22202 13120
rect 800 12712 22120 12992
rect 800 12584 22202 12712
rect 800 12304 22120 12584
rect 800 12176 22202 12304
rect 800 11896 22120 12176
rect 800 11768 22202 11896
rect 800 11632 22120 11768
rect 880 11488 22120 11632
rect 880 11360 22202 11488
rect 880 11352 22120 11360
rect 800 11080 22120 11352
rect 800 10952 22202 11080
rect 800 10672 22120 10952
rect 800 10544 22202 10672
rect 800 10264 22120 10544
rect 800 10136 22202 10264
rect 800 9856 22120 10136
rect 800 9728 22202 9856
rect 800 9448 22120 9728
rect 800 9320 22202 9448
rect 800 9040 22120 9320
rect 800 8912 22202 9040
rect 800 8632 22120 8912
rect 800 8504 22202 8632
rect 800 8224 22120 8504
rect 800 8096 22202 8224
rect 800 7816 22120 8096
rect 800 7688 22202 7816
rect 800 7408 22120 7688
rect 800 7280 22202 7408
rect 800 7000 22120 7280
rect 800 6872 22202 7000
rect 800 6592 22120 6872
rect 800 6464 22202 6592
rect 800 6184 22120 6464
rect 800 6056 22202 6184
rect 800 5776 22120 6056
rect 800 5648 22202 5776
rect 800 5368 22120 5648
rect 800 5240 22202 5368
rect 800 4960 22120 5240
rect 800 4832 22202 4960
rect 800 4552 22120 4832
rect 800 4424 22202 4552
rect 800 4144 22120 4424
rect 800 4016 22202 4144
rect 800 3736 22120 4016
rect 800 3608 22202 3736
rect 800 3328 22120 3608
rect 800 3200 22202 3328
rect 800 2920 22120 3200
rect 800 2792 22202 2920
rect 800 2512 22120 2792
rect 800 2384 22202 2512
rect 800 2104 22120 2384
rect 800 1976 22202 2104
rect 800 1696 22120 1976
rect 800 1568 22202 1696
rect 800 1395 22120 1568
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 17355 3571 19057 16013
<< labels >>
rlabel metal2 s 5722 22200 5778 23000 6 SC_IN_TOP
port 1 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 SC_OUT_BOT
port 2 nsew signal output
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal2 s 2042 0 2098 800 6 bottom_left_grid_pin_1_
port 5 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_head
port 6 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 ccff_tail
port 7 nsew signal output
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[0]
port 8 nsew signal input
rlabel metal3 s 22200 8712 23000 8832 6 chanx_right_in[10]
port 9 nsew signal input
rlabel metal3 s 22200 9120 23000 9240 6 chanx_right_in[11]
port 10 nsew signal input
rlabel metal3 s 22200 9528 23000 9648 6 chanx_right_in[12]
port 11 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 12 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 13 nsew signal input
rlabel metal3 s 22200 10752 23000 10872 6 chanx_right_in[15]
port 14 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[16]
port 15 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[17]
port 16 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[18]
port 17 nsew signal input
rlabel metal3 s 22200 12384 23000 12504 6 chanx_right_in[19]
port 18 nsew signal input
rlabel metal3 s 22200 5040 23000 5160 6 chanx_right_in[1]
port 19 nsew signal input
rlabel metal3 s 22200 5448 23000 5568 6 chanx_right_in[2]
port 20 nsew signal input
rlabel metal3 s 22200 5856 23000 5976 6 chanx_right_in[3]
port 21 nsew signal input
rlabel metal3 s 22200 6264 23000 6384 6 chanx_right_in[4]
port 22 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[5]
port 23 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[6]
port 24 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[7]
port 25 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[8]
port 26 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[9]
port 27 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_out[0]
port 28 nsew signal output
rlabel metal3 s 22200 16872 23000 16992 6 chanx_right_out[10]
port 29 nsew signal output
rlabel metal3 s 22200 17280 23000 17400 6 chanx_right_out[11]
port 30 nsew signal output
rlabel metal3 s 22200 17688 23000 17808 6 chanx_right_out[12]
port 31 nsew signal output
rlabel metal3 s 22200 18096 23000 18216 6 chanx_right_out[13]
port 32 nsew signal output
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[14]
port 33 nsew signal output
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[15]
port 34 nsew signal output
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[16]
port 35 nsew signal output
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[17]
port 36 nsew signal output
rlabel metal3 s 22200 20136 23000 20256 6 chanx_right_out[18]
port 37 nsew signal output
rlabel metal3 s 22200 20544 23000 20664 6 chanx_right_out[19]
port 38 nsew signal output
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[1]
port 39 nsew signal output
rlabel metal3 s 22200 13608 23000 13728 6 chanx_right_out[2]
port 40 nsew signal output
rlabel metal3 s 22200 14016 23000 14136 6 chanx_right_out[3]
port 41 nsew signal output
rlabel metal3 s 22200 14424 23000 14544 6 chanx_right_out[4]
port 42 nsew signal output
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[5]
port 43 nsew signal output
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[6]
port 44 nsew signal output
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[7]
port 45 nsew signal output
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[8]
port 46 nsew signal output
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[9]
port 47 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_in[0]
port 48 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 chany_bottom_in[10]
port 49 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[11]
port 50 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_in[12]
port 51 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[13]
port 52 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[14]
port 53 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[15]
port 54 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 chany_bottom_in[16]
port 55 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[17]
port 56 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 chany_bottom_in[18]
port 57 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 chany_bottom_in[19]
port 58 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 chany_bottom_in[1]
port 59 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_in[2]
port 60 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[3]
port 61 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[4]
port 62 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_in[5]
port 63 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_in[6]
port 64 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_in[7]
port 65 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_in[8]
port 66 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[9]
port 67 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_out[0]
port 68 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 chany_bottom_out[10]
port 69 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 chany_bottom_out[11]
port 70 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 chany_bottom_out[12]
port 71 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[13]
port 72 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 chany_bottom_out[14]
port 73 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[15]
port 74 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 chany_bottom_out[16]
port 75 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[17]
port 76 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 chany_bottom_out[18]
port 77 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[19]
port 78 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_out[1]
port 79 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_out[2]
port 80 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[3]
port 81 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_out[4]
port 82 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[5]
port 83 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 chany_bottom_out[6]
port 84 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_out[7]
port 85 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 chany_bottom_out[8]
port 86 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[9]
port 87 nsew signal output
rlabel metal3 s 22200 20952 23000 21072 6 prog_clk_0_E_in
port 88 nsew signal input
rlabel metal3 s 22200 1368 23000 1488 6 right_bottom_grid_pin_34_
port 89 nsew signal input
rlabel metal3 s 22200 1776 23000 1896 6 right_bottom_grid_pin_35_
port 90 nsew signal input
rlabel metal3 s 22200 2184 23000 2304 6 right_bottom_grid_pin_36_
port 91 nsew signal input
rlabel metal3 s 22200 2592 23000 2712 6 right_bottom_grid_pin_37_
port 92 nsew signal input
rlabel metal3 s 22200 3000 23000 3120 6 right_bottom_grid_pin_38_
port 93 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_39_
port 94 nsew signal input
rlabel metal3 s 22200 3816 23000 3936 6 right_bottom_grid_pin_40_
port 95 nsew signal input
rlabel metal3 s 22200 4224 23000 4344 6 right_bottom_grid_pin_41_
port 96 nsew signal input
rlabel metal3 s 22200 21360 23000 21480 6 right_top_grid_pin_1_
port 97 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 933860
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_0__2_/runs/sb_0__2_/results/signoff/sb_0__2_.magic.gds
string GDS_START 75876
<< end >>

