VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 115.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 30.710 10.640 32.310 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.700 10.640 58.300 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.690 10.640 84.290 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.680 10.640 110.280 103.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.715 10.640 19.315 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.705 10.640 45.305 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.695 10.640 71.295 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.685 10.640 97.285 103.600 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 25.200 115.000 25.800 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 45.600 115.000 46.200 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 47.640 115.000 48.240 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 49.680 115.000 50.280 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 51.720 115.000 52.320 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 53.760 115.000 54.360 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 55.800 115.000 56.400 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 57.840 115.000 58.440 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 59.880 115.000 60.480 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 61.920 115.000 62.520 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 63.960 115.000 64.560 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 27.240 115.000 27.840 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 29.280 115.000 29.880 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 31.320 115.000 31.920 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 33.360 115.000 33.960 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 35.400 115.000 36.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 37.440 115.000 38.040 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 39.480 115.000 40.080 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 41.520 115.000 42.120 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 43.560 115.000 44.160 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 66.000 115.000 66.600 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 86.400 115.000 87.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 88.440 115.000 89.040 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 90.480 115.000 91.080 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 92.520 115.000 93.120 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 94.560 115.000 95.160 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 96.600 115.000 97.200 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 98.640 115.000 99.240 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 100.680 115.000 101.280 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 102.720 115.000 103.320 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 104.760 115.000 105.360 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 68.040 115.000 68.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 70.080 115.000 70.680 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 72.120 115.000 72.720 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 74.160 115.000 74.760 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 76.200 115.000 76.800 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 78.240 115.000 78.840 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 80.280 115.000 80.880 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 82.320 115.000 82.920 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 84.360 115.000 84.960 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 111.000 4.970 115.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 111.000 32.570 115.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 111.000 35.330 115.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 111.000 38.090 115.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 111.000 40.850 115.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 111.000 43.610 115.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 111.000 46.370 115.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 111.000 49.130 115.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 111.000 51.890 115.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 111.000 54.650 115.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 111.000 57.410 115.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 111.000 7.730 115.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 111.000 10.490 115.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 111.000 13.250 115.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 111.000 16.010 115.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 111.000 18.770 115.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 111.000 21.530 115.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 111.000 24.290 115.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 111.000 27.050 115.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 111.000 29.810 115.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 111.000 60.170 115.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 111.000 87.770 115.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 111.000 90.530 115.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 111.000 93.290 115.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 111.000 96.050 115.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 111.000 98.810 115.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 111.000 101.570 115.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 111.000 104.330 115.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 111.000 107.090 115.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 111.000 109.850 115.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 111.000 112.610 115.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 111.000 62.930 115.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 111.000 65.690 115.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 111.000 68.450 115.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 111.000 71.210 115.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 111.000 73.970 115.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 111.000 76.730 115.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 111.000 79.490 115.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 111.000 82.250 115.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 111.000 85.010 115.000 ;
    END
  END chany_top_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 106.800 115.000 107.400 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 17.040 115.000 17.640 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 19.080 115.000 19.680 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 21.120 115.000 21.720 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 23.160 115.000 23.760 ;
    END
  END right_bottom_grid_pin_17_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 6.840 115.000 7.440 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 8.880 115.000 9.480 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 10.920 115.000 11.520 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 12.960 115.000 13.560 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 15.000 115.000 15.600 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 111.000 2.210 115.000 ;
    END
  END top_left_grid_pin_1_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 109.480 103.445 ;
      LAYER met1 ;
        RECT 1.910 10.640 112.630 103.600 ;
      LAYER met2 ;
        RECT 2.490 110.720 4.410 111.250 ;
        RECT 5.250 110.720 7.170 111.250 ;
        RECT 8.010 110.720 9.930 111.250 ;
        RECT 10.770 110.720 12.690 111.250 ;
        RECT 13.530 110.720 15.450 111.250 ;
        RECT 16.290 110.720 18.210 111.250 ;
        RECT 19.050 110.720 20.970 111.250 ;
        RECT 21.810 110.720 23.730 111.250 ;
        RECT 24.570 110.720 26.490 111.250 ;
        RECT 27.330 110.720 29.250 111.250 ;
        RECT 30.090 110.720 32.010 111.250 ;
        RECT 32.850 110.720 34.770 111.250 ;
        RECT 35.610 110.720 37.530 111.250 ;
        RECT 38.370 110.720 40.290 111.250 ;
        RECT 41.130 110.720 43.050 111.250 ;
        RECT 43.890 110.720 45.810 111.250 ;
        RECT 46.650 110.720 48.570 111.250 ;
        RECT 49.410 110.720 51.330 111.250 ;
        RECT 52.170 110.720 54.090 111.250 ;
        RECT 54.930 110.720 56.850 111.250 ;
        RECT 57.690 110.720 59.610 111.250 ;
        RECT 60.450 110.720 62.370 111.250 ;
        RECT 63.210 110.720 65.130 111.250 ;
        RECT 65.970 110.720 67.890 111.250 ;
        RECT 68.730 110.720 70.650 111.250 ;
        RECT 71.490 110.720 73.410 111.250 ;
        RECT 74.250 110.720 76.170 111.250 ;
        RECT 77.010 110.720 78.930 111.250 ;
        RECT 79.770 110.720 81.690 111.250 ;
        RECT 82.530 110.720 84.450 111.250 ;
        RECT 85.290 110.720 87.210 111.250 ;
        RECT 88.050 110.720 89.970 111.250 ;
        RECT 90.810 110.720 92.730 111.250 ;
        RECT 93.570 110.720 95.490 111.250 ;
        RECT 96.330 110.720 98.250 111.250 ;
        RECT 99.090 110.720 101.010 111.250 ;
        RECT 101.850 110.720 103.770 111.250 ;
        RECT 104.610 110.720 106.530 111.250 ;
        RECT 107.370 110.720 109.290 111.250 ;
        RECT 110.130 110.720 112.050 111.250 ;
        RECT 1.940 6.955 112.600 110.720 ;
      LAYER met3 ;
        RECT 4.000 106.400 110.600 107.265 ;
        RECT 4.000 105.760 111.010 106.400 ;
        RECT 4.000 104.360 110.600 105.760 ;
        RECT 4.000 103.720 111.010 104.360 ;
        RECT 4.000 102.320 110.600 103.720 ;
        RECT 4.000 101.680 111.010 102.320 ;
        RECT 4.000 100.280 110.600 101.680 ;
        RECT 4.000 99.640 111.010 100.280 ;
        RECT 4.000 98.240 110.600 99.640 ;
        RECT 4.000 97.600 111.010 98.240 ;
        RECT 4.000 96.200 110.600 97.600 ;
        RECT 4.000 95.560 111.010 96.200 ;
        RECT 4.000 94.160 110.600 95.560 ;
        RECT 4.000 93.520 111.010 94.160 ;
        RECT 4.000 92.120 110.600 93.520 ;
        RECT 4.000 91.480 111.010 92.120 ;
        RECT 4.000 90.080 110.600 91.480 ;
        RECT 4.000 89.440 111.010 90.080 ;
        RECT 4.000 88.040 110.600 89.440 ;
        RECT 4.000 87.400 111.010 88.040 ;
        RECT 4.000 86.720 110.600 87.400 ;
        RECT 4.400 86.000 110.600 86.720 ;
        RECT 4.400 85.360 111.010 86.000 ;
        RECT 4.400 85.320 110.600 85.360 ;
        RECT 4.000 83.960 110.600 85.320 ;
        RECT 4.000 83.320 111.010 83.960 ;
        RECT 4.000 81.920 110.600 83.320 ;
        RECT 4.000 81.280 111.010 81.920 ;
        RECT 4.000 79.880 110.600 81.280 ;
        RECT 4.000 79.240 111.010 79.880 ;
        RECT 4.000 77.840 110.600 79.240 ;
        RECT 4.000 77.200 111.010 77.840 ;
        RECT 4.000 75.800 110.600 77.200 ;
        RECT 4.000 75.160 111.010 75.800 ;
        RECT 4.000 73.760 110.600 75.160 ;
        RECT 4.000 73.120 111.010 73.760 ;
        RECT 4.000 71.720 110.600 73.120 ;
        RECT 4.000 71.080 111.010 71.720 ;
        RECT 4.000 69.680 110.600 71.080 ;
        RECT 4.000 69.040 111.010 69.680 ;
        RECT 4.000 67.640 110.600 69.040 ;
        RECT 4.000 67.000 111.010 67.640 ;
        RECT 4.000 65.600 110.600 67.000 ;
        RECT 4.000 64.960 111.010 65.600 ;
        RECT 4.000 63.560 110.600 64.960 ;
        RECT 4.000 62.920 111.010 63.560 ;
        RECT 4.000 61.520 110.600 62.920 ;
        RECT 4.000 60.880 111.010 61.520 ;
        RECT 4.000 59.480 110.600 60.880 ;
        RECT 4.000 58.840 111.010 59.480 ;
        RECT 4.000 57.440 110.600 58.840 ;
        RECT 4.000 56.800 111.010 57.440 ;
        RECT 4.000 55.400 110.600 56.800 ;
        RECT 4.000 54.760 111.010 55.400 ;
        RECT 4.000 53.360 110.600 54.760 ;
        RECT 4.000 52.720 111.010 53.360 ;
        RECT 4.000 51.320 110.600 52.720 ;
        RECT 4.000 50.680 111.010 51.320 ;
        RECT 4.000 49.280 110.600 50.680 ;
        RECT 4.000 48.640 111.010 49.280 ;
        RECT 4.000 47.240 110.600 48.640 ;
        RECT 4.000 46.600 111.010 47.240 ;
        RECT 4.000 45.200 110.600 46.600 ;
        RECT 4.000 44.560 111.010 45.200 ;
        RECT 4.000 43.160 110.600 44.560 ;
        RECT 4.000 42.520 111.010 43.160 ;
        RECT 4.000 41.120 110.600 42.520 ;
        RECT 4.000 40.480 111.010 41.120 ;
        RECT 4.000 39.080 110.600 40.480 ;
        RECT 4.000 38.440 111.010 39.080 ;
        RECT 4.000 37.040 110.600 38.440 ;
        RECT 4.000 36.400 111.010 37.040 ;
        RECT 4.000 35.000 110.600 36.400 ;
        RECT 4.000 34.360 111.010 35.000 ;
        RECT 4.000 32.960 110.600 34.360 ;
        RECT 4.000 32.320 111.010 32.960 ;
        RECT 4.000 30.920 110.600 32.320 ;
        RECT 4.000 30.280 111.010 30.920 ;
        RECT 4.000 29.600 110.600 30.280 ;
        RECT 4.400 28.880 110.600 29.600 ;
        RECT 4.400 28.240 111.010 28.880 ;
        RECT 4.400 28.200 110.600 28.240 ;
        RECT 4.000 26.840 110.600 28.200 ;
        RECT 4.000 26.200 111.010 26.840 ;
        RECT 4.000 24.800 110.600 26.200 ;
        RECT 4.000 24.160 111.010 24.800 ;
        RECT 4.000 22.760 110.600 24.160 ;
        RECT 4.000 22.120 111.010 22.760 ;
        RECT 4.000 20.720 110.600 22.120 ;
        RECT 4.000 20.080 111.010 20.720 ;
        RECT 4.000 18.680 110.600 20.080 ;
        RECT 4.000 18.040 111.010 18.680 ;
        RECT 4.000 16.640 110.600 18.040 ;
        RECT 4.000 16.000 111.010 16.640 ;
        RECT 4.000 14.600 110.600 16.000 ;
        RECT 4.000 13.960 111.010 14.600 ;
        RECT 4.000 12.560 110.600 13.960 ;
        RECT 4.000 11.920 111.010 12.560 ;
        RECT 4.000 10.520 110.600 11.920 ;
        RECT 4.000 9.880 111.010 10.520 ;
        RECT 4.000 8.480 110.600 9.880 ;
        RECT 4.000 7.840 111.010 8.480 ;
        RECT 4.000 6.975 110.600 7.840 ;
      LAYER met4 ;
        RECT 97.815 66.135 98.145 90.265 ;
  END
END sb_0__0_
END LIBRARY

