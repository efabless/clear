magic
tech sky130A
magscale 1 2
timestamp 1679320553
<< viali >>
rect 23213 54281 23247 54315
rect 24869 54281 24903 54315
rect 46121 54281 46155 54315
rect 3249 54213 3283 54247
rect 8401 54213 8435 54247
rect 10701 54213 10735 54247
rect 13553 54213 13587 54247
rect 15853 54213 15887 54247
rect 18705 54213 18739 54247
rect 42625 54213 42659 54247
rect 46029 54213 46063 54247
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9965 54145 9999 54179
rect 12541 54145 12575 54179
rect 15025 54145 15059 54179
rect 17693 54145 17727 54179
rect 20177 54145 20211 54179
rect 22753 54145 22787 54179
rect 23397 54145 23431 54179
rect 24041 54145 24075 54179
rect 25053 54145 25087 54179
rect 25697 54145 25731 54179
rect 26341 54145 26375 54179
rect 27353 54145 27387 54179
rect 27997 54145 28031 54179
rect 28641 54145 28675 54179
rect 29929 54145 29963 54179
rect 30573 54145 30607 54179
rect 31217 54145 31251 54179
rect 32505 54145 32539 54179
rect 33149 54145 33183 54179
rect 33793 54145 33827 54179
rect 35173 54145 35207 54179
rect 36645 54145 36679 54179
rect 37657 54145 37691 54179
rect 38301 54145 38335 54179
rect 38945 54145 38979 54179
rect 40233 54145 40267 54179
rect 40877 54145 40911 54179
rect 45201 54145 45235 54179
rect 46857 54145 46891 54179
rect 47777 54145 47811 54179
rect 48513 54145 48547 54179
rect 5457 54077 5491 54111
rect 20545 54077 20579 54111
rect 35449 54077 35483 54111
rect 23857 54009 23891 54043
rect 26157 54009 26191 54043
rect 28457 54009 28491 54043
rect 38117 54009 38151 54043
rect 38761 54009 38795 54043
rect 40049 54009 40083 54043
rect 40693 54009 40727 54043
rect 45385 54009 45419 54043
rect 47041 54009 47075 54043
rect 47961 54009 47995 54043
rect 22569 53941 22603 53975
rect 25513 53941 25547 53975
rect 27169 53941 27203 53975
rect 27813 53941 27847 53975
rect 29745 53941 29779 53975
rect 30389 53941 30423 53975
rect 31033 53941 31067 53975
rect 32321 53941 32355 53975
rect 32965 53941 32999 53975
rect 33609 53941 33643 53975
rect 36461 53941 36495 53975
rect 37473 53941 37507 53975
rect 43913 53941 43947 53975
rect 48697 53941 48731 53975
rect 23581 53669 23615 53703
rect 36461 53669 36495 53703
rect 48237 53669 48271 53703
rect 2881 53601 2915 53635
rect 6101 53601 6135 53635
rect 7849 53601 7883 53635
rect 11253 53601 11287 53635
rect 13369 53601 13403 53635
rect 16405 53601 16439 53635
rect 18337 53601 18371 53635
rect 34897 53601 34931 53635
rect 44465 53601 44499 53635
rect 2053 53533 2087 53567
rect 5457 53533 5491 53567
rect 7389 53533 7423 53567
rect 10701 53533 10735 53567
rect 12541 53533 12575 53567
rect 15853 53533 15887 53567
rect 17693 53533 17727 53567
rect 21189 53533 21223 53567
rect 23029 53533 23063 53567
rect 23765 53533 23799 53567
rect 28917 53533 28951 53567
rect 31493 53533 31527 53567
rect 34069 53533 34103 53567
rect 35173 53533 35207 53567
rect 36645 53533 36679 53567
rect 39221 53533 39255 53567
rect 44281 53533 44315 53567
rect 46765 53533 46799 53567
rect 48053 53533 48087 53567
rect 48697 53533 48731 53567
rect 21925 53465 21959 53499
rect 22845 53397 22879 53431
rect 28733 53397 28767 53431
rect 31309 53397 31343 53431
rect 33885 53397 33919 53431
rect 39037 53397 39071 53431
rect 46949 53397 46983 53431
rect 48881 53397 48915 53431
rect 23305 53193 23339 53227
rect 24041 53193 24075 53227
rect 23213 53125 23247 53159
rect 47869 53125 47903 53159
rect 2513 53057 2547 53091
rect 4721 53057 4755 53091
rect 7021 53057 7055 53091
rect 7665 53057 7699 53091
rect 9873 53057 9907 53091
rect 12817 53057 12851 53091
rect 15025 53057 15059 53091
rect 17877 53057 17911 53091
rect 19901 53057 19935 53091
rect 22201 53057 22235 53091
rect 23949 53057 23983 53091
rect 48789 53057 48823 53091
rect 2789 52989 2823 53023
rect 5089 52989 5123 53023
rect 7941 52989 7975 53023
rect 10241 52989 10275 53023
rect 13093 52989 13127 53023
rect 15393 52989 15427 53023
rect 18245 52989 18279 53023
rect 20177 52989 20211 53023
rect 48513 52989 48547 53023
rect 6837 52921 6871 52955
rect 22017 52853 22051 52887
rect 47961 52853 47995 52887
rect 22569 52649 22603 52683
rect 23397 52649 23431 52683
rect 20269 52581 20303 52615
rect 2145 52513 2179 52547
rect 4813 52513 4847 52547
rect 7297 52513 7331 52547
rect 9873 52513 9907 52547
rect 12449 52513 12483 52547
rect 15025 52513 15059 52547
rect 17601 52513 17635 52547
rect 48789 52513 48823 52547
rect 1685 52445 1719 52479
rect 4445 52445 4479 52479
rect 7021 52445 7055 52479
rect 9597 52445 9631 52479
rect 12173 52445 12207 52479
rect 14749 52445 14783 52479
rect 17325 52445 17359 52479
rect 22753 52445 22787 52479
rect 48053 52445 48087 52479
rect 48513 52445 48547 52479
rect 20085 52377 20119 52411
rect 23305 52377 23339 52411
rect 8493 52105 8527 52139
rect 8401 51969 8435 52003
rect 49341 51969 49375 52003
rect 49157 51765 49191 51799
rect 9321 51561 9355 51595
rect 2053 51425 2087 51459
rect 41705 51425 41739 51459
rect 1777 51357 1811 51391
rect 41429 51357 41463 51391
rect 43453 51357 43487 51391
rect 48513 51357 48547 51391
rect 48789 51357 48823 51391
rect 9229 51289 9263 51323
rect 9321 51017 9355 51051
rect 10149 51017 10183 51051
rect 13461 51017 13495 51051
rect 17049 51017 17083 51051
rect 22201 51017 22235 51051
rect 26249 51017 26283 51051
rect 27353 51017 27387 51051
rect 31493 50949 31527 50983
rect 1777 50881 1811 50915
rect 9229 50881 9263 50915
rect 10057 50881 10091 50915
rect 13369 50881 13403 50915
rect 16957 50881 16991 50915
rect 22109 50881 22143 50915
rect 26433 50881 26467 50915
rect 27537 50881 27571 50915
rect 28273 50881 28307 50915
rect 31401 50881 31435 50915
rect 49341 50881 49375 50915
rect 2053 50813 2087 50847
rect 31585 50813 31619 50847
rect 28089 50745 28123 50779
rect 31033 50677 31067 50711
rect 49157 50677 49191 50711
rect 13461 50473 13495 50507
rect 17601 50473 17635 50507
rect 22661 50473 22695 50507
rect 31125 50473 31159 50507
rect 8401 50405 8435 50439
rect 16957 50405 16991 50439
rect 29929 50405 29963 50439
rect 28365 50337 28399 50371
rect 30481 50337 30515 50371
rect 31769 50337 31803 50371
rect 16773 50269 16807 50303
rect 28181 50269 28215 50303
rect 8217 50201 8251 50235
rect 13369 50201 13403 50235
rect 17509 50201 17543 50235
rect 22569 50201 22603 50235
rect 27813 50133 27847 50167
rect 28273 50133 28307 50167
rect 30297 50133 30331 50167
rect 30389 50133 30423 50167
rect 31493 50133 31527 50167
rect 31585 50133 31619 50167
rect 13277 49929 13311 49963
rect 14105 49929 14139 49963
rect 16221 49929 16255 49963
rect 22201 49929 22235 49963
rect 29837 49929 29871 49963
rect 31033 49929 31067 49963
rect 31493 49929 31527 49963
rect 32689 49929 32723 49963
rect 33517 49929 33551 49963
rect 33977 49929 34011 49963
rect 34713 49929 34747 49963
rect 35173 49929 35207 49963
rect 15117 49861 15151 49895
rect 21465 49861 21499 49895
rect 30205 49861 30239 49895
rect 31401 49861 31435 49895
rect 33885 49861 33919 49895
rect 1777 49793 1811 49827
rect 13461 49793 13495 49827
rect 14013 49793 14047 49827
rect 14933 49793 14967 49827
rect 16129 49793 16163 49827
rect 21281 49793 21315 49827
rect 22109 49793 22143 49827
rect 30297 49793 30331 49827
rect 35081 49793 35115 49827
rect 49341 49793 49375 49827
rect 2053 49725 2087 49759
rect 27629 49725 27663 49759
rect 30389 49725 30423 49759
rect 31585 49725 31619 49759
rect 32781 49725 32815 49759
rect 32873 49725 32907 49759
rect 34161 49725 34195 49759
rect 35357 49725 35391 49759
rect 32321 49657 32355 49691
rect 49157 49657 49191 49691
rect 27892 49589 27926 49623
rect 29377 49589 29411 49623
rect 10057 49385 10091 49419
rect 13461 49385 13495 49419
rect 19993 49385 20027 49419
rect 28825 49385 28859 49419
rect 33517 49385 33551 49419
rect 34897 49385 34931 49419
rect 27169 49317 27203 49351
rect 2053 49249 2087 49283
rect 28089 49249 28123 49283
rect 28181 49249 28215 49283
rect 30297 49249 30331 49283
rect 35449 49249 35483 49283
rect 1777 49181 1811 49215
rect 25421 49181 25455 49215
rect 29009 49181 29043 49215
rect 31769 49181 31803 49215
rect 49065 49181 49099 49215
rect 9965 49113 9999 49147
rect 13369 49113 13403 49147
rect 19901 49113 19935 49147
rect 25697 49113 25731 49147
rect 27997 49113 28031 49147
rect 30113 49113 30147 49147
rect 30205 49113 30239 49147
rect 32045 49113 32079 49147
rect 35265 49113 35299 49147
rect 27629 49045 27663 49079
rect 29745 49045 29779 49079
rect 35357 49045 35391 49079
rect 49249 49045 49283 49079
rect 25237 48841 25271 48875
rect 26341 48841 26375 48875
rect 27629 48841 27663 48875
rect 30849 48841 30883 48875
rect 34989 48841 35023 48875
rect 35081 48841 35115 48875
rect 24225 48773 24259 48807
rect 29653 48773 29687 48807
rect 32689 48773 32723 48807
rect 24133 48705 24167 48739
rect 25421 48705 25455 48739
rect 26249 48705 26283 48739
rect 27537 48705 27571 48739
rect 29561 48705 29595 48739
rect 30757 48705 30791 48739
rect 24317 48637 24351 48671
rect 26433 48637 26467 48671
rect 27721 48637 27755 48671
rect 29837 48637 29871 48671
rect 31033 48637 31067 48671
rect 32413 48637 32447 48671
rect 34161 48637 34195 48671
rect 35173 48637 35207 48671
rect 25881 48569 25915 48603
rect 29193 48569 29227 48603
rect 23765 48501 23799 48535
rect 27169 48501 27203 48535
rect 30389 48501 30423 48535
rect 34621 48501 34655 48535
rect 34897 48297 34931 48331
rect 33057 48229 33091 48263
rect 2053 48161 2087 48195
rect 20361 48161 20395 48195
rect 27077 48161 27111 48195
rect 31033 48161 31067 48195
rect 33517 48161 33551 48195
rect 33701 48161 33735 48195
rect 35449 48161 35483 48195
rect 36875 48161 36909 48195
rect 1777 48093 1811 48127
rect 21741 48093 21775 48127
rect 22293 48093 22327 48127
rect 24777 48093 24811 48127
rect 30757 48093 30791 48127
rect 49341 48093 49375 48127
rect 22569 48025 22603 48059
rect 25053 48025 25087 48059
rect 27353 48025 27387 48059
rect 36645 48025 36679 48059
rect 36737 48025 36771 48059
rect 19717 47957 19751 47991
rect 20085 47957 20119 47991
rect 20177 47957 20211 47991
rect 24041 47957 24075 47991
rect 26525 47957 26559 47991
rect 28825 47957 28859 47991
rect 32505 47957 32539 47991
rect 33425 47957 33459 47991
rect 35265 47957 35299 47991
rect 35357 47957 35391 47991
rect 36093 47957 36127 47991
rect 36277 47957 36311 47991
rect 49157 47957 49191 47991
rect 12265 47753 12299 47787
rect 21465 47753 21499 47787
rect 22017 47753 22051 47787
rect 24961 47753 24995 47787
rect 35173 47753 35207 47787
rect 35541 47753 35575 47787
rect 38301 47753 38335 47787
rect 38669 47753 38703 47787
rect 19993 47685 20027 47719
rect 22477 47685 22511 47719
rect 25881 47685 25915 47719
rect 27537 47685 27571 47719
rect 27629 47685 27663 47719
rect 33241 47685 33275 47719
rect 1777 47617 1811 47651
rect 12449 47617 12483 47651
rect 22385 47617 22419 47651
rect 25789 47617 25823 47651
rect 29469 47617 29503 47651
rect 32965 47617 32999 47651
rect 38761 47617 38795 47651
rect 49341 47617 49375 47651
rect 2053 47549 2087 47583
rect 19717 47549 19751 47583
rect 22661 47549 22695 47583
rect 23213 47549 23247 47583
rect 23489 47549 23523 47583
rect 26065 47549 26099 47583
rect 27721 47549 27755 47583
rect 29745 47549 29779 47583
rect 31217 47549 31251 47583
rect 35633 47549 35667 47583
rect 35725 47549 35759 47583
rect 38945 47549 38979 47583
rect 27169 47481 27203 47515
rect 25421 47413 25455 47447
rect 34713 47413 34747 47447
rect 49157 47413 49191 47447
rect 18153 47209 18187 47243
rect 24961 47209 24995 47243
rect 27905 47209 27939 47243
rect 28365 47209 28399 47243
rect 30941 47209 30975 47243
rect 34897 47209 34931 47243
rect 38485 47209 38519 47243
rect 20545 47141 20579 47175
rect 23949 47141 23983 47175
rect 29745 47141 29779 47175
rect 36093 47141 36127 47175
rect 18797 47073 18831 47107
rect 21189 47073 21223 47107
rect 22477 47073 22511 47107
rect 25605 47073 25639 47107
rect 26157 47073 26191 47107
rect 28917 47073 28951 47107
rect 30297 47073 30331 47107
rect 31401 47073 31435 47107
rect 31493 47073 31527 47107
rect 32597 47073 32631 47107
rect 32689 47073 32723 47107
rect 33793 47073 33827 47107
rect 33977 47073 34011 47107
rect 35541 47073 35575 47107
rect 36553 47073 36587 47107
rect 36645 47073 36679 47107
rect 39037 47073 39071 47107
rect 18521 47005 18555 47039
rect 20085 47005 20119 47039
rect 21005 47005 21039 47039
rect 22201 47005 22235 47039
rect 25329 47005 25363 47039
rect 28733 47005 28767 47039
rect 32505 47005 32539 47039
rect 33701 47005 33735 47039
rect 35265 47005 35299 47039
rect 35357 47005 35391 47039
rect 38853 47005 38887 47039
rect 18613 46937 18647 46971
rect 20913 46937 20947 46971
rect 25421 46937 25455 46971
rect 26433 46937 26467 46971
rect 30113 46937 30147 46971
rect 30205 46937 30239 46971
rect 31309 46937 31343 46971
rect 36461 46937 36495 46971
rect 38945 46937 38979 46971
rect 28825 46869 28859 46903
rect 32137 46869 32171 46903
rect 33333 46869 33367 46903
rect 11989 46665 12023 46699
rect 23765 46665 23799 46699
rect 26617 46665 26651 46699
rect 27997 46665 28031 46699
rect 29193 46665 29227 46699
rect 29285 46665 29319 46699
rect 32689 46665 32723 46699
rect 22293 46597 22327 46631
rect 27905 46597 27939 46631
rect 30297 46597 30331 46631
rect 1777 46529 1811 46563
rect 12173 46529 12207 46563
rect 24869 46529 24903 46563
rect 30021 46529 30055 46563
rect 34529 46529 34563 46563
rect 49065 46529 49099 46563
rect 2053 46461 2087 46495
rect 19717 46461 19751 46495
rect 19993 46461 20027 46495
rect 22017 46461 22051 46495
rect 25145 46461 25179 46495
rect 28181 46461 28215 46495
rect 29469 46461 29503 46495
rect 31769 46461 31803 46495
rect 32781 46461 32815 46495
rect 32873 46461 32907 46495
rect 34805 46461 34839 46495
rect 36277 46461 36311 46495
rect 27537 46393 27571 46427
rect 49249 46393 49283 46427
rect 21465 46325 21499 46359
rect 28825 46325 28859 46359
rect 32321 46325 32355 46359
rect 11069 46121 11103 46155
rect 19441 46121 19475 46155
rect 21998 46121 22032 46155
rect 23489 46121 23523 46155
rect 25053 46121 25087 46155
rect 30021 46121 30055 46155
rect 26249 46053 26283 46087
rect 31033 46053 31067 46087
rect 2053 45985 2087 46019
rect 21005 45985 21039 46019
rect 21189 45985 21223 46019
rect 21741 45985 21775 46019
rect 25697 45985 25731 46019
rect 26709 45985 26743 46019
rect 26801 45985 26835 46019
rect 27445 45985 27479 46019
rect 30573 45985 30607 46019
rect 31493 45985 31527 46019
rect 31585 45985 31619 46019
rect 33425 45985 33459 46019
rect 35173 45985 35207 46019
rect 38025 45985 38059 46019
rect 1777 45917 1811 45951
rect 19625 45917 19659 45951
rect 25421 45917 25455 45951
rect 26617 45917 26651 45951
rect 30481 45917 30515 45951
rect 31401 45917 31435 45951
rect 32321 45917 32355 45951
rect 33149 45917 33183 45951
rect 34161 45917 34195 45951
rect 37841 45917 37875 45951
rect 49065 45917 49099 45951
rect 10977 45849 11011 45883
rect 20913 45849 20947 45883
rect 27721 45849 27755 45883
rect 30389 45849 30423 45883
rect 33241 45849 33275 45883
rect 35449 45849 35483 45883
rect 20545 45781 20579 45815
rect 25513 45781 25547 45815
rect 29193 45781 29227 45815
rect 32781 45781 32815 45815
rect 36921 45781 36955 45815
rect 37473 45781 37507 45815
rect 37933 45781 37967 45815
rect 49249 45781 49283 45815
rect 22753 45577 22787 45611
rect 25145 45577 25179 45611
rect 25881 45577 25915 45611
rect 32965 45577 32999 45611
rect 33793 45577 33827 45611
rect 34161 45577 34195 45611
rect 7665 45509 7699 45543
rect 22661 45509 22695 45543
rect 23949 45509 23983 45543
rect 26341 45509 26375 45543
rect 27537 45509 27571 45543
rect 30113 45509 30147 45543
rect 33057 45509 33091 45543
rect 39681 45509 39715 45543
rect 7481 45441 7515 45475
rect 12173 45441 12207 45475
rect 13369 45441 13403 45475
rect 18245 45441 18279 45475
rect 19717 45441 19751 45475
rect 23857 45441 23891 45475
rect 25053 45441 25087 45475
rect 26249 45441 26283 45475
rect 27629 45441 27663 45475
rect 28733 45441 28767 45475
rect 31401 45441 31435 45475
rect 35725 45441 35759 45475
rect 36553 45441 36587 45475
rect 37841 45441 37875 45475
rect 39589 45441 39623 45475
rect 19993 45373 20027 45407
rect 22845 45373 22879 45407
rect 24041 45373 24075 45407
rect 25329 45373 25363 45407
rect 26525 45373 26559 45407
rect 27721 45373 27755 45407
rect 28825 45373 28859 45407
rect 28917 45373 28951 45407
rect 30205 45373 30239 45407
rect 30297 45373 30331 45407
rect 31493 45373 31527 45407
rect 31677 45373 31711 45407
rect 33149 45373 33183 45407
rect 34253 45373 34287 45407
rect 34437 45373 34471 45407
rect 36645 45373 36679 45407
rect 36737 45373 36771 45407
rect 37933 45373 37967 45407
rect 38025 45373 38059 45407
rect 39773 45373 39807 45407
rect 11989 45305 12023 45339
rect 18061 45305 18095 45339
rect 21465 45305 21499 45339
rect 23489 45305 23523 45339
rect 28365 45305 28399 45339
rect 31033 45305 31067 45339
rect 39221 45305 39255 45339
rect 13185 45237 13219 45271
rect 18889 45237 18923 45271
rect 22293 45237 22327 45271
rect 24685 45237 24719 45271
rect 27169 45237 27203 45271
rect 29745 45237 29779 45271
rect 32597 45237 32631 45271
rect 36185 45237 36219 45271
rect 37473 45237 37507 45271
rect 7297 45033 7331 45067
rect 12725 45033 12759 45067
rect 18153 45033 18187 45067
rect 26801 45033 26835 45067
rect 29745 45033 29779 45067
rect 36645 45033 36679 45067
rect 26341 44965 26375 44999
rect 27997 44965 28031 44999
rect 36737 44965 36771 44999
rect 49249 44965 49283 44999
rect 2053 44897 2087 44931
rect 18797 44897 18831 44931
rect 23765 44897 23799 44931
rect 23949 44897 23983 44931
rect 27261 44897 27295 44931
rect 27353 44897 27387 44931
rect 30389 44897 30423 44931
rect 31677 44897 31711 44931
rect 33425 44897 33459 44931
rect 34161 44897 34195 44931
rect 34897 44897 34931 44931
rect 37289 44897 37323 44931
rect 38025 44897 38059 44931
rect 38209 44897 38243 44931
rect 38945 44897 38979 44931
rect 1777 44829 1811 44863
rect 12909 44829 12943 44863
rect 18521 44829 18555 44863
rect 19901 44829 19935 44863
rect 22385 44829 22419 44863
rect 24593 44829 24627 44863
rect 27169 44829 27203 44863
rect 28181 44829 28215 44863
rect 28825 44829 28859 44863
rect 31401 44829 31435 44863
rect 33241 44829 33275 44863
rect 37105 44829 37139 44863
rect 38853 44829 38887 44863
rect 49065 44829 49099 44863
rect 7205 44761 7239 44795
rect 20177 44761 20211 44795
rect 24869 44761 24903 44795
rect 30113 44761 30147 44795
rect 31493 44761 31527 44795
rect 33149 44761 33183 44795
rect 35173 44761 35207 44795
rect 37197 44761 37231 44795
rect 37933 44761 37967 44795
rect 18613 44693 18647 44727
rect 21649 44693 21683 44727
rect 23305 44693 23339 44727
rect 23673 44693 23707 44727
rect 30205 44693 30239 44727
rect 31033 44693 31067 44727
rect 32781 44693 32815 44727
rect 37565 44693 37599 44727
rect 38393 44693 38427 44727
rect 38761 44693 38795 44727
rect 3893 44489 3927 44523
rect 10241 44489 10275 44523
rect 15485 44489 15519 44523
rect 17785 44489 17819 44523
rect 21097 44489 21131 44523
rect 22017 44489 22051 44523
rect 25605 44489 25639 44523
rect 28365 44489 28399 44523
rect 28733 44489 28767 44523
rect 29745 44489 29779 44523
rect 31401 44489 31435 44523
rect 32597 44489 32631 44523
rect 34253 44489 34287 44523
rect 34989 44489 35023 44523
rect 36185 44489 36219 44523
rect 36277 44489 36311 44523
rect 37933 44489 37967 44523
rect 39681 44489 39715 44523
rect 49157 44489 49191 44523
rect 5549 44421 5583 44455
rect 6837 44421 6871 44455
rect 22385 44421 22419 44455
rect 27537 44421 27571 44455
rect 31309 44421 31343 44455
rect 34161 44421 34195 44455
rect 1777 44353 1811 44387
rect 3801 44353 3835 44387
rect 5365 44353 5399 44387
rect 10425 44353 10459 44387
rect 15669 44353 15703 44387
rect 16313 44353 16347 44387
rect 17969 44353 18003 44387
rect 21189 44353 21223 44387
rect 25789 44353 25823 44387
rect 27629 44353 27663 44387
rect 30113 44353 30147 44387
rect 32965 44353 32999 44387
rect 35357 44353 35391 44387
rect 37841 44353 37875 44387
rect 40049 44353 40083 44387
rect 49341 44353 49375 44387
rect 2053 44285 2087 44319
rect 18429 44285 18463 44319
rect 18705 44285 18739 44319
rect 21281 44285 21315 44319
rect 22477 44285 22511 44319
rect 22661 44285 22695 44319
rect 23305 44285 23339 44319
rect 23581 44285 23615 44319
rect 25053 44285 25087 44319
rect 27721 44285 27755 44319
rect 28825 44285 28859 44319
rect 28917 44285 28951 44319
rect 30205 44285 30239 44319
rect 30297 44285 30331 44319
rect 31493 44285 31527 44319
rect 33057 44285 33091 44319
rect 33241 44285 33275 44319
rect 34345 44285 34379 44319
rect 35449 44285 35483 44319
rect 35633 44285 35667 44319
rect 36461 44285 36495 44319
rect 38025 44285 38059 44319
rect 40141 44285 40175 44319
rect 40233 44285 40267 44319
rect 16129 44217 16163 44251
rect 33793 44217 33827 44251
rect 37473 44217 37507 44251
rect 6929 44149 6963 44183
rect 20177 44149 20211 44183
rect 20729 44149 20763 44183
rect 27169 44149 27203 44183
rect 30941 44149 30975 44183
rect 35817 44149 35851 44183
rect 7849 43945 7883 43979
rect 12909 43945 12943 43979
rect 16129 43945 16163 43979
rect 18889 43945 18923 43979
rect 26617 43945 26651 43979
rect 27997 43945 28031 43979
rect 4721 43877 4755 43911
rect 5733 43877 5767 43911
rect 12265 43877 12299 43911
rect 39037 43877 39071 43911
rect 17141 43809 17175 43843
rect 20177 43809 20211 43843
rect 22293 43809 22327 43843
rect 23397 43809 23431 43843
rect 24869 43809 24903 43843
rect 28641 43809 28675 43843
rect 30297 43809 30331 43843
rect 31309 43809 31343 43843
rect 34161 43809 34195 43843
rect 35081 43809 35115 43843
rect 35357 43809 35391 43843
rect 37289 43809 37323 43843
rect 5549 43741 5583 43775
rect 12081 43741 12115 43775
rect 15669 43741 15703 43775
rect 16313 43741 16347 43775
rect 22109 43741 22143 43775
rect 23305 43741 23339 43775
rect 30205 43741 30239 43775
rect 34069 43741 34103 43775
rect 4537 43673 4571 43707
rect 7757 43673 7791 43707
rect 12817 43673 12851 43707
rect 17417 43673 17451 43707
rect 22017 43673 22051 43707
rect 25145 43673 25179 43707
rect 28365 43673 28399 43707
rect 30113 43673 30147 43707
rect 31585 43673 31619 43707
rect 37565 43673 37599 43707
rect 19533 43605 19567 43639
rect 19901 43605 19935 43639
rect 19993 43605 20027 43639
rect 21649 43605 21683 43639
rect 22845 43605 22879 43639
rect 23213 43605 23247 43639
rect 28457 43605 28491 43639
rect 29745 43605 29779 43639
rect 33057 43605 33091 43639
rect 33609 43605 33643 43639
rect 33977 43605 34011 43639
rect 36829 43605 36863 43639
rect 5641 43401 5675 43435
rect 8677 43401 8711 43435
rect 15577 43401 15611 43435
rect 15945 43401 15979 43435
rect 18889 43401 18923 43435
rect 21465 43401 21499 43435
rect 26433 43401 26467 43435
rect 27169 43401 27203 43435
rect 31217 43401 31251 43435
rect 35909 43401 35943 43435
rect 36001 43401 36035 43435
rect 49249 43401 49283 43435
rect 19993 43333 20027 43367
rect 22753 43333 22787 43367
rect 24961 43333 24995 43367
rect 1777 43265 1811 43299
rect 5549 43265 5583 43299
rect 8585 43265 8619 43299
rect 16037 43265 16071 43299
rect 18981 43265 19015 43299
rect 19717 43265 19751 43299
rect 27353 43265 27387 43299
rect 29469 43265 29503 43299
rect 32321 43265 32355 43299
rect 35081 43265 35115 43299
rect 49157 43265 49191 43299
rect 2053 43197 2087 43231
rect 16221 43197 16255 43231
rect 19165 43197 19199 43231
rect 22477 43197 22511 43231
rect 24685 43197 24719 43231
rect 29745 43197 29779 43231
rect 32597 43197 32631 43231
rect 36185 43197 36219 43231
rect 18521 43061 18555 43095
rect 24225 43061 24259 43095
rect 34069 43061 34103 43095
rect 35541 43061 35575 43095
rect 25973 42857 26007 42891
rect 26709 42857 26743 42891
rect 27708 42857 27742 42891
rect 35436 42857 35470 42891
rect 18153 42789 18187 42823
rect 2053 42721 2087 42755
rect 18613 42721 18647 42755
rect 18797 42721 18831 42755
rect 20269 42721 20303 42755
rect 23305 42721 23339 42755
rect 25237 42721 25271 42755
rect 27445 42721 27479 42755
rect 30481 42721 30515 42755
rect 31125 42721 31159 42755
rect 32873 42721 32907 42755
rect 33793 42721 33827 42755
rect 33885 42721 33919 42755
rect 35173 42721 35207 42755
rect 1777 42653 1811 42687
rect 15301 42653 15335 42687
rect 17049 42653 17083 42687
rect 17693 42653 17727 42687
rect 18521 42653 18555 42687
rect 19625 42653 19659 42687
rect 24961 42653 24995 42687
rect 26893 42653 26927 42687
rect 49065 42653 49099 42687
rect 15117 42585 15151 42619
rect 20545 42585 20579 42619
rect 22477 42585 22511 42619
rect 29745 42585 29779 42619
rect 31401 42585 31435 42619
rect 16865 42517 16899 42551
rect 17509 42517 17543 42551
rect 19441 42517 19475 42551
rect 22017 42517 22051 42551
rect 24593 42517 24627 42551
rect 25053 42517 25087 42551
rect 29193 42517 29227 42551
rect 33333 42517 33367 42551
rect 33701 42517 33735 42551
rect 36921 42517 36955 42551
rect 49249 42517 49283 42551
rect 11897 42313 11931 42347
rect 26157 42313 26191 42347
rect 29101 42313 29135 42347
rect 29193 42313 29227 42347
rect 31677 42313 31711 42347
rect 35081 42313 35115 42347
rect 19809 42245 19843 42279
rect 27169 42245 27203 42279
rect 30205 42245 30239 42279
rect 33609 42245 33643 42279
rect 36461 42245 36495 42279
rect 37933 42245 37967 42279
rect 11805 42177 11839 42211
rect 16313 42177 16347 42211
rect 16865 42177 16899 42211
rect 20545 42177 20579 42211
rect 22017 42177 22051 42211
rect 37841 42177 37875 42211
rect 17141 42109 17175 42143
rect 22293 42109 22327 42143
rect 24409 42109 24443 42143
rect 27905 42109 27939 42143
rect 29285 42109 29319 42143
rect 29936 42109 29970 42143
rect 33333 42109 33367 42143
rect 36553 42109 36587 42143
rect 36645 42109 36679 42143
rect 38025 42109 38059 42143
rect 18613 42041 18647 42075
rect 28733 42041 28767 42075
rect 16129 41973 16163 42007
rect 21373 41973 21407 42007
rect 23765 41973 23799 42007
rect 24672 41973 24706 42007
rect 36093 41973 36127 42007
rect 37473 41973 37507 42007
rect 11989 41769 12023 41803
rect 15025 41769 15059 41803
rect 22096 41769 22130 41803
rect 27629 41769 27663 41803
rect 31493 41769 31527 41803
rect 33701 41769 33735 41803
rect 35160 41769 35194 41803
rect 36645 41769 36679 41803
rect 13093 41701 13127 41735
rect 20729 41701 20763 41735
rect 26617 41701 26651 41735
rect 2053 41633 2087 41667
rect 15669 41633 15703 41667
rect 19901 41633 19935 41667
rect 20085 41633 20119 41667
rect 21281 41633 21315 41667
rect 21465 41633 21499 41667
rect 21833 41633 21867 41667
rect 23581 41633 23615 41667
rect 24869 41633 24903 41667
rect 28181 41633 28215 41667
rect 29745 41633 29779 41667
rect 30021 41633 30055 41667
rect 31953 41633 31987 41667
rect 32229 41633 32263 41667
rect 34897 41633 34931 41667
rect 1777 41565 1811 41599
rect 12173 41565 12207 41599
rect 13277 41565 13311 41599
rect 15393 41565 15427 41599
rect 16405 41565 16439 41599
rect 17233 41565 17267 41599
rect 18889 41565 18923 41599
rect 19809 41565 19843 41599
rect 24777 41565 24811 41599
rect 28089 41565 28123 41599
rect 29009 41565 29043 41599
rect 49065 41565 49099 41599
rect 15485 41497 15519 41531
rect 21189 41497 21223 41531
rect 25145 41497 25179 41531
rect 17049 41429 17083 41463
rect 19441 41429 19475 41463
rect 20821 41429 20855 41463
rect 24593 41429 24627 41463
rect 27077 41429 27111 41463
rect 27997 41429 28031 41463
rect 49249 41429 49283 41463
rect 13277 41225 13311 41259
rect 22385 41225 22419 41259
rect 23581 41225 23615 41259
rect 24777 41225 24811 41259
rect 25237 41225 25271 41259
rect 27721 41225 27755 41259
rect 28089 41225 28123 41259
rect 29561 41225 29595 41259
rect 30665 41225 30699 41259
rect 30757 41225 30791 41259
rect 31585 41225 31619 41259
rect 32321 41225 32355 41259
rect 36553 41225 36587 41259
rect 12633 41157 12667 41191
rect 13185 41157 13219 41191
rect 18245 41157 18279 41191
rect 23949 41157 23983 41191
rect 29653 41157 29687 41191
rect 33977 41157 34011 41191
rect 1777 41089 1811 41123
rect 15485 41089 15519 41123
rect 18889 41089 18923 41123
rect 21281 41089 21315 41123
rect 22753 41089 22787 41123
rect 25145 41089 25179 41123
rect 32689 41089 32723 41123
rect 32781 41089 32815 41123
rect 35725 41089 35759 41123
rect 36461 41089 36495 41123
rect 37473 41089 37507 41123
rect 49341 41089 49375 41123
rect 2053 41021 2087 41055
rect 19165 41021 19199 41055
rect 22845 41021 22879 41055
rect 23029 41021 23063 41055
rect 24041 41021 24075 41055
rect 24225 41021 24259 41055
rect 25421 41021 25455 41055
rect 28181 41021 28215 41055
rect 28273 41021 28307 41055
rect 29745 41021 29779 41055
rect 30849 41021 30883 41055
rect 32965 41021 32999 41055
rect 33701 41021 33735 41055
rect 36645 41021 36679 41055
rect 37749 41021 37783 41055
rect 29193 40953 29227 40987
rect 15301 40885 15335 40919
rect 18337 40885 18371 40919
rect 20637 40885 20671 40919
rect 30297 40885 30331 40919
rect 33517 40885 33551 40919
rect 36093 40885 36127 40919
rect 39221 40885 39255 40919
rect 49157 40885 49191 40919
rect 12265 40681 12299 40715
rect 17877 40681 17911 40715
rect 19441 40681 19475 40715
rect 26801 40681 26835 40715
rect 28089 40681 28123 40715
rect 38209 40681 38243 40715
rect 13093 40613 13127 40647
rect 30941 40613 30975 40647
rect 19901 40545 19935 40579
rect 19993 40545 20027 40579
rect 20637 40545 20671 40579
rect 22661 40545 22695 40579
rect 23857 40545 23891 40579
rect 27353 40545 27387 40579
rect 28733 40545 28767 40579
rect 30297 40545 30331 40579
rect 31401 40545 31435 40579
rect 31493 40545 31527 40579
rect 33149 40545 33183 40579
rect 37197 40545 37231 40579
rect 37657 40545 37691 40579
rect 38761 40545 38795 40579
rect 13277 40477 13311 40511
rect 15669 40477 15703 40511
rect 16129 40477 16163 40511
rect 18429 40477 18463 40511
rect 23765 40477 23799 40511
rect 25421 40477 25455 40511
rect 28457 40477 28491 40511
rect 30113 40477 30147 40511
rect 31309 40477 31343 40511
rect 32413 40477 32447 40511
rect 35173 40477 35207 40511
rect 38577 40477 38611 40511
rect 12173 40409 12207 40443
rect 16405 40409 16439 40443
rect 18613 40409 18647 40443
rect 19809 40409 19843 40443
rect 20913 40409 20947 40443
rect 26249 40409 26283 40443
rect 27261 40409 27295 40443
rect 35449 40409 35483 40443
rect 23305 40341 23339 40375
rect 23673 40341 23707 40375
rect 27169 40341 27203 40375
rect 28549 40341 28583 40375
rect 29745 40341 29779 40375
rect 30205 40341 30239 40375
rect 38669 40341 38703 40375
rect 14289 40137 14323 40171
rect 18153 40137 18187 40171
rect 18521 40137 18555 40171
rect 21373 40137 21407 40171
rect 22293 40137 22327 40171
rect 26341 40137 26375 40171
rect 27537 40137 27571 40171
rect 30297 40137 30331 40171
rect 36277 40137 36311 40171
rect 38669 40137 38703 40171
rect 19901 40069 19935 40103
rect 22661 40069 22695 40103
rect 23857 40069 23891 40103
rect 31401 40069 31435 40103
rect 39037 40069 39071 40103
rect 1777 40001 1811 40035
rect 14657 40001 14691 40035
rect 14749 40001 14783 40035
rect 15577 40001 15611 40035
rect 16129 40001 16163 40035
rect 23949 40001 23983 40035
rect 24593 40001 24627 40035
rect 31493 40001 31527 40035
rect 32321 40001 32355 40035
rect 34529 40001 34563 40035
rect 39129 40001 39163 40035
rect 49065 40001 49099 40035
rect 2053 39933 2087 39967
rect 14933 39933 14967 39967
rect 18613 39933 18647 39967
rect 18797 39933 18831 39967
rect 19625 39933 19659 39967
rect 22753 39933 22787 39967
rect 22845 39933 22879 39967
rect 24041 39933 24075 39967
rect 24869 39933 24903 39967
rect 27629 39933 27663 39967
rect 27721 39933 27755 39967
rect 28549 39933 28583 39967
rect 28825 39933 28859 39967
rect 31585 39933 31619 39967
rect 32597 39933 32631 39967
rect 34805 39933 34839 39967
rect 39313 39933 39347 39967
rect 17601 39865 17635 39899
rect 31033 39865 31067 39899
rect 38117 39865 38151 39899
rect 16221 39797 16255 39831
rect 23489 39797 23523 39831
rect 27169 39797 27203 39831
rect 34069 39797 34103 39831
rect 49249 39797 49283 39831
rect 13369 39593 13403 39627
rect 14933 39593 14967 39627
rect 17417 39593 17451 39627
rect 18153 39593 18187 39627
rect 24593 39593 24627 39627
rect 25881 39593 25915 39627
rect 26893 39593 26927 39627
rect 29101 39593 29135 39627
rect 31572 39593 31606 39627
rect 33057 39593 33091 39627
rect 23029 39525 23063 39559
rect 29745 39525 29779 39559
rect 38853 39525 38887 39559
rect 10701 39457 10735 39491
rect 15669 39457 15703 39491
rect 18705 39457 18739 39491
rect 20361 39457 20395 39491
rect 21465 39457 21499 39491
rect 23581 39457 23615 39491
rect 25145 39457 25179 39491
rect 26525 39457 26559 39491
rect 27353 39457 27387 39491
rect 30297 39457 30331 39491
rect 31309 39457 31343 39491
rect 34161 39457 34195 39491
rect 38577 39457 38611 39491
rect 39405 39457 39439 39491
rect 1777 39389 1811 39423
rect 12725 39389 12759 39423
rect 20085 39389 20119 39423
rect 22845 39389 22879 39423
rect 24961 39389 24995 39423
rect 25789 39389 25823 39423
rect 26249 39389 26283 39423
rect 34989 39389 35023 39423
rect 38393 39389 38427 39423
rect 2513 39321 2547 39355
rect 10977 39321 11011 39355
rect 13277 39321 13311 39355
rect 15945 39321 15979 39355
rect 18521 39321 18555 39355
rect 21281 39321 21315 39355
rect 21373 39321 21407 39355
rect 23489 39321 23523 39355
rect 27629 39321 27663 39355
rect 30113 39321 30147 39355
rect 34069 39321 34103 39355
rect 35265 39321 35299 39355
rect 37013 39321 37047 39355
rect 37473 39321 37507 39355
rect 39313 39321 39347 39355
rect 49157 39321 49191 39355
rect 18613 39253 18647 39287
rect 19717 39253 19751 39287
rect 20177 39253 20211 39287
rect 20913 39253 20947 39287
rect 22569 39253 22603 39287
rect 23397 39253 23431 39287
rect 25053 39253 25087 39287
rect 26341 39253 26375 39287
rect 30205 39253 30239 39287
rect 33609 39253 33643 39287
rect 33977 39253 34011 39287
rect 38025 39253 38059 39287
rect 38485 39253 38519 39287
rect 39221 39253 39255 39287
rect 49249 39253 49283 39287
rect 15485 39049 15519 39083
rect 15853 39049 15887 39083
rect 16957 39049 16991 39083
rect 17325 39049 17359 39083
rect 17969 39049 18003 39083
rect 18429 39049 18463 39083
rect 21465 39049 21499 39083
rect 23765 39049 23799 39083
rect 24225 39049 24259 39083
rect 24685 39049 24719 39083
rect 27537 39049 27571 39083
rect 30205 39049 30239 39083
rect 31033 39049 31067 39083
rect 34437 39049 34471 39083
rect 36921 39049 36955 39083
rect 39129 39049 39163 39083
rect 17417 38981 17451 39015
rect 15025 38913 15059 38947
rect 18337 38913 18371 38947
rect 19717 38913 19751 38947
rect 22017 38913 22051 38947
rect 24593 38913 24627 38947
rect 31401 38913 31435 38947
rect 33149 38913 33183 38947
rect 34345 38913 34379 38947
rect 35173 38913 35207 38947
rect 38117 38913 38151 38947
rect 39037 38913 39071 38947
rect 15945 38845 15979 38879
rect 16129 38845 16163 38879
rect 17601 38845 17635 38879
rect 18521 38845 18555 38879
rect 19993 38845 20027 38879
rect 22293 38845 22327 38879
rect 24777 38845 24811 38879
rect 27629 38845 27663 38879
rect 27721 38845 27755 38879
rect 28457 38845 28491 38879
rect 28733 38845 28767 38879
rect 31493 38845 31527 38879
rect 31677 38845 31711 38879
rect 33241 38845 33275 38879
rect 33425 38845 33459 38879
rect 34529 38845 34563 38879
rect 35449 38845 35483 38879
rect 39221 38845 39255 38879
rect 25605 38777 25639 38811
rect 14841 38709 14875 38743
rect 27169 38709 27203 38743
rect 32781 38709 32815 38743
rect 33977 38709 34011 38743
rect 38669 38709 38703 38743
rect 8401 38505 8435 38539
rect 12449 38505 12483 38539
rect 16865 38505 16899 38539
rect 19533 38505 19567 38539
rect 22109 38505 22143 38539
rect 25145 38505 25179 38539
rect 26341 38505 26375 38539
rect 37473 38505 37507 38539
rect 16221 38437 16255 38471
rect 23305 38437 23339 38471
rect 36277 38437 36311 38471
rect 38301 38437 38335 38471
rect 2053 38369 2087 38403
rect 13001 38369 13035 38403
rect 14473 38369 14507 38403
rect 20177 38369 20211 38403
rect 22753 38369 22787 38403
rect 23949 38369 23983 38403
rect 25789 38369 25823 38403
rect 27537 38369 27571 38403
rect 27629 38369 27663 38403
rect 33517 38369 33551 38403
rect 33701 38369 33735 38403
rect 36829 38369 36863 38403
rect 38025 38369 38059 38403
rect 38761 38369 38795 38403
rect 38945 38369 38979 38403
rect 1777 38301 1811 38335
rect 12909 38301 12943 38335
rect 16773 38301 16807 38335
rect 18705 38301 18739 38335
rect 19901 38301 19935 38335
rect 19993 38301 20027 38335
rect 23765 38301 23799 38335
rect 29101 38301 29135 38335
rect 29745 38301 29779 38335
rect 32229 38301 32263 38335
rect 37933 38301 37967 38335
rect 8309 38233 8343 38267
rect 14749 38233 14783 38267
rect 17325 38233 17359 38267
rect 17969 38233 18003 38267
rect 20729 38233 20763 38267
rect 21465 38233 21499 38267
rect 22477 38233 22511 38267
rect 28273 38233 28307 38267
rect 30021 38233 30055 38267
rect 34897 38233 34931 38267
rect 35633 38233 35667 38267
rect 37841 38233 37875 38267
rect 49157 38233 49191 38267
rect 12817 38165 12851 38199
rect 17417 38165 17451 38199
rect 22569 38165 22603 38199
rect 23673 38165 23707 38199
rect 25513 38165 25547 38199
rect 25605 38165 25639 38199
rect 27077 38165 27111 38199
rect 27445 38165 27479 38199
rect 31493 38165 31527 38199
rect 33057 38165 33091 38199
rect 33425 38165 33459 38199
rect 36645 38165 36679 38199
rect 36737 38165 36771 38199
rect 38669 38165 38703 38199
rect 49249 38165 49283 38199
rect 17969 37961 18003 37995
rect 20729 37961 20763 37995
rect 21097 37961 21131 37995
rect 25697 37961 25731 37995
rect 28917 37961 28951 37995
rect 31493 37961 31527 37995
rect 38669 37961 38703 37995
rect 39129 37961 39163 37995
rect 8493 37893 8527 37927
rect 19349 37893 19383 37927
rect 20269 37893 20303 37927
rect 21189 37893 21223 37927
rect 24961 37893 24995 37927
rect 37841 37893 37875 37927
rect 1777 37825 1811 37859
rect 13001 37825 13035 37859
rect 14565 37825 14599 37859
rect 17509 37825 17543 37859
rect 18337 37825 18371 37859
rect 22017 37825 22051 37859
rect 24869 37825 24903 37859
rect 26065 37825 26099 37859
rect 27169 37825 27203 37859
rect 29745 37825 29779 37859
rect 32505 37825 32539 37859
rect 35633 37825 35667 37859
rect 37933 37825 37967 37859
rect 39037 37825 39071 37859
rect 49341 37825 49375 37859
rect 2053 37757 2087 37791
rect 14841 37757 14875 37791
rect 18429 37757 18463 37791
rect 18613 37757 18647 37791
rect 19441 37757 19475 37791
rect 19533 37757 19567 37791
rect 21281 37757 21315 37791
rect 22293 37757 22327 37791
rect 24041 37757 24075 37791
rect 25053 37757 25087 37791
rect 26157 37757 26191 37791
rect 26249 37757 26283 37791
rect 27445 37757 27479 37791
rect 30021 37757 30055 37791
rect 32781 37757 32815 37791
rect 35725 37757 35759 37791
rect 35817 37757 35851 37791
rect 38025 37757 38059 37791
rect 39221 37757 39255 37791
rect 24501 37689 24535 37723
rect 35265 37689 35299 37723
rect 49157 37689 49191 37723
rect 8585 37621 8619 37655
rect 16313 37621 16347 37655
rect 18981 37621 19015 37655
rect 34253 37621 34287 37655
rect 34713 37621 34747 37655
rect 37473 37621 37507 37655
rect 21741 37417 21775 37451
rect 34253 37417 34287 37451
rect 13645 37281 13679 37315
rect 14933 37281 14967 37315
rect 15117 37281 15151 37315
rect 16129 37281 16163 37315
rect 18613 37281 18647 37315
rect 20361 37281 20395 37315
rect 23581 37281 23615 37315
rect 26801 37281 26835 37315
rect 30941 37281 30975 37315
rect 33425 37281 33459 37315
rect 35633 37281 35667 37315
rect 38117 37281 38151 37315
rect 13369 37213 13403 37247
rect 15853 37213 15887 37247
rect 20085 37213 20119 37247
rect 21097 37213 21131 37247
rect 23397 37213 23431 37247
rect 27445 37213 27479 37247
rect 30665 37213 30699 37247
rect 35357 37213 35391 37247
rect 37933 37213 37967 37247
rect 13461 37145 13495 37179
rect 18429 37145 18463 37179
rect 28181 37145 28215 37179
rect 33241 37145 33275 37179
rect 13001 37077 13035 37111
rect 14473 37077 14507 37111
rect 14841 37077 14875 37111
rect 17601 37077 17635 37111
rect 18061 37077 18095 37111
rect 18521 37077 18555 37111
rect 19717 37077 19751 37111
rect 20177 37077 20211 37111
rect 22937 37077 22971 37111
rect 23305 37077 23339 37111
rect 26249 37077 26283 37111
rect 26617 37077 26651 37111
rect 26709 37077 26743 37111
rect 32413 37077 32447 37111
rect 32873 37077 32907 37111
rect 33333 37077 33367 37111
rect 37105 37077 37139 37111
rect 37565 37077 37599 37111
rect 38025 37077 38059 37111
rect 12817 36873 12851 36907
rect 18613 36873 18647 36907
rect 19533 36873 19567 36907
rect 21097 36873 21131 36907
rect 22477 36873 22511 36907
rect 34161 36873 34195 36907
rect 36737 36873 36771 36907
rect 38761 36873 38795 36907
rect 13829 36805 13863 36839
rect 29193 36805 29227 36839
rect 35265 36805 35299 36839
rect 1777 36737 1811 36771
rect 12725 36737 12759 36771
rect 13553 36737 13587 36771
rect 16313 36737 16347 36771
rect 19441 36737 19475 36771
rect 22385 36737 22419 36771
rect 23581 36737 23615 36771
rect 26157 36737 26191 36771
rect 26249 36737 26283 36771
rect 27169 36737 27203 36771
rect 29653 36737 29687 36771
rect 38669 36737 38703 36771
rect 49065 36737 49099 36771
rect 2053 36669 2087 36703
rect 13001 36669 13035 36703
rect 16865 36669 16899 36703
rect 17141 36669 17175 36703
rect 19717 36669 19751 36703
rect 21189 36669 21223 36703
rect 21373 36669 21407 36703
rect 22661 36669 22695 36703
rect 23857 36669 23891 36703
rect 25329 36669 25363 36703
rect 26341 36669 26375 36703
rect 27445 36669 27479 36703
rect 29929 36669 29963 36703
rect 31401 36669 31435 36703
rect 32413 36669 32447 36703
rect 32689 36669 32723 36703
rect 34989 36669 35023 36703
rect 38853 36669 38887 36703
rect 16129 36601 16163 36635
rect 19073 36601 19107 36635
rect 20729 36601 20763 36635
rect 49249 36601 49283 36635
rect 12357 36533 12391 36567
rect 15301 36533 15335 36567
rect 22017 36533 22051 36567
rect 25789 36533 25823 36567
rect 38301 36533 38335 36567
rect 8493 36329 8527 36363
rect 9137 36329 9171 36363
rect 15577 36329 15611 36363
rect 21189 36329 21223 36363
rect 24041 36329 24075 36363
rect 26341 36329 26375 36363
rect 36737 36329 36771 36363
rect 49249 36329 49283 36363
rect 12173 36261 12207 36295
rect 18153 36261 18187 36295
rect 29193 36261 29227 36295
rect 31769 36261 31803 36295
rect 9689 36193 9723 36227
rect 13461 36193 13495 36227
rect 13645 36193 13679 36227
rect 15117 36193 15151 36227
rect 16129 36193 16163 36227
rect 16865 36193 16899 36227
rect 16957 36193 16991 36227
rect 18797 36193 18831 36227
rect 19441 36193 19475 36227
rect 22293 36193 22327 36227
rect 24593 36193 24627 36227
rect 27445 36193 27479 36227
rect 27721 36193 27755 36227
rect 30021 36193 30055 36227
rect 32781 36193 32815 36227
rect 37197 36193 37231 36227
rect 37473 36193 37507 36227
rect 1777 36125 1811 36159
rect 9505 36125 9539 36159
rect 11989 36125 12023 36159
rect 13369 36125 13403 36159
rect 17601 36125 17635 36159
rect 18613 36125 18647 36159
rect 33425 36125 33459 36159
rect 34989 36125 35023 36159
rect 49065 36125 49099 36159
rect 2789 36057 2823 36091
rect 8401 36057 8435 36091
rect 14933 36057 14967 36091
rect 15945 36057 15979 36091
rect 16037 36057 16071 36091
rect 18521 36057 18555 36091
rect 19717 36057 19751 36091
rect 22569 36057 22603 36091
rect 24869 36057 24903 36091
rect 30297 36057 30331 36091
rect 32597 36057 32631 36091
rect 32689 36057 32723 36091
rect 34161 36057 34195 36091
rect 35265 36057 35299 36091
rect 9597 35989 9631 36023
rect 13001 35989 13035 36023
rect 14565 35989 14599 36023
rect 15025 35989 15059 36023
rect 16405 35989 16439 36023
rect 16773 35989 16807 36023
rect 32229 35989 32263 36023
rect 38945 35989 38979 36023
rect 9413 35785 9447 35819
rect 14841 35785 14875 35819
rect 15945 35785 15979 35819
rect 17877 35785 17911 35819
rect 35909 35785 35943 35819
rect 9321 35717 9355 35751
rect 15853 35717 15887 35751
rect 19809 35717 19843 35751
rect 23213 35717 23247 35751
rect 32321 35717 32355 35751
rect 18245 35649 18279 35683
rect 22201 35649 22235 35683
rect 28273 35649 28307 35683
rect 30849 35649 30883 35683
rect 38209 35649 38243 35683
rect 9597 35581 9631 35615
rect 13093 35581 13127 35615
rect 13369 35581 13403 35615
rect 16129 35581 16163 35615
rect 18337 35581 18371 35615
rect 18429 35581 18463 35615
rect 19533 35581 19567 35615
rect 23305 35581 23339 35615
rect 23397 35581 23431 35615
rect 24133 35581 24167 35615
rect 24409 35581 24443 35615
rect 25881 35581 25915 35615
rect 28549 35581 28583 35615
rect 30941 35581 30975 35615
rect 31033 35581 31067 35615
rect 33057 35581 33091 35615
rect 34161 35581 34195 35615
rect 34437 35581 34471 35615
rect 17417 35513 17451 35547
rect 22845 35513 22879 35547
rect 30021 35513 30055 35547
rect 8953 35445 8987 35479
rect 15485 35445 15519 35479
rect 21281 35445 21315 35479
rect 30481 35445 30515 35479
rect 38025 35445 38059 35479
rect 16681 35241 16715 35275
rect 22385 35241 22419 35275
rect 23305 35241 23339 35275
rect 26433 35241 26467 35275
rect 30941 35241 30975 35275
rect 33425 35241 33459 35275
rect 16037 35173 16071 35207
rect 27537 35173 27571 35207
rect 29745 35173 29779 35207
rect 32137 35173 32171 35207
rect 2053 35105 2087 35139
rect 11805 35105 11839 35139
rect 13553 35105 13587 35139
rect 14289 35105 14323 35139
rect 17141 35105 17175 35139
rect 17325 35105 17359 35139
rect 18337 35105 18371 35139
rect 18521 35105 18555 35139
rect 19993 35105 20027 35139
rect 20637 35105 20671 35139
rect 20913 35105 20947 35139
rect 23765 35105 23799 35139
rect 23949 35105 23983 35139
rect 24685 35105 24719 35139
rect 27997 35105 28031 35139
rect 28181 35105 28215 35139
rect 30297 35105 30331 35139
rect 31585 35105 31619 35139
rect 32597 35105 32631 35139
rect 32689 35105 32723 35139
rect 33977 35105 34011 35139
rect 36645 35105 36679 35139
rect 1777 35037 1811 35071
rect 10885 35037 10919 35071
rect 13369 35037 13403 35071
rect 18245 35037 18279 35071
rect 19809 35037 19843 35071
rect 27905 35037 27939 35071
rect 29009 35037 29043 35071
rect 30113 35037 30147 35071
rect 33793 35037 33827 35071
rect 34897 35037 34931 35071
rect 40233 35037 40267 35071
rect 49065 35037 49099 35071
rect 11621 34969 11655 35003
rect 14565 34969 14599 35003
rect 17049 34969 17083 35003
rect 23673 34969 23707 35003
rect 24961 34969 24995 35003
rect 31309 34969 31343 35003
rect 35173 34969 35207 35003
rect 10977 34901 11011 34935
rect 13001 34901 13035 34935
rect 13461 34901 13495 34935
rect 17877 34901 17911 34935
rect 19441 34901 19475 34935
rect 19901 34901 19935 34935
rect 30205 34901 30239 34935
rect 31401 34901 31435 34935
rect 32505 34901 32539 34935
rect 33885 34901 33919 34935
rect 40049 34901 40083 34935
rect 49249 34901 49283 34935
rect 14289 34697 14323 34731
rect 14657 34697 14691 34731
rect 14749 34697 14783 34731
rect 15945 34697 15979 34731
rect 23765 34697 23799 34731
rect 26157 34697 26191 34731
rect 28917 34697 28951 34731
rect 32781 34697 32815 34731
rect 38301 34697 38335 34731
rect 41153 34697 41187 34731
rect 49157 34697 49191 34731
rect 13553 34629 13587 34663
rect 16957 34629 16991 34663
rect 22293 34629 22327 34663
rect 24685 34629 24719 34663
rect 1777 34561 1811 34595
rect 13461 34561 13495 34595
rect 16037 34561 16071 34595
rect 17141 34561 17175 34595
rect 18245 34561 18279 34595
rect 18337 34561 18371 34595
rect 19073 34561 19107 34595
rect 27169 34561 27203 34595
rect 29929 34561 29963 34595
rect 32689 34561 32723 34595
rect 38209 34561 38243 34595
rect 41337 34561 41371 34595
rect 49341 34561 49375 34595
rect 2053 34493 2087 34527
rect 13645 34493 13679 34527
rect 14933 34493 14967 34527
rect 16221 34493 16255 34527
rect 18429 34493 18463 34527
rect 20821 34493 20855 34527
rect 22017 34493 22051 34527
rect 24409 34493 24443 34527
rect 31677 34493 31711 34527
rect 32965 34493 32999 34527
rect 34529 34493 34563 34527
rect 38393 34493 38427 34527
rect 15577 34425 15611 34459
rect 17877 34425 17911 34459
rect 37841 34425 37875 34459
rect 13093 34357 13127 34391
rect 19336 34357 19370 34391
rect 27432 34357 27466 34391
rect 30186 34357 30220 34391
rect 32321 34357 32355 34391
rect 33701 34357 33735 34391
rect 34792 34357 34826 34391
rect 36277 34357 36311 34391
rect 14289 34153 14323 34187
rect 17233 34153 17267 34187
rect 20256 34153 20290 34187
rect 21741 34153 21775 34187
rect 24593 34153 24627 34187
rect 25973 34153 26007 34187
rect 28089 34153 28123 34187
rect 35725 34153 35759 34187
rect 29745 34085 29779 34119
rect 35081 34085 35115 34119
rect 11897 34017 11931 34051
rect 12081 34017 12115 34051
rect 14933 34017 14967 34051
rect 15485 34017 15519 34051
rect 18613 34017 18647 34051
rect 18705 34017 18739 34051
rect 19993 34017 20027 34051
rect 25145 34017 25179 34051
rect 28733 34017 28767 34051
rect 30205 34017 30239 34051
rect 30297 34017 30331 34051
rect 31585 34017 31619 34051
rect 32873 34017 32907 34051
rect 11805 33949 11839 33983
rect 13737 33949 13771 33983
rect 14657 33949 14691 33983
rect 18521 33949 18555 33983
rect 22937 33949 22971 33983
rect 23765 33949 23799 33983
rect 24961 33949 24995 33983
rect 25053 33949 25087 33983
rect 27629 33949 27663 33983
rect 28549 33949 28583 33983
rect 30113 33949 30147 33983
rect 31309 33949 31343 33983
rect 32597 33949 32631 33983
rect 15761 33881 15795 33915
rect 22201 33881 22235 33915
rect 28457 33881 28491 33915
rect 11437 33813 11471 33847
rect 14749 33813 14783 33847
rect 18153 33813 18187 33847
rect 30941 33813 30975 33847
rect 31401 33813 31435 33847
rect 34345 33813 34379 33847
rect 14381 33609 14415 33643
rect 14749 33609 14783 33643
rect 17785 33609 17819 33643
rect 20729 33609 20763 33643
rect 21097 33609 21131 33643
rect 26065 33609 26099 33643
rect 16037 33541 16071 33575
rect 18613 33541 18647 33575
rect 19349 33541 19383 33575
rect 21189 33541 21223 33575
rect 27445 33541 27479 33575
rect 1777 33473 1811 33507
rect 15945 33473 15979 33507
rect 17877 33473 17911 33507
rect 24317 33473 24351 33507
rect 27169 33473 27203 33507
rect 29561 33473 29595 33507
rect 30021 33473 30055 33507
rect 32505 33473 32539 33507
rect 39681 33473 39715 33507
rect 41061 33473 41095 33507
rect 49157 33473 49191 33507
rect 2053 33405 2087 33439
rect 14841 33405 14875 33439
rect 14933 33405 14967 33439
rect 16221 33405 16255 33439
rect 17969 33405 18003 33439
rect 21281 33405 21315 33439
rect 22017 33405 22051 33439
rect 22293 33405 22327 33439
rect 24593 33405 24627 33439
rect 30297 33405 30331 33439
rect 33057 33405 33091 33439
rect 33333 33405 33367 33439
rect 49341 33405 49375 33439
rect 15577 33337 15611 33371
rect 34805 33337 34839 33371
rect 39497 33337 39531 33371
rect 17417 33269 17451 33303
rect 23765 33269 23799 33303
rect 28917 33269 28951 33303
rect 31769 33269 31803 33303
rect 40877 33269 40911 33303
rect 19625 33065 19659 33099
rect 23121 33065 23155 33099
rect 24593 33065 24627 33099
rect 27629 33065 27663 33099
rect 49249 33065 49283 33099
rect 20177 32997 20211 33031
rect 32137 32997 32171 33031
rect 2053 32929 2087 32963
rect 15945 32929 15979 32963
rect 20729 32929 20763 32963
rect 21649 32929 21683 32963
rect 25237 32929 25271 32963
rect 28273 32929 28307 32963
rect 30021 32929 30055 32963
rect 32597 32929 32631 32963
rect 1777 32861 1811 32895
rect 14841 32861 14875 32895
rect 20545 32861 20579 32895
rect 21373 32861 21407 32895
rect 24041 32861 24075 32895
rect 24961 32861 24995 32895
rect 27997 32861 28031 32895
rect 29193 32861 29227 32895
rect 29745 32861 29779 32895
rect 49065 32861 49099 32895
rect 16221 32793 16255 32827
rect 28089 32793 28123 32827
rect 32873 32793 32907 32827
rect 17693 32725 17727 32759
rect 20637 32725 20671 32759
rect 25053 32725 25087 32759
rect 31493 32725 31527 32759
rect 34345 32725 34379 32759
rect 12909 32521 12943 32555
rect 21005 32521 21039 32555
rect 22017 32521 22051 32555
rect 22477 32521 22511 32555
rect 30941 32521 30975 32555
rect 32321 32521 32355 32555
rect 36645 32521 36679 32555
rect 12449 32453 12483 32487
rect 13277 32453 13311 32487
rect 14565 32453 14599 32487
rect 19533 32453 19567 32487
rect 23949 32453 23983 32487
rect 28549 32453 28583 32487
rect 12633 32385 12667 32419
rect 14289 32385 14323 32419
rect 17417 32385 17451 32419
rect 19257 32385 19291 32419
rect 22385 32385 22419 32419
rect 30849 32385 30883 32419
rect 32689 32385 32723 32419
rect 33885 32385 33919 32419
rect 36553 32385 36587 32419
rect 13369 32317 13403 32351
rect 13553 32317 13587 32351
rect 17509 32317 17543 32351
rect 17693 32317 17727 32351
rect 22569 32317 22603 32351
rect 23673 32317 23707 32351
rect 28273 32317 28307 32351
rect 30021 32317 30055 32351
rect 31033 32317 31067 32351
rect 32781 32317 32815 32351
rect 32965 32317 32999 32351
rect 33977 32317 34011 32351
rect 34069 32317 34103 32351
rect 36737 32317 36771 32351
rect 30481 32249 30515 32283
rect 33517 32249 33551 32283
rect 12725 32181 12759 32215
rect 14197 32181 14231 32215
rect 16037 32181 16071 32215
rect 17049 32181 17083 32215
rect 25421 32181 25455 32215
rect 36185 32181 36219 32215
rect 16589 31977 16623 32011
rect 18797 31977 18831 32011
rect 21097 31977 21131 32011
rect 24041 31977 24075 32011
rect 28273 31977 28307 32011
rect 31953 31977 31987 32011
rect 33149 31977 33183 32011
rect 25881 31909 25915 31943
rect 31493 31909 31527 31943
rect 49249 31909 49283 31943
rect 2053 31841 2087 31875
rect 14841 31841 14875 31875
rect 17325 31841 17359 31875
rect 20269 31841 20303 31875
rect 20453 31841 20487 31875
rect 21649 31841 21683 31875
rect 22293 31841 22327 31875
rect 22569 31841 22603 31875
rect 26341 31841 26375 31875
rect 26525 31841 26559 31875
rect 28733 31841 28767 31875
rect 28917 31841 28951 31875
rect 29745 31841 29779 31875
rect 32413 31841 32447 31875
rect 32505 31841 32539 31875
rect 33701 31841 33735 31875
rect 1777 31773 1811 31807
rect 8033 31773 8067 31807
rect 10977 31773 11011 31807
rect 17049 31773 17083 31807
rect 27813 31773 27847 31807
rect 33609 31773 33643 31807
rect 49065 31773 49099 31807
rect 7849 31705 7883 31739
rect 15117 31705 15151 31739
rect 20177 31705 20211 31739
rect 21557 31705 21591 31739
rect 30021 31705 30055 31739
rect 33517 31705 33551 31739
rect 11069 31637 11103 31671
rect 19809 31637 19843 31671
rect 21465 31637 21499 31671
rect 26249 31637 26283 31671
rect 28641 31637 28675 31671
rect 32321 31637 32355 31671
rect 13185 31433 13219 31467
rect 13553 31433 13587 31467
rect 13645 31433 13679 31467
rect 14749 31433 14783 31467
rect 15945 31433 15979 31467
rect 16037 31433 16071 31467
rect 17417 31433 17451 31467
rect 27629 31433 27663 31467
rect 29561 31433 29595 31467
rect 17509 31365 17543 31399
rect 44465 31365 44499 31399
rect 1777 31297 1811 31331
rect 10701 31297 10735 31331
rect 18245 31297 18279 31331
rect 20821 31297 20855 31331
rect 28641 31297 28675 31331
rect 29653 31297 29687 31331
rect 32505 31297 32539 31331
rect 38393 31297 38427 31331
rect 49341 31297 49375 31331
rect 2053 31229 2087 31263
rect 13737 31229 13771 31263
rect 14841 31229 14875 31263
rect 15025 31229 15059 31263
rect 16221 31229 16255 31263
rect 17601 31229 17635 31263
rect 18521 31229 18555 31263
rect 20913 31229 20947 31263
rect 21097 31229 21131 31263
rect 27721 31229 27755 31263
rect 27905 31229 27939 31263
rect 29837 31229 29871 31263
rect 14381 31161 14415 31195
rect 19993 31161 20027 31195
rect 27261 31161 27295 31195
rect 44649 31161 44683 31195
rect 49157 31161 49191 31195
rect 10793 31093 10827 31127
rect 15577 31093 15611 31127
rect 17049 31093 17083 31127
rect 20453 31093 20487 31127
rect 23397 31093 23431 31127
rect 24409 31093 24443 31127
rect 29193 31093 29227 31127
rect 38209 31093 38243 31127
rect 24593 30889 24627 30923
rect 26157 30889 26191 30923
rect 14933 30753 14967 30787
rect 15025 30753 15059 30787
rect 17877 30753 17911 30787
rect 20913 30753 20947 30787
rect 21005 30753 21039 30787
rect 23765 30753 23799 30787
rect 23949 30753 23983 30787
rect 25237 30753 25271 30787
rect 26801 30753 26835 30787
rect 13737 30685 13771 30719
rect 14841 30685 14875 30719
rect 15853 30685 15887 30719
rect 24961 30685 24995 30719
rect 26525 30685 26559 30719
rect 45293 30685 45327 30719
rect 12817 30617 12851 30651
rect 13553 30617 13587 30651
rect 16129 30617 16163 30651
rect 20821 30617 20855 30651
rect 25053 30617 25087 30651
rect 45477 30617 45511 30651
rect 12909 30549 12943 30583
rect 14473 30549 14507 30583
rect 20453 30549 20487 30583
rect 23305 30549 23339 30583
rect 23673 30549 23707 30583
rect 26617 30549 26651 30583
rect 23213 30345 23247 30379
rect 23305 30277 23339 30311
rect 1777 30209 1811 30243
rect 17417 30209 17451 30243
rect 19717 30209 19751 30243
rect 22201 30209 22235 30243
rect 37657 30209 37691 30243
rect 49065 30209 49099 30243
rect 2053 30141 2087 30175
rect 14105 30141 14139 30175
rect 14381 30141 14415 30175
rect 18153 30141 18187 30175
rect 19993 30141 20027 30175
rect 21465 30141 21499 30175
rect 23397 30141 23431 30175
rect 15853 30005 15887 30039
rect 22845 30005 22879 30039
rect 29285 30005 29319 30039
rect 37473 30005 37507 30039
rect 49249 30005 49283 30039
rect 27169 29801 27203 29835
rect 2053 29665 2087 29699
rect 18889 29665 18923 29699
rect 20177 29665 20211 29699
rect 21925 29665 21959 29699
rect 29009 29665 29043 29699
rect 49341 29665 49375 29699
rect 1777 29597 1811 29631
rect 14657 29597 14691 29631
rect 16865 29597 16899 29631
rect 19901 29597 19935 29631
rect 22569 29597 22603 29631
rect 28825 29597 28859 29631
rect 29929 29597 29963 29631
rect 46581 29597 46615 29631
rect 14933 29529 14967 29563
rect 17141 29529 17175 29563
rect 25881 29529 25915 29563
rect 45845 29529 45879 29563
rect 46765 29529 46799 29563
rect 49157 29529 49191 29563
rect 16405 29461 16439 29495
rect 28457 29461 28491 29495
rect 28917 29461 28951 29495
rect 45937 29461 45971 29495
rect 15577 29257 15611 29291
rect 16037 29257 16071 29291
rect 21465 29257 21499 29291
rect 22017 29257 22051 29291
rect 22385 29257 22419 29291
rect 24961 29257 24995 29291
rect 28733 29257 28767 29291
rect 29101 29257 29135 29291
rect 24501 29189 24535 29223
rect 25421 29189 25455 29223
rect 15945 29121 15979 29155
rect 17325 29121 17359 29155
rect 19717 29121 19751 29155
rect 22477 29121 22511 29155
rect 25329 29121 25363 29155
rect 16221 29053 16255 29087
rect 17601 29053 17635 29087
rect 19073 29053 19107 29087
rect 22661 29053 22695 29087
rect 25605 29053 25639 29087
rect 29193 29053 29227 29087
rect 29285 29053 29319 29087
rect 19980 28917 20014 28951
rect 18889 28713 18923 28747
rect 2053 28577 2087 28611
rect 15945 28577 15979 28611
rect 17141 28577 17175 28611
rect 17417 28577 17451 28611
rect 21557 28577 21591 28611
rect 1777 28509 1811 28543
rect 15761 28509 15795 28543
rect 19533 28509 19567 28543
rect 21281 28509 21315 28543
rect 37289 28509 37323 28543
rect 49065 28509 49099 28543
rect 20269 28441 20303 28475
rect 15393 28373 15427 28407
rect 15853 28373 15887 28407
rect 20913 28373 20947 28407
rect 21373 28373 21407 28407
rect 37105 28373 37139 28407
rect 49249 28373 49283 28407
rect 15301 28169 15335 28203
rect 16957 28169 16991 28203
rect 17417 28169 17451 28203
rect 18521 28169 18555 28203
rect 18889 28169 18923 28203
rect 19717 28169 19751 28203
rect 14289 28101 14323 28135
rect 15761 28101 15795 28135
rect 45201 28101 45235 28135
rect 1777 28033 1811 28067
rect 15669 28033 15703 28067
rect 17325 28033 17359 28067
rect 20085 28033 20119 28067
rect 49341 28033 49375 28067
rect 2053 27965 2087 27999
rect 15945 27965 15979 27999
rect 17509 27965 17543 27999
rect 18981 27965 19015 27999
rect 19073 27965 19107 27999
rect 20177 27965 20211 27999
rect 20361 27965 20395 27999
rect 49157 27897 49191 27931
rect 14749 27829 14783 27863
rect 45293 27829 45327 27863
rect 15393 27557 15427 27591
rect 15853 27489 15887 27523
rect 16037 27489 16071 27523
rect 17049 27489 17083 27523
rect 17233 27489 17267 27523
rect 18705 27489 18739 27523
rect 15761 27421 15795 27455
rect 16957 27421 16991 27455
rect 18521 27421 18555 27455
rect 18613 27353 18647 27387
rect 38945 27353 38979 27387
rect 39129 27353 39163 27387
rect 16589 27285 16623 27319
rect 18153 27285 18187 27319
rect 21097 27081 21131 27115
rect 21189 27013 21223 27047
rect 44557 27013 44591 27047
rect 1685 26945 1719 26979
rect 47961 26945 47995 26979
rect 21373 26877 21407 26911
rect 49157 26877 49191 26911
rect 44741 26809 44775 26843
rect 1777 26741 1811 26775
rect 20729 26741 20763 26775
rect 18153 26469 18187 26503
rect 18613 26401 18647 26435
rect 18797 26401 18831 26435
rect 48421 26401 48455 26435
rect 1869 26333 1903 26367
rect 18521 26333 18555 26367
rect 47961 26333 47995 26367
rect 1685 26265 1719 26299
rect 38853 25925 38887 25959
rect 38209 25857 38243 25891
rect 39037 25721 39071 25755
rect 38025 25653 38059 25687
rect 1869 25313 1903 25347
rect 1593 25245 1627 25279
rect 47961 25245 47995 25279
rect 49157 25245 49191 25279
rect 1685 24769 1719 24803
rect 39589 24769 39623 24803
rect 39957 24769 39991 24803
rect 47961 24769 47995 24803
rect 39313 24701 39347 24735
rect 49157 24701 49191 24735
rect 39773 24633 39807 24667
rect 1961 24565 1995 24599
rect 40049 24565 40083 24599
rect 15853 24157 15887 24191
rect 37657 24157 37691 24191
rect 44097 24157 44131 24191
rect 44281 24089 44315 24123
rect 15669 24021 15703 24055
rect 37473 24021 37507 24055
rect 1869 23749 1903 23783
rect 39129 23749 39163 23783
rect 1685 23681 1719 23715
rect 36921 23681 36955 23715
rect 47961 23681 47995 23715
rect 49157 23613 49191 23647
rect 39313 23545 39347 23579
rect 36737 23477 36771 23511
rect 1869 23137 1903 23171
rect 1593 23069 1627 23103
rect 47961 23069 47995 23103
rect 49157 23001 49191 23035
rect 43913 21981 43947 22015
rect 47961 21981 47995 22015
rect 49157 21981 49191 22015
rect 1685 21913 1719 21947
rect 44097 21913 44131 21947
rect 1961 21845 1995 21879
rect 1685 21505 1719 21539
rect 37565 21505 37599 21539
rect 47961 21505 47995 21539
rect 49157 21437 49191 21471
rect 37749 21369 37783 21403
rect 1961 21301 1995 21335
rect 40141 20825 40175 20859
rect 40325 20825 40359 20859
rect 1685 20417 1719 20451
rect 47961 20417 47995 20451
rect 49157 20349 49191 20383
rect 1961 20213 1995 20247
rect 47961 19805 47995 19839
rect 1685 19737 1719 19771
rect 49157 19737 49191 19771
rect 1777 19669 1811 19703
rect 17785 19465 17819 19499
rect 22109 19465 22143 19499
rect 44465 19397 44499 19431
rect 17969 19329 18003 19363
rect 22293 19329 22327 19363
rect 38669 19329 38703 19363
rect 38853 19193 38887 19227
rect 44649 19193 44683 19227
rect 1593 18717 1627 18751
rect 20177 18717 20211 18751
rect 40141 18717 40175 18751
rect 47961 18717 47995 18751
rect 49157 18717 49191 18751
rect 40325 18649 40359 18683
rect 1777 18581 1811 18615
rect 19993 18581 20027 18615
rect 1593 18241 1627 18275
rect 47961 18241 47995 18275
rect 49157 18173 49191 18207
rect 1777 18037 1811 18071
rect 38025 17629 38059 17663
rect 38209 17561 38243 17595
rect 1685 17153 1719 17187
rect 2053 17153 2087 17187
rect 38117 17153 38151 17187
rect 47961 17153 47995 17187
rect 49157 17085 49191 17119
rect 38301 17017 38335 17051
rect 1869 16609 1903 16643
rect 38117 16609 38151 16643
rect 44373 16609 44407 16643
rect 44189 16541 44223 16575
rect 47961 16541 47995 16575
rect 1685 16473 1719 16507
rect 37933 16473 37967 16507
rect 49157 16473 49191 16507
rect 24961 16133 24995 16167
rect 38209 16065 38243 16099
rect 38853 16065 38887 16099
rect 24777 15997 24811 16031
rect 25237 15997 25271 16031
rect 38393 15929 38427 15963
rect 26709 15521 26743 15555
rect 26249 15453 26283 15487
rect 47961 15453 47995 15487
rect 49157 15453 49191 15487
rect 1685 15385 1719 15419
rect 26433 15385 26467 15419
rect 1961 15317 1995 15351
rect 28181 15045 28215 15079
rect 43729 15045 43763 15079
rect 1685 14977 1719 15011
rect 47961 14977 47995 15011
rect 27997 14909 28031 14943
rect 29377 14909 29411 14943
rect 49157 14909 49191 14943
rect 1961 14773 1995 14807
rect 43821 14773 43855 14807
rect 30389 14433 30423 14467
rect 29837 14365 29871 14399
rect 30021 14297 30055 14331
rect 1593 13889 1627 13923
rect 37565 13889 37599 13923
rect 47961 13889 47995 13923
rect 37749 13821 37783 13855
rect 49157 13821 49191 13855
rect 1777 13753 1811 13787
rect 1869 13345 1903 13379
rect 18245 13345 18279 13379
rect 1593 13277 1627 13311
rect 18429 13277 18463 13311
rect 37657 13277 37691 13311
rect 47961 13277 47995 13311
rect 37841 13209 37875 13243
rect 49157 13209 49191 13243
rect 18889 13141 18923 13175
rect 23535 12937 23569 12971
rect 23464 12801 23498 12835
rect 38301 12801 38335 12835
rect 38393 12597 38427 12631
rect 24731 12393 24765 12427
rect 25467 12393 25501 12427
rect 26755 12393 26789 12427
rect 24628 12189 24662 12223
rect 25364 12189 25398 12223
rect 26652 12189 26686 12223
rect 47961 12189 47995 12223
rect 49157 12189 49191 12223
rect 1685 12121 1719 12155
rect 1961 12053 1995 12087
rect 1685 11713 1719 11747
rect 19993 11713 20027 11747
rect 47961 11713 47995 11747
rect 20177 11645 20211 11679
rect 49157 11645 49191 11679
rect 1961 11577 1995 11611
rect 20637 11509 20671 11543
rect 36737 11237 36771 11271
rect 21925 11169 21959 11203
rect 22109 11169 22143 11203
rect 24593 11169 24627 11203
rect 24777 11169 24811 11203
rect 37381 11101 37415 11135
rect 22569 11033 22603 11067
rect 25237 11033 25271 11067
rect 37565 11033 37599 11067
rect 1685 10625 1719 10659
rect 37565 10625 37599 10659
rect 38209 10625 38243 10659
rect 47961 10625 47995 10659
rect 49157 10557 49191 10591
rect 37749 10489 37783 10523
rect 1961 10421 1995 10455
rect 26065 10081 26099 10115
rect 47961 10013 47995 10047
rect 1685 9945 1719 9979
rect 26341 9945 26375 9979
rect 49157 9945 49191 9979
rect 1777 9877 1811 9911
rect 27813 9877 27847 9911
rect 22017 9537 22051 9571
rect 36277 9537 36311 9571
rect 22293 9469 22327 9503
rect 36461 9401 36495 9435
rect 23765 9333 23799 9367
rect 1593 8925 1627 8959
rect 47961 8925 47995 8959
rect 49157 8925 49191 8959
rect 1777 8789 1811 8823
rect 25605 8585 25639 8619
rect 1593 8449 1627 8483
rect 25145 8449 25179 8483
rect 27169 8449 27203 8483
rect 32689 8449 32723 8483
rect 47961 8449 47995 8483
rect 32965 8381 32999 8415
rect 49157 8381 49191 8415
rect 1777 8313 1811 8347
rect 25421 8245 25455 8279
rect 27445 8245 27479 8279
rect 27629 8245 27663 8279
rect 34437 8245 34471 8279
rect 23029 8041 23063 8075
rect 23397 8041 23431 8075
rect 22937 7837 22971 7871
rect 1685 7361 1719 7395
rect 30757 7361 30791 7395
rect 47961 7361 47995 7395
rect 49157 7293 49191 7327
rect 31217 7225 31251 7259
rect 1961 7157 1995 7191
rect 30297 7157 30331 7191
rect 31033 7157 31067 7191
rect 19533 6749 19567 6783
rect 47961 6749 47995 6783
rect 1685 6681 1719 6715
rect 49157 6681 49191 6715
rect 1777 6613 1811 6647
rect 19625 6613 19659 6647
rect 13001 5797 13035 5831
rect 11253 5729 11287 5763
rect 21373 5661 21407 5695
rect 24685 5661 24719 5695
rect 26617 5661 26651 5695
rect 47961 5661 47995 5695
rect 49157 5661 49191 5695
rect 1685 5593 1719 5627
rect 11529 5593 11563 5627
rect 21557 5593 21591 5627
rect 24869 5593 24903 5627
rect 26801 5593 26835 5627
rect 1961 5525 1995 5559
rect 13553 5253 13587 5287
rect 1685 5185 1719 5219
rect 47961 5185 47995 5219
rect 49157 5117 49191 5151
rect 1961 4981 1995 5015
rect 13645 4981 13679 5015
rect 17601 4641 17635 4675
rect 15301 4573 15335 4607
rect 19533 4573 19567 4607
rect 17417 4505 17451 4539
rect 15393 4437 15427 4471
rect 19625 4437 19659 4471
rect 1593 4097 1627 4131
rect 47961 4097 47995 4131
rect 49157 4029 49191 4063
rect 1777 3893 1811 3927
rect 47961 3485 47995 3519
rect 1685 3417 1719 3451
rect 49157 3417 49191 3451
rect 1777 3349 1811 3383
rect 28825 3009 28859 3043
rect 29285 2941 29319 2975
rect 7021 2465 7055 2499
rect 9689 2465 9723 2499
rect 12725 2465 12759 2499
rect 15485 2465 15519 2499
rect 19901 2465 19935 2499
rect 22661 2465 22695 2499
rect 25697 2465 25731 2499
rect 38945 2465 38979 2499
rect 42901 2465 42935 2499
rect 2513 2397 2547 2431
rect 6745 2397 6779 2431
rect 9321 2397 9355 2431
rect 12357 2397 12391 2431
rect 15117 2397 15151 2431
rect 19625 2397 19659 2431
rect 22201 2397 22235 2431
rect 25237 2397 25271 2431
rect 32505 2397 32539 2431
rect 35449 2397 35483 2431
rect 35725 2397 35759 2431
rect 38669 2397 38703 2431
rect 42625 2397 42659 2431
rect 47961 2397 47995 2431
rect 45477 2329 45511 2363
rect 49157 2329 49191 2363
rect 2329 2261 2363 2295
rect 32321 2261 32355 2295
rect 45569 2261 45603 2295
<< metal1 >>
rect 30558 54612 30564 54664
rect 30616 54652 30622 54664
rect 37458 54652 37464 54664
rect 30616 54624 37464 54652
rect 30616 54612 30622 54624
rect 37458 54612 37464 54624
rect 37516 54612 37522 54664
rect 32490 54544 32496 54596
rect 32548 54584 32554 54596
rect 45830 54584 45836 54596
rect 32548 54556 45836 54584
rect 32548 54544 32554 54556
rect 45830 54544 45836 54556
rect 45888 54544 45894 54596
rect 34514 54476 34520 54528
rect 34572 54516 34578 54528
rect 40678 54516 40684 54528
rect 34572 54488 40684 54516
rect 34572 54476 34578 54488
rect 40678 54476 40684 54488
rect 40736 54476 40742 54528
rect 1104 54426 49864 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 27950 54426
rect 28002 54374 28014 54426
rect 28066 54374 28078 54426
rect 28130 54374 28142 54426
rect 28194 54374 28206 54426
rect 28258 54374 37950 54426
rect 38002 54374 38014 54426
rect 38066 54374 38078 54426
rect 38130 54374 38142 54426
rect 38194 54374 38206 54426
rect 38258 54374 47950 54426
rect 48002 54374 48014 54426
rect 48066 54374 48078 54426
rect 48130 54374 48142 54426
rect 48194 54374 48206 54426
rect 48258 54374 49864 54426
rect 1104 54352 49864 54374
rect 23201 54315 23259 54321
rect 23201 54281 23213 54315
rect 23247 54281 23259 54315
rect 23201 54275 23259 54281
rect 24857 54315 24915 54321
rect 24857 54281 24869 54315
rect 24903 54312 24915 54315
rect 30098 54312 30104 54324
rect 24903 54284 30104 54312
rect 24903 54281 24915 54284
rect 24857 54275 24915 54281
rect 3237 54247 3295 54253
rect 3237 54213 3249 54247
rect 3283 54244 3295 54247
rect 3510 54244 3516 54256
rect 3283 54216 3516 54244
rect 3283 54213 3295 54216
rect 3237 54207 3295 54213
rect 3510 54204 3516 54216
rect 3568 54204 3574 54256
rect 5534 54244 5540 54256
rect 3804 54216 5540 54244
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 3804 54176 3832 54216
rect 5534 54204 5540 54216
rect 5592 54204 5598 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 8662 54244 8668 54256
rect 8435 54216 8668 54244
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 8662 54204 8668 54216
rect 8720 54204 8726 54256
rect 10594 54204 10600 54256
rect 10652 54244 10658 54256
rect 10689 54247 10747 54253
rect 10689 54244 10701 54247
rect 10652 54216 10701 54244
rect 10652 54204 10658 54216
rect 10689 54213 10701 54216
rect 10735 54213 10747 54247
rect 10689 54207 10747 54213
rect 13541 54247 13599 54253
rect 13541 54213 13553 54247
rect 13587 54244 13599 54247
rect 13814 54244 13820 54256
rect 13587 54216 13820 54244
rect 13587 54213 13599 54216
rect 13541 54207 13599 54213
rect 13814 54204 13820 54216
rect 13872 54204 13878 54256
rect 15746 54204 15752 54256
rect 15804 54244 15810 54256
rect 15841 54247 15899 54253
rect 15841 54244 15853 54247
rect 15804 54216 15853 54244
rect 15804 54204 15810 54216
rect 15841 54213 15853 54216
rect 15887 54213 15899 54247
rect 15841 54207 15899 54213
rect 18693 54247 18751 54253
rect 18693 54213 18705 54247
rect 18739 54244 18751 54247
rect 18966 54244 18972 54256
rect 18739 54216 18972 54244
rect 18739 54213 18751 54216
rect 18693 54207 18751 54213
rect 18966 54204 18972 54216
rect 19024 54204 19030 54256
rect 20714 54244 20720 54256
rect 20088 54216 20720 54244
rect 2271 54148 3832 54176
rect 4801 54179 4859 54185
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4801 54145 4813 54179
rect 4847 54176 4859 54179
rect 4890 54176 4896 54188
rect 4847 54148 4896 54176
rect 4847 54145 4859 54148
rect 4801 54139 4859 54145
rect 4890 54136 4896 54148
rect 4948 54136 4954 54188
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54145 7435 54179
rect 7377 54139 7435 54145
rect 9953 54179 10011 54185
rect 9953 54145 9965 54179
rect 9999 54176 10011 54179
rect 10502 54176 10508 54188
rect 9999 54148 10508 54176
rect 9999 54145 10011 54148
rect 9953 54139 10011 54145
rect 5442 54068 5448 54120
rect 5500 54068 5506 54120
rect 7392 54108 7420 54139
rect 10502 54136 10508 54148
rect 10560 54136 10566 54188
rect 12529 54179 12587 54185
rect 12529 54145 12541 54179
rect 12575 54176 12587 54179
rect 13722 54176 13728 54188
rect 12575 54148 13728 54176
rect 12575 54145 12587 54148
rect 12529 54139 12587 54145
rect 13722 54136 13728 54148
rect 13780 54136 13786 54188
rect 15010 54136 15016 54188
rect 15068 54136 15074 54188
rect 17681 54179 17739 54185
rect 17681 54145 17693 54179
rect 17727 54176 17739 54179
rect 20088 54176 20116 54216
rect 20714 54204 20720 54216
rect 20772 54204 20778 54256
rect 23216 54244 23244 54275
rect 30098 54272 30104 54284
rect 30156 54272 30162 54324
rect 32214 54272 32220 54324
rect 32272 54312 32278 54324
rect 32272 54284 45554 54312
rect 32272 54272 32278 54284
rect 28258 54244 28264 54256
rect 23216 54216 28264 54244
rect 28258 54204 28264 54216
rect 28316 54204 28322 54256
rect 30190 54204 30196 54256
rect 30248 54244 30254 54256
rect 33686 54244 33692 54256
rect 30248 54216 33692 54244
rect 30248 54204 30254 54216
rect 33686 54204 33692 54216
rect 33744 54204 33750 54256
rect 35250 54204 35256 54256
rect 35308 54244 35314 54256
rect 35308 54216 36952 54244
rect 35308 54204 35314 54216
rect 17727 54148 20116 54176
rect 20165 54179 20223 54185
rect 17727 54145 17739 54148
rect 17681 54139 17739 54145
rect 20165 54145 20177 54179
rect 20211 54176 20223 54179
rect 22741 54179 22799 54185
rect 20211 54148 22048 54176
rect 20211 54145 20223 54148
rect 20165 54139 20223 54145
rect 15378 54108 15384 54120
rect 7392 54080 15384 54108
rect 15378 54068 15384 54080
rect 15436 54068 15442 54120
rect 20254 54068 20260 54120
rect 20312 54108 20318 54120
rect 20533 54111 20591 54117
rect 20533 54108 20545 54111
rect 20312 54080 20545 54108
rect 20312 54068 20318 54080
rect 20533 54077 20545 54080
rect 20579 54077 20591 54111
rect 22020 54108 22048 54148
rect 22741 54145 22753 54179
rect 22787 54176 22799 54179
rect 22830 54176 22836 54188
rect 22787 54148 22836 54176
rect 22787 54145 22799 54148
rect 22741 54139 22799 54145
rect 22830 54136 22836 54148
rect 22888 54136 22894 54188
rect 23385 54179 23443 54185
rect 23385 54145 23397 54179
rect 23431 54176 23443 54179
rect 23474 54176 23480 54188
rect 23431 54148 23480 54176
rect 23431 54145 23443 54148
rect 23385 54139 23443 54145
rect 23474 54136 23480 54148
rect 23532 54136 23538 54188
rect 24029 54179 24087 54185
rect 24029 54145 24041 54179
rect 24075 54176 24087 54179
rect 24118 54176 24124 54188
rect 24075 54148 24124 54176
rect 24075 54145 24087 54148
rect 24029 54139 24087 54145
rect 24118 54136 24124 54148
rect 24176 54136 24182 54188
rect 24762 54136 24768 54188
rect 24820 54176 24826 54188
rect 25041 54179 25099 54185
rect 25041 54176 25053 54179
rect 24820 54148 25053 54176
rect 24820 54136 24826 54148
rect 25041 54145 25053 54148
rect 25087 54145 25099 54179
rect 25041 54139 25099 54145
rect 25406 54136 25412 54188
rect 25464 54176 25470 54188
rect 25685 54179 25743 54185
rect 25685 54176 25697 54179
rect 25464 54148 25697 54176
rect 25464 54136 25470 54148
rect 25685 54145 25697 54148
rect 25731 54145 25743 54179
rect 25685 54139 25743 54145
rect 26234 54136 26240 54188
rect 26292 54176 26298 54188
rect 26329 54179 26387 54185
rect 26329 54176 26341 54179
rect 26292 54148 26341 54176
rect 26292 54136 26298 54148
rect 26329 54145 26341 54148
rect 26375 54145 26387 54179
rect 26329 54139 26387 54145
rect 26694 54136 26700 54188
rect 26752 54176 26758 54188
rect 27341 54179 27399 54185
rect 27341 54176 27353 54179
rect 26752 54148 27353 54176
rect 26752 54136 26758 54148
rect 27341 54145 27353 54148
rect 27387 54145 27399 54179
rect 27341 54139 27399 54145
rect 27430 54136 27436 54188
rect 27488 54176 27494 54188
rect 27985 54179 28043 54185
rect 27985 54176 27997 54179
rect 27488 54148 27997 54176
rect 27488 54136 27494 54148
rect 27985 54145 27997 54148
rect 28031 54145 28043 54179
rect 27985 54139 28043 54145
rect 28350 54136 28356 54188
rect 28408 54176 28414 54188
rect 28629 54179 28687 54185
rect 28629 54176 28641 54179
rect 28408 54148 28641 54176
rect 28408 54136 28414 54148
rect 28629 54145 28641 54148
rect 28675 54145 28687 54179
rect 28629 54139 28687 54145
rect 29270 54136 29276 54188
rect 29328 54176 29334 54188
rect 29917 54179 29975 54185
rect 29917 54176 29929 54179
rect 29328 54148 29929 54176
rect 29328 54136 29334 54148
rect 29917 54145 29929 54148
rect 29963 54145 29975 54179
rect 29917 54139 29975 54145
rect 30282 54136 30288 54188
rect 30340 54176 30346 54188
rect 30561 54179 30619 54185
rect 30561 54176 30573 54179
rect 30340 54148 30573 54176
rect 30340 54136 30346 54148
rect 30561 54145 30573 54148
rect 30607 54145 30619 54179
rect 30561 54139 30619 54145
rect 30650 54136 30656 54188
rect 30708 54176 30714 54188
rect 31205 54179 31263 54185
rect 31205 54176 31217 54179
rect 30708 54148 31217 54176
rect 30708 54136 30714 54148
rect 31205 54145 31217 54148
rect 31251 54145 31263 54179
rect 31205 54139 31263 54145
rect 31846 54136 31852 54188
rect 31904 54176 31910 54188
rect 32493 54179 32551 54185
rect 32493 54176 32505 54179
rect 31904 54148 32505 54176
rect 31904 54136 31910 54148
rect 32493 54145 32505 54148
rect 32539 54145 32551 54179
rect 32493 54139 32551 54145
rect 32582 54136 32588 54188
rect 32640 54176 32646 54188
rect 33137 54179 33195 54185
rect 33137 54176 33149 54179
rect 32640 54148 33149 54176
rect 32640 54136 32646 54148
rect 33137 54145 33149 54148
rect 33183 54145 33195 54179
rect 33137 54139 33195 54145
rect 33226 54136 33232 54188
rect 33284 54176 33290 54188
rect 33781 54179 33839 54185
rect 33781 54176 33793 54179
rect 33284 54148 33793 54176
rect 33284 54136 33290 54148
rect 33781 54145 33793 54148
rect 33827 54145 33839 54179
rect 33781 54139 33839 54145
rect 35066 54136 35072 54188
rect 35124 54176 35130 54188
rect 35161 54179 35219 54185
rect 35161 54176 35173 54179
rect 35124 54148 35173 54176
rect 35124 54136 35130 54148
rect 35161 54145 35173 54148
rect 35207 54145 35219 54179
rect 35161 54139 35219 54145
rect 35894 54136 35900 54188
rect 35952 54176 35958 54188
rect 36633 54179 36691 54185
rect 36633 54176 36645 54179
rect 35952 54148 36645 54176
rect 35952 54136 35958 54148
rect 36633 54145 36645 54148
rect 36679 54145 36691 54179
rect 36633 54139 36691 54145
rect 23566 54108 23572 54120
rect 22020 54080 23572 54108
rect 20533 54071 20591 54077
rect 23566 54068 23572 54080
rect 23624 54068 23630 54120
rect 27706 54108 27712 54120
rect 23860 54080 27712 54108
rect 23860 54049 23888 54080
rect 27706 54068 27712 54080
rect 27764 54068 27770 54120
rect 28810 54108 28816 54120
rect 27816 54080 28816 54108
rect 23845 54043 23903 54049
rect 23845 54009 23857 54043
rect 23891 54009 23903 54043
rect 23845 54003 23903 54009
rect 26145 54043 26203 54049
rect 26145 54009 26157 54043
rect 26191 54040 26203 54043
rect 27816 54040 27844 54080
rect 28810 54068 28816 54080
rect 28868 54068 28874 54120
rect 29730 54068 29736 54120
rect 29788 54108 29794 54120
rect 35437 54111 35495 54117
rect 35437 54108 35449 54111
rect 29788 54080 35449 54108
rect 29788 54068 29794 54080
rect 35437 54077 35449 54080
rect 35483 54077 35495 54111
rect 36924 54108 36952 54216
rect 37182 54204 37188 54256
rect 37240 54244 37246 54256
rect 37240 54216 39068 54244
rect 37240 54204 37246 54216
rect 36998 54136 37004 54188
rect 37056 54176 37062 54188
rect 37645 54179 37703 54185
rect 37645 54176 37657 54179
rect 37056 54148 37657 54176
rect 37056 54136 37062 54148
rect 37645 54145 37657 54148
rect 37691 54145 37703 54179
rect 37645 54139 37703 54145
rect 37734 54136 37740 54188
rect 37792 54176 37798 54188
rect 38289 54179 38347 54185
rect 38289 54176 38301 54179
rect 37792 54148 38301 54176
rect 37792 54136 37798 54148
rect 38289 54145 38301 54148
rect 38335 54145 38347 54179
rect 38289 54139 38347 54145
rect 38378 54136 38384 54188
rect 38436 54176 38442 54188
rect 38933 54179 38991 54185
rect 38933 54176 38945 54179
rect 38436 54148 38945 54176
rect 38436 54136 38442 54148
rect 38933 54145 38945 54148
rect 38979 54145 38991 54179
rect 38933 54139 38991 54145
rect 39040 54108 39068 54216
rect 39114 54204 39120 54256
rect 39172 54244 39178 54256
rect 40770 54244 40776 54256
rect 39172 54216 40776 54244
rect 39172 54204 39178 54216
rect 40770 54204 40776 54216
rect 40828 54204 40834 54256
rect 42150 54204 42156 54256
rect 42208 54244 42214 54256
rect 42613 54247 42671 54253
rect 42613 54244 42625 54247
rect 42208 54216 42625 54244
rect 42208 54204 42214 54216
rect 42613 54213 42625 54216
rect 42659 54213 42671 54247
rect 42613 54207 42671 54213
rect 39574 54136 39580 54188
rect 39632 54176 39638 54188
rect 40221 54179 40279 54185
rect 40221 54176 40233 54179
rect 39632 54148 40233 54176
rect 39632 54136 39638 54148
rect 40221 54145 40233 54148
rect 40267 54145 40279 54179
rect 40221 54139 40279 54145
rect 40310 54136 40316 54188
rect 40368 54176 40374 54188
rect 40865 54179 40923 54185
rect 40865 54176 40877 54179
rect 40368 54148 40877 54176
rect 40368 54136 40374 54148
rect 40865 54145 40877 54148
rect 40911 54145 40923 54179
rect 40865 54139 40923 54145
rect 44726 54136 44732 54188
rect 44784 54176 44790 54188
rect 45189 54179 45247 54185
rect 45189 54176 45201 54179
rect 44784 54148 45201 54176
rect 44784 54136 44790 54148
rect 45189 54145 45201 54148
rect 45235 54145 45247 54179
rect 45526 54176 45554 54284
rect 45830 54272 45836 54324
rect 45888 54312 45894 54324
rect 46109 54315 46167 54321
rect 46109 54312 46121 54315
rect 45888 54284 46121 54312
rect 45888 54272 45894 54284
rect 46109 54281 46121 54284
rect 46155 54281 46167 54315
rect 46109 54275 46167 54281
rect 45646 54204 45652 54256
rect 45704 54244 45710 54256
rect 46017 54247 46075 54253
rect 46017 54244 46029 54247
rect 45704 54216 46029 54244
rect 45704 54204 45710 54216
rect 46017 54213 46029 54216
rect 46063 54213 46075 54247
rect 46017 54207 46075 54213
rect 45526 54148 46060 54176
rect 45189 54139 45247 54145
rect 46032 54108 46060 54148
rect 46106 54136 46112 54188
rect 46164 54176 46170 54188
rect 46845 54179 46903 54185
rect 46845 54176 46857 54179
rect 46164 54148 46857 54176
rect 46164 54136 46170 54148
rect 46845 54145 46857 54148
rect 46891 54145 46903 54179
rect 46845 54139 46903 54145
rect 47302 54136 47308 54188
rect 47360 54176 47366 54188
rect 47765 54179 47823 54185
rect 47765 54176 47777 54179
rect 47360 54148 47777 54176
rect 47360 54136 47366 54148
rect 47765 54145 47777 54148
rect 47811 54145 47823 54179
rect 47765 54139 47823 54145
rect 47854 54136 47860 54188
rect 47912 54176 47918 54188
rect 48501 54179 48559 54185
rect 48501 54176 48513 54179
rect 47912 54148 48513 54176
rect 47912 54136 47918 54148
rect 48501 54145 48513 54148
rect 48547 54145 48559 54179
rect 48501 54139 48559 54145
rect 36924 54080 38792 54108
rect 39040 54080 40080 54108
rect 35437 54071 35495 54077
rect 26191 54012 27844 54040
rect 26191 54009 26203 54012
rect 26145 54003 26203 54009
rect 27890 54000 27896 54052
rect 27948 54040 27954 54052
rect 28445 54043 28503 54049
rect 28445 54040 28457 54043
rect 27948 54012 28457 54040
rect 27948 54000 27954 54012
rect 28445 54009 28457 54012
rect 28491 54009 28503 54043
rect 28445 54003 28503 54009
rect 31938 54000 31944 54052
rect 31996 54040 32002 54052
rect 38764 54049 38792 54080
rect 40052 54049 40080 54080
rect 40144 54080 45554 54108
rect 46032 54080 47992 54108
rect 38105 54043 38163 54049
rect 38105 54040 38117 54043
rect 31996 54012 38117 54040
rect 31996 54000 32002 54012
rect 38105 54009 38117 54012
rect 38151 54009 38163 54043
rect 38105 54003 38163 54009
rect 38749 54043 38807 54049
rect 38749 54009 38761 54043
rect 38795 54009 38807 54043
rect 38749 54003 38807 54009
rect 40037 54043 40095 54049
rect 40037 54009 40049 54043
rect 40083 54009 40095 54043
rect 40037 54003 40095 54009
rect 22557 53975 22615 53981
rect 22557 53941 22569 53975
rect 22603 53972 22615 53975
rect 25406 53972 25412 53984
rect 22603 53944 25412 53972
rect 22603 53941 22615 53944
rect 22557 53935 22615 53941
rect 25406 53932 25412 53944
rect 25464 53932 25470 53984
rect 25501 53975 25559 53981
rect 25501 53941 25513 53975
rect 25547 53972 25559 53975
rect 26050 53972 26056 53984
rect 25547 53944 26056 53972
rect 25547 53941 25559 53944
rect 25501 53935 25559 53941
rect 26050 53932 26056 53944
rect 26108 53932 26114 53984
rect 27157 53975 27215 53981
rect 27157 53941 27169 53975
rect 27203 53972 27215 53975
rect 27430 53972 27436 53984
rect 27203 53944 27436 53972
rect 27203 53941 27215 53944
rect 27157 53935 27215 53941
rect 27430 53932 27436 53944
rect 27488 53932 27494 53984
rect 27801 53975 27859 53981
rect 27801 53941 27813 53975
rect 27847 53972 27859 53975
rect 28350 53972 28356 53984
rect 27847 53944 28356 53972
rect 27847 53941 27859 53944
rect 27801 53935 27859 53941
rect 28350 53932 28356 53944
rect 28408 53932 28414 53984
rect 29086 53932 29092 53984
rect 29144 53972 29150 53984
rect 29733 53975 29791 53981
rect 29733 53972 29745 53975
rect 29144 53944 29745 53972
rect 29144 53932 29150 53944
rect 29733 53941 29745 53944
rect 29779 53941 29791 53975
rect 29733 53935 29791 53941
rect 30374 53932 30380 53984
rect 30432 53932 30438 53984
rect 30742 53932 30748 53984
rect 30800 53972 30806 53984
rect 31021 53975 31079 53981
rect 31021 53972 31033 53975
rect 30800 53944 31033 53972
rect 30800 53932 30806 53944
rect 31021 53941 31033 53944
rect 31067 53941 31079 53975
rect 31021 53935 31079 53941
rect 32306 53932 32312 53984
rect 32364 53932 32370 53984
rect 32582 53932 32588 53984
rect 32640 53972 32646 53984
rect 32953 53975 33011 53981
rect 32953 53972 32965 53975
rect 32640 53944 32965 53972
rect 32640 53932 32646 53944
rect 32953 53941 32965 53944
rect 32999 53941 33011 53975
rect 32953 53935 33011 53941
rect 33594 53932 33600 53984
rect 33652 53932 33658 53984
rect 33686 53932 33692 53984
rect 33744 53972 33750 53984
rect 36449 53975 36507 53981
rect 36449 53972 36461 53975
rect 33744 53944 36461 53972
rect 33744 53932 33750 53944
rect 36449 53941 36461 53944
rect 36495 53941 36507 53975
rect 36449 53935 36507 53941
rect 37458 53932 37464 53984
rect 37516 53932 37522 53984
rect 37550 53932 37556 53984
rect 37608 53972 37614 53984
rect 40144 53972 40172 54080
rect 40678 54000 40684 54052
rect 40736 54000 40742 54052
rect 40770 54000 40776 54052
rect 40828 54040 40834 54052
rect 45373 54043 45431 54049
rect 45373 54040 45385 54043
rect 40828 54012 45385 54040
rect 40828 54000 40834 54012
rect 45373 54009 45385 54012
rect 45419 54009 45431 54043
rect 45526 54040 45554 54080
rect 47964 54049 47992 54080
rect 47029 54043 47087 54049
rect 47029 54040 47041 54043
rect 45526 54012 47041 54040
rect 45373 54003 45431 54009
rect 47029 54009 47041 54012
rect 47075 54009 47087 54043
rect 47029 54003 47087 54009
rect 47949 54043 48007 54049
rect 47949 54009 47961 54043
rect 47995 54009 48007 54043
rect 47949 54003 48007 54009
rect 37608 53944 40172 53972
rect 37608 53932 37614 53944
rect 43898 53932 43904 53984
rect 43956 53932 43962 53984
rect 48682 53932 48688 53984
rect 48740 53932 48746 53984
rect 1104 53882 49864 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 32950 53882
rect 33002 53830 33014 53882
rect 33066 53830 33078 53882
rect 33130 53830 33142 53882
rect 33194 53830 33206 53882
rect 33258 53830 42950 53882
rect 43002 53830 43014 53882
rect 43066 53830 43078 53882
rect 43130 53830 43142 53882
rect 43194 53830 43206 53882
rect 43258 53830 49864 53882
rect 1104 53808 49864 53830
rect 22094 53700 22100 53712
rect 15856 53672 22100 53700
rect 2866 53592 2872 53644
rect 2924 53592 2930 53644
rect 6086 53592 6092 53644
rect 6144 53592 6150 53644
rect 7834 53592 7840 53644
rect 7892 53592 7898 53644
rect 11238 53592 11244 53644
rect 11296 53592 11302 53644
rect 13354 53592 13360 53644
rect 13412 53592 13418 53644
rect 2038 53524 2044 53576
rect 2096 53524 2102 53576
rect 5445 53567 5503 53573
rect 5445 53533 5457 53567
rect 5491 53533 5503 53567
rect 5445 53527 5503 53533
rect 7377 53567 7435 53573
rect 7377 53533 7389 53567
rect 7423 53564 7435 53567
rect 8478 53564 8484 53576
rect 7423 53536 8484 53564
rect 7423 53533 7435 53536
rect 7377 53527 7435 53533
rect 5460 53496 5488 53527
rect 8478 53524 8484 53536
rect 8536 53524 8542 53576
rect 10689 53567 10747 53573
rect 10689 53533 10701 53567
rect 10735 53533 10747 53567
rect 10689 53527 10747 53533
rect 12529 53567 12587 53573
rect 12529 53533 12541 53567
rect 12575 53564 12587 53567
rect 15194 53564 15200 53576
rect 12575 53536 15200 53564
rect 12575 53533 12587 53536
rect 12529 53527 12587 53533
rect 8386 53496 8392 53508
rect 5460 53468 8392 53496
rect 8386 53456 8392 53468
rect 8444 53456 8450 53508
rect 10704 53496 10732 53527
rect 15194 53524 15200 53536
rect 15252 53524 15258 53576
rect 15856 53573 15884 53672
rect 22094 53660 22100 53672
rect 22152 53660 22158 53712
rect 23569 53703 23627 53709
rect 23569 53669 23581 53703
rect 23615 53669 23627 53703
rect 23569 53663 23627 53669
rect 16390 53592 16396 53644
rect 16448 53592 16454 53644
rect 18322 53592 18328 53644
rect 18380 53592 18386 53644
rect 23584 53632 23612 53663
rect 29454 53660 29460 53712
rect 29512 53700 29518 53712
rect 36449 53703 36507 53709
rect 36449 53700 36461 53703
rect 29512 53672 36461 53700
rect 29512 53660 29518 53672
rect 36449 53669 36461 53672
rect 36495 53669 36507 53703
rect 36449 53663 36507 53669
rect 38654 53660 38660 53712
rect 38712 53700 38718 53712
rect 48225 53703 48283 53709
rect 48225 53700 48237 53703
rect 38712 53672 48237 53700
rect 38712 53660 38718 53672
rect 48225 53669 48237 53672
rect 48271 53669 48283 53703
rect 48225 53663 48283 53669
rect 21192 53604 23612 53632
rect 21192 53573 21220 53604
rect 34422 53592 34428 53644
rect 34480 53632 34486 53644
rect 34885 53635 34943 53641
rect 34885 53632 34897 53635
rect 34480 53604 34897 53632
rect 34480 53592 34486 53604
rect 34885 53601 34897 53604
rect 34931 53601 34943 53635
rect 34885 53595 34943 53601
rect 38286 53592 38292 53644
rect 38344 53632 38350 53644
rect 44453 53635 44511 53641
rect 44453 53632 44465 53635
rect 38344 53604 44465 53632
rect 38344 53592 38350 53604
rect 44453 53601 44465 53604
rect 44499 53601 44511 53635
rect 44453 53595 44511 53601
rect 15841 53567 15899 53573
rect 15841 53533 15853 53567
rect 15887 53533 15899 53567
rect 15841 53527 15899 53533
rect 17681 53567 17739 53573
rect 17681 53533 17693 53567
rect 17727 53533 17739 53567
rect 17681 53527 17739 53533
rect 21177 53567 21235 53573
rect 21177 53533 21189 53567
rect 21223 53533 21235 53567
rect 21177 53527 21235 53533
rect 13538 53496 13544 53508
rect 10704 53468 13544 53496
rect 13538 53456 13544 53468
rect 13596 53456 13602 53508
rect 17696 53428 17724 53527
rect 22186 53524 22192 53576
rect 22244 53564 22250 53576
rect 23017 53567 23075 53573
rect 23017 53564 23029 53567
rect 22244 53536 23029 53564
rect 22244 53524 22250 53536
rect 23017 53533 23029 53536
rect 23063 53533 23075 53567
rect 23017 53527 23075 53533
rect 23753 53567 23811 53573
rect 23753 53533 23765 53567
rect 23799 53564 23811 53567
rect 26234 53564 26240 53576
rect 23799 53536 26240 53564
rect 23799 53533 23811 53536
rect 23753 53527 23811 53533
rect 26234 53524 26240 53536
rect 26292 53524 26298 53576
rect 28626 53524 28632 53576
rect 28684 53564 28690 53576
rect 28905 53567 28963 53573
rect 28905 53564 28917 53567
rect 28684 53536 28917 53564
rect 28684 53524 28690 53536
rect 28905 53533 28917 53536
rect 28951 53533 28963 53567
rect 28905 53527 28963 53533
rect 31202 53524 31208 53576
rect 31260 53564 31266 53576
rect 31481 53567 31539 53573
rect 31481 53564 31493 53567
rect 31260 53536 31493 53564
rect 31260 53524 31266 53536
rect 31481 53533 31493 53536
rect 31527 53533 31539 53567
rect 31481 53527 31539 53533
rect 33778 53524 33784 53576
rect 33836 53564 33842 53576
rect 34057 53567 34115 53573
rect 34057 53564 34069 53567
rect 33836 53536 34069 53564
rect 33836 53524 33842 53536
rect 34057 53533 34069 53536
rect 34103 53533 34115 53567
rect 34057 53527 34115 53533
rect 35161 53567 35219 53573
rect 35161 53533 35173 53567
rect 35207 53533 35219 53567
rect 35161 53527 35219 53533
rect 20898 53456 20904 53508
rect 20956 53496 20962 53508
rect 21913 53499 21971 53505
rect 21913 53496 21925 53499
rect 20956 53468 21925 53496
rect 20956 53456 20962 53468
rect 21913 53465 21925 53468
rect 21959 53465 21971 53499
rect 21913 53459 21971 53465
rect 29638 53456 29644 53508
rect 29696 53496 29702 53508
rect 35176 53496 35204 53527
rect 36354 53524 36360 53576
rect 36412 53564 36418 53576
rect 36633 53567 36691 53573
rect 36633 53564 36645 53567
rect 36412 53536 36645 53564
rect 36412 53524 36418 53536
rect 36633 53533 36645 53536
rect 36679 53533 36691 53567
rect 36633 53527 36691 53533
rect 38930 53524 38936 53576
rect 38988 53564 38994 53576
rect 39209 53567 39267 53573
rect 39209 53564 39221 53567
rect 38988 53536 39221 53564
rect 38988 53524 38994 53536
rect 39209 53533 39221 53536
rect 39255 53533 39267 53567
rect 39209 53527 39267 53533
rect 44082 53524 44088 53576
rect 44140 53564 44146 53576
rect 44269 53567 44327 53573
rect 44269 53564 44281 53567
rect 44140 53536 44281 53564
rect 44140 53524 44146 53536
rect 44269 53533 44281 53536
rect 44315 53533 44327 53567
rect 44269 53527 44327 53533
rect 46658 53524 46664 53576
rect 46716 53564 46722 53576
rect 46753 53567 46811 53573
rect 46753 53564 46765 53567
rect 46716 53536 46765 53564
rect 46716 53524 46722 53536
rect 46753 53533 46765 53536
rect 46799 53533 46811 53567
rect 46753 53527 46811 53533
rect 48041 53567 48099 53573
rect 48041 53533 48053 53567
rect 48087 53564 48099 53567
rect 48314 53564 48320 53576
rect 48087 53536 48320 53564
rect 48087 53533 48099 53536
rect 48041 53527 48099 53533
rect 48314 53524 48320 53536
rect 48372 53524 48378 53576
rect 48590 53524 48596 53576
rect 48648 53564 48654 53576
rect 48685 53567 48743 53573
rect 48685 53564 48697 53567
rect 48648 53536 48697 53564
rect 48648 53524 48654 53536
rect 48685 53533 48697 53536
rect 48731 53533 48743 53567
rect 48685 53527 48743 53533
rect 29696 53468 35204 53496
rect 29696 53456 29702 53468
rect 37366 53456 37372 53508
rect 37424 53496 37430 53508
rect 37424 53468 45554 53496
rect 37424 53456 37430 53468
rect 22646 53428 22652 53440
rect 17696 53400 22652 53428
rect 22646 53388 22652 53400
rect 22704 53388 22710 53440
rect 22833 53431 22891 53437
rect 22833 53397 22845 53431
rect 22879 53428 22891 53431
rect 23382 53428 23388 53440
rect 22879 53400 23388 53428
rect 22879 53397 22891 53400
rect 22833 53391 22891 53397
rect 23382 53388 23388 53400
rect 23440 53388 23446 53440
rect 28626 53388 28632 53440
rect 28684 53428 28690 53440
rect 28721 53431 28779 53437
rect 28721 53428 28733 53431
rect 28684 53400 28733 53428
rect 28684 53388 28690 53400
rect 28721 53397 28733 53400
rect 28767 53397 28779 53431
rect 28721 53391 28779 53397
rect 30466 53388 30472 53440
rect 30524 53428 30530 53440
rect 31297 53431 31355 53437
rect 31297 53428 31309 53431
rect 30524 53400 31309 53428
rect 30524 53388 30530 53400
rect 31297 53397 31309 53400
rect 31343 53397 31355 53431
rect 31297 53391 31355 53397
rect 31754 53388 31760 53440
rect 31812 53428 31818 53440
rect 33873 53431 33931 53437
rect 33873 53428 33885 53431
rect 31812 53400 33885 53428
rect 31812 53388 31818 53400
rect 33873 53397 33885 53400
rect 33919 53397 33931 53431
rect 33873 53391 33931 53397
rect 39022 53388 39028 53440
rect 39080 53388 39086 53440
rect 45526 53428 45554 53468
rect 46937 53431 46995 53437
rect 46937 53428 46949 53431
rect 45526 53400 46949 53428
rect 46937 53397 46949 53400
rect 46983 53397 46995 53431
rect 46937 53391 46995 53397
rect 48866 53388 48872 53440
rect 48924 53388 48930 53440
rect 1104 53338 49864 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 27950 53338
rect 28002 53286 28014 53338
rect 28066 53286 28078 53338
rect 28130 53286 28142 53338
rect 28194 53286 28206 53338
rect 28258 53286 37950 53338
rect 38002 53286 38014 53338
rect 38066 53286 38078 53338
rect 38130 53286 38142 53338
rect 38194 53286 38206 53338
rect 38258 53286 47950 53338
rect 48002 53286 48014 53338
rect 48066 53286 48078 53338
rect 48130 53286 48142 53338
rect 48194 53286 48206 53338
rect 48258 53286 49864 53338
rect 1104 53264 49864 53286
rect 20714 53184 20720 53236
rect 20772 53224 20778 53236
rect 23293 53227 23351 53233
rect 23293 53224 23305 53227
rect 20772 53196 23305 53224
rect 20772 53184 20778 53196
rect 23293 53193 23305 53196
rect 23339 53193 23351 53227
rect 23293 53187 23351 53193
rect 23566 53184 23572 53236
rect 23624 53224 23630 53236
rect 24029 53227 24087 53233
rect 24029 53224 24041 53227
rect 23624 53196 24041 53224
rect 23624 53184 23630 53196
rect 24029 53193 24041 53196
rect 24075 53193 24087 53227
rect 24029 53187 24087 53193
rect 2222 53116 2228 53168
rect 2280 53156 2286 53168
rect 16206 53156 16212 53168
rect 2280 53128 2820 53156
rect 2280 53116 2286 53128
rect 2501 53091 2559 53097
rect 2501 53057 2513 53091
rect 2547 53057 2559 53091
rect 2501 53051 2559 53057
rect 2516 52952 2544 53051
rect 2792 53029 2820 53128
rect 12820 53128 16212 53156
rect 4709 53091 4767 53097
rect 4709 53057 4721 53091
rect 4755 53088 4767 53091
rect 5810 53088 5816 53100
rect 4755 53060 5816 53088
rect 4755 53057 4767 53060
rect 4709 53051 4767 53057
rect 5810 53048 5816 53060
rect 5868 53048 5874 53100
rect 7009 53091 7067 53097
rect 7009 53057 7021 53091
rect 7055 53057 7067 53091
rect 7009 53051 7067 53057
rect 7653 53091 7711 53097
rect 7653 53057 7665 53091
rect 7699 53088 7711 53091
rect 9674 53088 9680 53100
rect 7699 53060 9680 53088
rect 7699 53057 7711 53060
rect 7653 53051 7711 53057
rect 2777 53023 2835 53029
rect 2777 52989 2789 53023
rect 2823 52989 2835 53023
rect 2777 52983 2835 52989
rect 4798 52980 4804 53032
rect 4856 53020 4862 53032
rect 5077 53023 5135 53029
rect 5077 53020 5089 53023
rect 4856 52992 5089 53020
rect 4856 52980 4862 52992
rect 5077 52989 5089 52992
rect 5123 52989 5135 53023
rect 5077 52983 5135 52989
rect 6825 52955 6883 52961
rect 6825 52952 6837 52955
rect 2516 52924 6837 52952
rect 6825 52921 6837 52924
rect 6871 52921 6883 52955
rect 7024 52952 7052 53051
rect 9674 53048 9680 53060
rect 9732 53048 9738 53100
rect 9861 53091 9919 53097
rect 9861 53057 9873 53091
rect 9907 53088 9919 53091
rect 12434 53088 12440 53100
rect 9907 53060 12440 53088
rect 9907 53057 9919 53060
rect 9861 53051 9919 53057
rect 12434 53048 12440 53060
rect 12492 53048 12498 53100
rect 12820 53097 12848 53128
rect 16206 53116 16212 53128
rect 16264 53116 16270 53168
rect 23201 53159 23259 53165
rect 23201 53125 23213 53159
rect 23247 53156 23259 53159
rect 24854 53156 24860 53168
rect 23247 53128 24860 53156
rect 23247 53125 23259 53128
rect 23201 53119 23259 53125
rect 24854 53116 24860 53128
rect 24912 53116 24918 53168
rect 47762 53116 47768 53168
rect 47820 53156 47826 53168
rect 47857 53159 47915 53165
rect 47857 53156 47869 53159
rect 47820 53128 47869 53156
rect 47820 53116 47826 53128
rect 47857 53125 47869 53128
rect 47903 53125 47915 53159
rect 47857 53119 47915 53125
rect 12805 53091 12863 53097
rect 12805 53057 12817 53091
rect 12851 53057 12863 53091
rect 12805 53051 12863 53057
rect 15013 53091 15071 53097
rect 15013 53057 15025 53091
rect 15059 53088 15071 53091
rect 15286 53088 15292 53100
rect 15059 53060 15292 53088
rect 15059 53057 15071 53060
rect 15013 53051 15071 53057
rect 15286 53048 15292 53060
rect 15344 53048 15350 53100
rect 17865 53091 17923 53097
rect 17865 53057 17877 53091
rect 17911 53088 17923 53091
rect 19334 53088 19340 53100
rect 17911 53060 19340 53088
rect 17911 53057 17923 53060
rect 17865 53051 17923 53057
rect 19334 53048 19340 53060
rect 19392 53048 19398 53100
rect 19886 53048 19892 53100
rect 19944 53048 19950 53100
rect 21542 53048 21548 53100
rect 21600 53088 21606 53100
rect 22189 53091 22247 53097
rect 22189 53088 22201 53091
rect 21600 53060 22201 53088
rect 21600 53048 21606 53060
rect 22189 53057 22201 53060
rect 22235 53057 22247 53091
rect 22189 53051 22247 53057
rect 23937 53091 23995 53097
rect 23937 53057 23949 53091
rect 23983 53088 23995 53091
rect 27338 53088 27344 53100
rect 23983 53060 27344 53088
rect 23983 53057 23995 53060
rect 23937 53051 23995 53057
rect 27338 53048 27344 53060
rect 27396 53048 27402 53100
rect 48777 53091 48835 53097
rect 48777 53088 48789 53091
rect 47964 53060 48789 53088
rect 7374 52980 7380 53032
rect 7432 53020 7438 53032
rect 7929 53023 7987 53029
rect 7929 53020 7941 53023
rect 7432 52992 7941 53020
rect 7432 52980 7438 52992
rect 7929 52989 7941 52992
rect 7975 52989 7987 53023
rect 7929 52983 7987 52989
rect 9950 52980 9956 53032
rect 10008 53020 10014 53032
rect 10229 53023 10287 53029
rect 10229 53020 10241 53023
rect 10008 52992 10241 53020
rect 10008 52980 10014 52992
rect 10229 52989 10241 52992
rect 10275 52989 10287 53023
rect 10229 52983 10287 52989
rect 12526 52980 12532 53032
rect 12584 53020 12590 53032
rect 13081 53023 13139 53029
rect 13081 53020 13093 53023
rect 12584 52992 13093 53020
rect 12584 52980 12590 52992
rect 13081 52989 13093 52992
rect 13127 52989 13139 53023
rect 13081 52983 13139 52989
rect 15102 52980 15108 53032
rect 15160 53020 15166 53032
rect 15381 53023 15439 53029
rect 15381 53020 15393 53023
rect 15160 52992 15393 53020
rect 15160 52980 15166 52992
rect 15381 52989 15393 52992
rect 15427 52989 15439 53023
rect 15381 52983 15439 52989
rect 17678 52980 17684 53032
rect 17736 53020 17742 53032
rect 18233 53023 18291 53029
rect 18233 53020 18245 53023
rect 17736 52992 18245 53020
rect 17736 52980 17742 52992
rect 18233 52989 18245 52992
rect 18279 52989 18291 53023
rect 18233 52983 18291 52989
rect 19610 52980 19616 53032
rect 19668 53020 19674 53032
rect 20165 53023 20223 53029
rect 20165 53020 20177 53023
rect 19668 52992 20177 53020
rect 19668 52980 19674 52992
rect 20165 52989 20177 52992
rect 20211 52989 20223 53023
rect 20165 52983 20223 52989
rect 33686 52980 33692 53032
rect 33744 53020 33750 53032
rect 47964 53020 47992 53060
rect 48777 53057 48789 53060
rect 48823 53057 48835 53091
rect 48777 53051 48835 53057
rect 33744 52992 47992 53020
rect 33744 52980 33750 52992
rect 48498 52980 48504 53032
rect 48556 52980 48562 53032
rect 12802 52952 12808 52964
rect 7024 52924 12808 52952
rect 6825 52915 6883 52921
rect 12802 52912 12808 52924
rect 12860 52912 12866 52964
rect 22005 52887 22063 52893
rect 22005 52853 22017 52887
rect 22051 52884 22063 52887
rect 25314 52884 25320 52896
rect 22051 52856 25320 52884
rect 22051 52853 22063 52856
rect 22005 52847 22063 52853
rect 25314 52844 25320 52856
rect 25372 52844 25378 52896
rect 46198 52844 46204 52896
rect 46256 52884 46262 52896
rect 47949 52887 48007 52893
rect 47949 52884 47961 52887
rect 46256 52856 47961 52884
rect 46256 52844 46262 52856
rect 47949 52853 47961 52856
rect 47995 52853 48007 52887
rect 47949 52847 48007 52853
rect 1104 52794 49864 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 32950 52794
rect 33002 52742 33014 52794
rect 33066 52742 33078 52794
rect 33130 52742 33142 52794
rect 33194 52742 33206 52794
rect 33258 52742 42950 52794
rect 43002 52742 43014 52794
rect 43066 52742 43078 52794
rect 43130 52742 43142 52794
rect 43194 52742 43206 52794
rect 43258 52742 49864 52794
rect 1104 52720 49864 52742
rect 19886 52640 19892 52692
rect 19944 52680 19950 52692
rect 22557 52683 22615 52689
rect 22557 52680 22569 52683
rect 19944 52652 22569 52680
rect 19944 52640 19950 52652
rect 22557 52649 22569 52652
rect 22603 52649 22615 52683
rect 22557 52643 22615 52649
rect 22646 52640 22652 52692
rect 22704 52680 22710 52692
rect 23385 52683 23443 52689
rect 23385 52680 23397 52683
rect 22704 52652 23397 52680
rect 22704 52640 22710 52652
rect 23385 52649 23397 52652
rect 23431 52649 23443 52683
rect 23385 52643 23443 52649
rect 15378 52572 15384 52624
rect 15436 52612 15442 52624
rect 20257 52615 20315 52621
rect 20257 52612 20269 52615
rect 15436 52584 20269 52612
rect 15436 52572 15442 52584
rect 20257 52581 20269 52584
rect 20303 52581 20315 52615
rect 20257 52575 20315 52581
rect 1578 52504 1584 52556
rect 1636 52544 1642 52556
rect 2133 52547 2191 52553
rect 2133 52544 2145 52547
rect 1636 52516 2145 52544
rect 1636 52504 1642 52516
rect 2133 52513 2145 52516
rect 2179 52513 2191 52547
rect 2133 52507 2191 52513
rect 4154 52504 4160 52556
rect 4212 52544 4218 52556
rect 4801 52547 4859 52553
rect 4801 52544 4813 52547
rect 4212 52516 4813 52544
rect 4212 52504 4218 52516
rect 4801 52513 4813 52516
rect 4847 52513 4859 52547
rect 4801 52507 4859 52513
rect 6730 52504 6736 52556
rect 6788 52544 6794 52556
rect 7285 52547 7343 52553
rect 7285 52544 7297 52547
rect 6788 52516 7297 52544
rect 6788 52504 6794 52516
rect 7285 52513 7297 52516
rect 7331 52513 7343 52547
rect 7285 52507 7343 52513
rect 9306 52504 9312 52556
rect 9364 52544 9370 52556
rect 9861 52547 9919 52553
rect 9861 52544 9873 52547
rect 9364 52516 9873 52544
rect 9364 52504 9370 52516
rect 9861 52513 9873 52516
rect 9907 52513 9919 52547
rect 9861 52507 9919 52513
rect 11882 52504 11888 52556
rect 11940 52544 11946 52556
rect 12437 52547 12495 52553
rect 12437 52544 12449 52547
rect 11940 52516 12449 52544
rect 11940 52504 11946 52516
rect 12437 52513 12449 52516
rect 12483 52513 12495 52547
rect 12437 52507 12495 52513
rect 14458 52504 14464 52556
rect 14516 52544 14522 52556
rect 15013 52547 15071 52553
rect 15013 52544 15025 52547
rect 14516 52516 15025 52544
rect 14516 52504 14522 52516
rect 15013 52513 15025 52516
rect 15059 52513 15071 52547
rect 15013 52507 15071 52513
rect 17034 52504 17040 52556
rect 17092 52544 17098 52556
rect 17589 52547 17647 52553
rect 17589 52544 17601 52547
rect 17092 52516 17601 52544
rect 17092 52504 17098 52516
rect 17589 52513 17601 52516
rect 17635 52513 17647 52547
rect 24762 52544 24768 52556
rect 17589 52507 17647 52513
rect 22756 52516 24768 52544
rect 1670 52436 1676 52488
rect 1728 52436 1734 52488
rect 4433 52479 4491 52485
rect 4433 52445 4445 52479
rect 4479 52476 4491 52479
rect 4706 52476 4712 52488
rect 4479 52448 4712 52476
rect 4479 52445 4491 52448
rect 4433 52439 4491 52445
rect 4706 52436 4712 52448
rect 4764 52436 4770 52488
rect 7009 52479 7067 52485
rect 7009 52445 7021 52479
rect 7055 52476 7067 52479
rect 8294 52476 8300 52488
rect 7055 52448 8300 52476
rect 7055 52445 7067 52448
rect 7009 52439 7067 52445
rect 8294 52436 8300 52448
rect 8352 52436 8358 52488
rect 9585 52479 9643 52485
rect 9585 52445 9597 52479
rect 9631 52476 9643 52479
rect 9766 52476 9772 52488
rect 9631 52448 9772 52476
rect 9631 52445 9643 52448
rect 9585 52439 9643 52445
rect 9766 52436 9772 52448
rect 9824 52436 9830 52488
rect 12161 52479 12219 52485
rect 12161 52445 12173 52479
rect 12207 52476 12219 52479
rect 13814 52476 13820 52488
rect 12207 52448 13820 52476
rect 12207 52445 12219 52448
rect 12161 52439 12219 52445
rect 13814 52436 13820 52448
rect 13872 52436 13878 52488
rect 14737 52479 14795 52485
rect 14737 52445 14749 52479
rect 14783 52476 14795 52479
rect 16850 52476 16856 52488
rect 14783 52448 16856 52476
rect 14783 52445 14795 52448
rect 14737 52439 14795 52445
rect 16850 52436 16856 52448
rect 16908 52436 16914 52488
rect 17313 52479 17371 52485
rect 17313 52445 17325 52479
rect 17359 52476 17371 52479
rect 19426 52476 19432 52488
rect 17359 52448 19432 52476
rect 17359 52445 17371 52448
rect 17313 52439 17371 52445
rect 19426 52436 19432 52448
rect 19484 52436 19490 52488
rect 22756 52485 22784 52516
rect 24762 52504 24768 52516
rect 24820 52504 24826 52556
rect 36354 52504 36360 52556
rect 36412 52544 36418 52556
rect 48777 52547 48835 52553
rect 48777 52544 48789 52547
rect 36412 52516 48789 52544
rect 36412 52504 36418 52516
rect 48777 52513 48789 52516
rect 48823 52513 48835 52547
rect 48777 52507 48835 52513
rect 22741 52479 22799 52485
rect 22741 52445 22753 52479
rect 22787 52445 22799 52479
rect 48041 52479 48099 52485
rect 22741 52439 22799 52445
rect 23216 52448 23428 52476
rect 20073 52411 20131 52417
rect 20073 52377 20085 52411
rect 20119 52408 20131 52411
rect 23216 52408 23244 52448
rect 20119 52380 23244 52408
rect 23293 52411 23351 52417
rect 20119 52377 20131 52380
rect 20073 52371 20131 52377
rect 23293 52377 23305 52411
rect 23339 52377 23351 52411
rect 23400 52408 23428 52448
rect 48041 52445 48053 52479
rect 48087 52476 48099 52479
rect 48498 52476 48504 52488
rect 48087 52448 48504 52476
rect 48087 52445 48099 52448
rect 48041 52439 48099 52445
rect 48498 52436 48504 52448
rect 48556 52436 48562 52488
rect 35526 52408 35532 52420
rect 23400 52380 35532 52408
rect 23293 52371 23351 52377
rect 23308 52340 23336 52371
rect 35526 52368 35532 52380
rect 35584 52368 35590 52420
rect 24946 52340 24952 52352
rect 23308 52312 24952 52340
rect 24946 52300 24952 52312
rect 25004 52300 25010 52352
rect 1104 52250 49864 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 27950 52250
rect 28002 52198 28014 52250
rect 28066 52198 28078 52250
rect 28130 52198 28142 52250
rect 28194 52198 28206 52250
rect 28258 52198 37950 52250
rect 38002 52198 38014 52250
rect 38066 52198 38078 52250
rect 38130 52198 38142 52250
rect 38194 52198 38206 52250
rect 38258 52198 47950 52250
rect 48002 52198 48014 52250
rect 48066 52198 48078 52250
rect 48130 52198 48142 52250
rect 48194 52198 48206 52250
rect 48258 52198 49864 52250
rect 1104 52176 49864 52198
rect 5810 52096 5816 52148
rect 5868 52136 5874 52148
rect 8481 52139 8539 52145
rect 8481 52136 8493 52139
rect 5868 52108 8493 52136
rect 5868 52096 5874 52108
rect 8481 52105 8493 52108
rect 8527 52105 8539 52139
rect 8481 52099 8539 52105
rect 8389 52003 8447 52009
rect 8389 51969 8401 52003
rect 8435 52000 8447 52003
rect 10686 52000 10692 52012
rect 8435 51972 10692 52000
rect 8435 51969 8447 51972
rect 8389 51963 8447 51969
rect 10686 51960 10692 51972
rect 10744 51960 10750 52012
rect 49234 51960 49240 52012
rect 49292 52000 49298 52012
rect 49329 52003 49387 52009
rect 49329 52000 49341 52003
rect 49292 51972 49341 52000
rect 49292 51960 49298 51972
rect 49329 51969 49341 51972
rect 49375 51969 49387 52003
rect 49329 51963 49387 51969
rect 38930 51756 38936 51808
rect 38988 51796 38994 51808
rect 43438 51796 43444 51808
rect 38988 51768 43444 51796
rect 38988 51756 38994 51768
rect 43438 51756 43444 51768
rect 43496 51756 43502 51808
rect 49142 51756 49148 51808
rect 49200 51756 49206 51808
rect 1104 51706 49864 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 32950 51706
rect 33002 51654 33014 51706
rect 33066 51654 33078 51706
rect 33130 51654 33142 51706
rect 33194 51654 33206 51706
rect 33258 51654 42950 51706
rect 43002 51654 43014 51706
rect 43066 51654 43078 51706
rect 43130 51654 43142 51706
rect 43194 51654 43206 51706
rect 43258 51654 49864 51706
rect 1104 51632 49864 51654
rect 4890 51552 4896 51604
rect 4948 51592 4954 51604
rect 9309 51595 9367 51601
rect 9309 51592 9321 51595
rect 4948 51564 9321 51592
rect 4948 51552 4954 51564
rect 9309 51561 9321 51564
rect 9355 51561 9367 51595
rect 9309 51555 9367 51561
rect 42150 51552 42156 51604
rect 42208 51592 42214 51604
rect 43898 51592 43904 51604
rect 42208 51564 43904 51592
rect 42208 51552 42214 51564
rect 43898 51552 43904 51564
rect 43956 51552 43962 51604
rect 1302 51416 1308 51468
rect 1360 51456 1366 51468
rect 2041 51459 2099 51465
rect 2041 51456 2053 51459
rect 1360 51428 2053 51456
rect 1360 51416 1366 51428
rect 2041 51425 2053 51428
rect 2087 51425 2099 51459
rect 2041 51419 2099 51425
rect 41693 51459 41751 51465
rect 41693 51425 41705 51459
rect 41739 51456 41751 51459
rect 49142 51456 49148 51468
rect 41739 51428 49148 51456
rect 41739 51425 41751 51428
rect 41693 51419 41751 51425
rect 49142 51416 49148 51428
rect 49200 51416 49206 51468
rect 1765 51391 1823 51397
rect 1765 51357 1777 51391
rect 1811 51388 1823 51391
rect 7558 51388 7564 51400
rect 1811 51360 7564 51388
rect 1811 51357 1823 51360
rect 1765 51351 1823 51357
rect 7558 51348 7564 51360
rect 7616 51348 7622 51400
rect 37274 51348 37280 51400
rect 37332 51388 37338 51400
rect 41417 51391 41475 51397
rect 41417 51388 41429 51391
rect 37332 51360 41429 51388
rect 37332 51348 37338 51360
rect 41417 51357 41429 51360
rect 41463 51357 41475 51391
rect 41417 51351 41475 51357
rect 43438 51348 43444 51400
rect 43496 51348 43502 51400
rect 48498 51348 48504 51400
rect 48556 51348 48562 51400
rect 48777 51391 48835 51397
rect 48777 51357 48789 51391
rect 48823 51357 48835 51391
rect 48777 51351 48835 51357
rect 9217 51323 9275 51329
rect 9217 51289 9229 51323
rect 9263 51320 9275 51323
rect 10962 51320 10968 51332
rect 9263 51292 10968 51320
rect 9263 51289 9275 51292
rect 9217 51283 9275 51289
rect 10962 51280 10968 51292
rect 11020 51280 11026 51332
rect 39298 51280 39304 51332
rect 39356 51320 39362 51332
rect 42150 51320 42156 51332
rect 39356 51292 42156 51320
rect 39356 51280 39362 51292
rect 42150 51280 42156 51292
rect 42208 51280 42214 51332
rect 23934 51212 23940 51264
rect 23992 51252 23998 51264
rect 48792 51252 48820 51351
rect 23992 51224 48820 51252
rect 23992 51212 23998 51224
rect 1104 51162 49864 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 27950 51162
rect 28002 51110 28014 51162
rect 28066 51110 28078 51162
rect 28130 51110 28142 51162
rect 28194 51110 28206 51162
rect 28258 51110 37950 51162
rect 38002 51110 38014 51162
rect 38066 51110 38078 51162
rect 38130 51110 38142 51162
rect 38194 51110 38206 51162
rect 38258 51110 47950 51162
rect 48002 51110 48014 51162
rect 48066 51110 48078 51162
rect 48130 51110 48142 51162
rect 48194 51110 48206 51162
rect 48258 51110 49864 51162
rect 1104 51088 49864 51110
rect 8294 51008 8300 51060
rect 8352 51048 8358 51060
rect 9309 51051 9367 51057
rect 9309 51048 9321 51051
rect 8352 51020 9321 51048
rect 8352 51008 8358 51020
rect 9309 51017 9321 51020
rect 9355 51017 9367 51051
rect 9309 51011 9367 51017
rect 9674 51008 9680 51060
rect 9732 51048 9738 51060
rect 10137 51051 10195 51057
rect 10137 51048 10149 51051
rect 9732 51020 10149 51048
rect 9732 51008 9738 51020
rect 10137 51017 10149 51020
rect 10183 51017 10195 51051
rect 10137 51011 10195 51017
rect 10502 51008 10508 51060
rect 10560 51048 10566 51060
rect 13449 51051 13507 51057
rect 13449 51048 13461 51051
rect 10560 51020 13461 51048
rect 10560 51008 10566 51020
rect 13449 51017 13461 51020
rect 13495 51017 13507 51051
rect 13449 51011 13507 51017
rect 15194 51008 15200 51060
rect 15252 51048 15258 51060
rect 17037 51051 17095 51057
rect 17037 51048 17049 51051
rect 15252 51020 17049 51048
rect 15252 51008 15258 51020
rect 17037 51017 17049 51020
rect 17083 51017 17095 51051
rect 17037 51011 17095 51017
rect 19334 51008 19340 51060
rect 19392 51048 19398 51060
rect 22189 51051 22247 51057
rect 22189 51048 22201 51051
rect 19392 51020 22201 51048
rect 19392 51008 19398 51020
rect 22189 51017 22201 51020
rect 22235 51017 22247 51051
rect 22189 51011 22247 51017
rect 26234 51008 26240 51060
rect 26292 51008 26298 51060
rect 27338 51008 27344 51060
rect 27396 51008 27402 51060
rect 31481 50983 31539 50989
rect 31481 50949 31493 50983
rect 31527 50980 31539 50983
rect 35158 50980 35164 50992
rect 31527 50952 35164 50980
rect 31527 50949 31539 50952
rect 31481 50943 31539 50949
rect 35158 50940 35164 50952
rect 35216 50940 35222 50992
rect 1765 50915 1823 50921
rect 1765 50881 1777 50915
rect 1811 50912 1823 50915
rect 5626 50912 5632 50924
rect 1811 50884 5632 50912
rect 1811 50881 1823 50884
rect 1765 50875 1823 50881
rect 5626 50872 5632 50884
rect 5684 50872 5690 50924
rect 9217 50915 9275 50921
rect 9217 50881 9229 50915
rect 9263 50912 9275 50915
rect 9950 50912 9956 50924
rect 9263 50884 9956 50912
rect 9263 50881 9275 50884
rect 9217 50875 9275 50881
rect 9950 50872 9956 50884
rect 10008 50872 10014 50924
rect 10045 50915 10103 50921
rect 10045 50881 10057 50915
rect 10091 50912 10103 50915
rect 11606 50912 11612 50924
rect 10091 50884 11612 50912
rect 10091 50881 10103 50884
rect 10045 50875 10103 50881
rect 11606 50872 11612 50884
rect 11664 50872 11670 50924
rect 13357 50915 13415 50921
rect 13357 50881 13369 50915
rect 13403 50912 13415 50915
rect 14918 50912 14924 50924
rect 13403 50884 14924 50912
rect 13403 50881 13415 50884
rect 13357 50875 13415 50881
rect 14918 50872 14924 50884
rect 14976 50872 14982 50924
rect 16945 50915 17003 50921
rect 16945 50881 16957 50915
rect 16991 50912 17003 50915
rect 19242 50912 19248 50924
rect 16991 50884 19248 50912
rect 16991 50881 17003 50884
rect 16945 50875 17003 50881
rect 19242 50872 19248 50884
rect 19300 50872 19306 50924
rect 22097 50915 22155 50921
rect 22097 50881 22109 50915
rect 22143 50912 22155 50915
rect 24486 50912 24492 50924
rect 22143 50884 24492 50912
rect 22143 50881 22155 50884
rect 22097 50875 22155 50881
rect 24486 50872 24492 50884
rect 24544 50872 24550 50924
rect 26421 50915 26479 50921
rect 26421 50881 26433 50915
rect 26467 50881 26479 50915
rect 26421 50875 26479 50881
rect 1302 50804 1308 50856
rect 1360 50844 1366 50856
rect 2041 50847 2099 50853
rect 2041 50844 2053 50847
rect 1360 50816 2053 50844
rect 1360 50804 1366 50816
rect 2041 50813 2053 50816
rect 2087 50813 2099 50847
rect 26436 50844 26464 50875
rect 27522 50872 27528 50924
rect 27580 50872 27586 50924
rect 28261 50915 28319 50921
rect 28261 50881 28273 50915
rect 28307 50912 28319 50915
rect 31294 50912 31300 50924
rect 28307 50884 31300 50912
rect 28307 50881 28319 50884
rect 28261 50875 28319 50881
rect 31294 50872 31300 50884
rect 31352 50872 31358 50924
rect 31389 50915 31447 50921
rect 31389 50881 31401 50915
rect 31435 50912 31447 50915
rect 32306 50912 32312 50924
rect 31435 50884 32312 50912
rect 31435 50881 31447 50884
rect 31389 50875 31447 50881
rect 32306 50872 32312 50884
rect 32364 50872 32370 50924
rect 49326 50872 49332 50924
rect 49384 50872 49390 50924
rect 28902 50844 28908 50856
rect 26436 50816 28908 50844
rect 2041 50807 2099 50813
rect 28902 50804 28908 50816
rect 28960 50804 28966 50856
rect 29086 50804 29092 50856
rect 29144 50844 29150 50856
rect 31573 50847 31631 50853
rect 31573 50844 31585 50847
rect 29144 50816 31585 50844
rect 29144 50804 29150 50816
rect 31573 50813 31585 50816
rect 31619 50813 31631 50847
rect 31573 50807 31631 50813
rect 24854 50736 24860 50788
rect 24912 50776 24918 50788
rect 28077 50779 28135 50785
rect 28077 50776 28089 50779
rect 24912 50748 28089 50776
rect 24912 50736 24918 50748
rect 28077 50745 28089 50748
rect 28123 50745 28135 50779
rect 28077 50739 28135 50745
rect 28184 50748 31616 50776
rect 26694 50668 26700 50720
rect 26752 50708 26758 50720
rect 28184 50708 28212 50748
rect 31588 50720 31616 50748
rect 26752 50680 28212 50708
rect 26752 50668 26758 50680
rect 30374 50668 30380 50720
rect 30432 50708 30438 50720
rect 30558 50708 30564 50720
rect 30432 50680 30564 50708
rect 30432 50668 30438 50680
rect 30558 50668 30564 50680
rect 30616 50668 30622 50720
rect 31018 50668 31024 50720
rect 31076 50668 31082 50720
rect 31570 50668 31576 50720
rect 31628 50668 31634 50720
rect 42794 50668 42800 50720
rect 42852 50708 42858 50720
rect 49145 50711 49203 50717
rect 49145 50708 49157 50711
rect 42852 50680 49157 50708
rect 42852 50668 42858 50680
rect 49145 50677 49157 50680
rect 49191 50677 49203 50711
rect 49145 50671 49203 50677
rect 1104 50618 49864 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 32950 50618
rect 33002 50566 33014 50618
rect 33066 50566 33078 50618
rect 33130 50566 33142 50618
rect 33194 50566 33206 50618
rect 33258 50566 42950 50618
rect 43002 50566 43014 50618
rect 43066 50566 43078 50618
rect 43130 50566 43142 50618
rect 43194 50566 43206 50618
rect 43258 50566 49864 50618
rect 1104 50544 49864 50566
rect 12434 50464 12440 50516
rect 12492 50504 12498 50516
rect 13449 50507 13507 50513
rect 13449 50504 13461 50507
rect 12492 50476 13461 50504
rect 12492 50464 12498 50476
rect 13449 50473 13461 50476
rect 13495 50473 13507 50507
rect 13449 50467 13507 50473
rect 16850 50464 16856 50516
rect 16908 50504 16914 50516
rect 17589 50507 17647 50513
rect 17589 50504 17601 50507
rect 16908 50476 17601 50504
rect 16908 50464 16914 50476
rect 17589 50473 17601 50476
rect 17635 50473 17647 50507
rect 17589 50467 17647 50473
rect 19426 50464 19432 50516
rect 19484 50504 19490 50516
rect 22649 50507 22707 50513
rect 22649 50504 22661 50507
rect 19484 50476 22661 50504
rect 19484 50464 19490 50476
rect 22649 50473 22661 50476
rect 22695 50473 22707 50507
rect 22649 50467 22707 50473
rect 27522 50464 27528 50516
rect 27580 50504 27586 50516
rect 31113 50507 31171 50513
rect 31113 50504 31125 50507
rect 27580 50476 31125 50504
rect 27580 50464 27586 50476
rect 31113 50473 31125 50476
rect 31159 50473 31171 50507
rect 31113 50467 31171 50473
rect 32306 50464 32312 50516
rect 32364 50504 32370 50516
rect 32950 50504 32956 50516
rect 32364 50476 32956 50504
rect 32364 50464 32370 50476
rect 32950 50464 32956 50476
rect 33008 50464 33014 50516
rect 8386 50396 8392 50448
rect 8444 50396 8450 50448
rect 13722 50396 13728 50448
rect 13780 50436 13786 50448
rect 16945 50439 17003 50445
rect 16945 50436 16957 50439
rect 13780 50408 16957 50436
rect 13780 50396 13786 50408
rect 16945 50405 16957 50408
rect 16991 50405 17003 50439
rect 16945 50399 17003 50405
rect 27614 50396 27620 50448
rect 27672 50436 27678 50448
rect 29917 50439 29975 50445
rect 29917 50436 29929 50439
rect 27672 50408 29929 50436
rect 27672 50396 27678 50408
rect 29917 50405 29929 50408
rect 29963 50405 29975 50439
rect 29917 50399 29975 50405
rect 30006 50396 30012 50448
rect 30064 50436 30070 50448
rect 35250 50436 35256 50448
rect 30064 50408 30512 50436
rect 30064 50396 30070 50408
rect 13814 50328 13820 50380
rect 13872 50368 13878 50380
rect 15102 50368 15108 50380
rect 13872 50340 15108 50368
rect 13872 50328 13878 50340
rect 15102 50328 15108 50340
rect 15160 50328 15166 50380
rect 25866 50328 25872 50380
rect 25924 50368 25930 50380
rect 30484 50377 30512 50408
rect 31036 50408 35256 50436
rect 28353 50371 28411 50377
rect 28353 50368 28365 50371
rect 25924 50340 28365 50368
rect 25924 50328 25930 50340
rect 28353 50337 28365 50340
rect 28399 50337 28411 50371
rect 28353 50331 28411 50337
rect 30469 50371 30527 50377
rect 30469 50337 30481 50371
rect 30515 50337 30527 50371
rect 30469 50331 30527 50337
rect 16761 50303 16819 50309
rect 16761 50269 16773 50303
rect 16807 50300 16819 50303
rect 18322 50300 18328 50312
rect 16807 50272 18328 50300
rect 16807 50269 16819 50272
rect 16761 50263 16819 50269
rect 18322 50260 18328 50272
rect 18380 50260 18386 50312
rect 28169 50303 28227 50309
rect 28169 50269 28181 50303
rect 28215 50300 28227 50303
rect 30558 50300 30564 50312
rect 28215 50272 30564 50300
rect 28215 50269 28227 50272
rect 28169 50263 28227 50269
rect 30558 50260 30564 50272
rect 30616 50260 30622 50312
rect 8205 50235 8263 50241
rect 8205 50201 8217 50235
rect 8251 50232 8263 50235
rect 9582 50232 9588 50244
rect 8251 50204 9588 50232
rect 8251 50201 8263 50204
rect 8205 50195 8263 50201
rect 9582 50192 9588 50204
rect 9640 50192 9646 50244
rect 13357 50235 13415 50241
rect 13357 50201 13369 50235
rect 13403 50232 13415 50235
rect 14826 50232 14832 50244
rect 13403 50204 14832 50232
rect 13403 50201 13415 50204
rect 13357 50195 13415 50201
rect 14826 50192 14832 50204
rect 14884 50192 14890 50244
rect 17494 50192 17500 50244
rect 17552 50192 17558 50244
rect 22557 50235 22615 50241
rect 22557 50201 22569 50235
rect 22603 50232 22615 50235
rect 25590 50232 25596 50244
rect 22603 50204 25596 50232
rect 22603 50201 22615 50204
rect 22557 50195 22615 50201
rect 25590 50192 25596 50204
rect 25648 50192 25654 50244
rect 30650 50232 30656 50244
rect 28276 50204 30656 50232
rect 22462 50124 22468 50176
rect 22520 50164 22526 50176
rect 28276 50173 28304 50204
rect 30650 50192 30656 50204
rect 30708 50192 30714 50244
rect 27801 50167 27859 50173
rect 27801 50164 27813 50167
rect 22520 50136 27813 50164
rect 22520 50124 22526 50136
rect 27801 50133 27813 50136
rect 27847 50133 27859 50167
rect 27801 50127 27859 50133
rect 28261 50167 28319 50173
rect 28261 50133 28273 50167
rect 28307 50133 28319 50167
rect 28261 50127 28319 50133
rect 30282 50124 30288 50176
rect 30340 50124 30346 50176
rect 30377 50167 30435 50173
rect 30377 50133 30389 50167
rect 30423 50164 30435 50167
rect 31036 50164 31064 50408
rect 35250 50396 35256 50408
rect 35308 50396 35314 50448
rect 31757 50371 31815 50377
rect 31757 50337 31769 50371
rect 31803 50368 31815 50371
rect 33502 50368 33508 50380
rect 31803 50340 33508 50368
rect 31803 50337 31815 50340
rect 31757 50331 31815 50337
rect 33502 50328 33508 50340
rect 33560 50328 33566 50380
rect 31662 50192 31668 50244
rect 31720 50232 31726 50244
rect 34514 50232 34520 50244
rect 31720 50204 34520 50232
rect 31720 50192 31726 50204
rect 34514 50192 34520 50204
rect 34572 50192 34578 50244
rect 30423 50136 31064 50164
rect 30423 50133 30435 50136
rect 30377 50127 30435 50133
rect 31110 50124 31116 50176
rect 31168 50164 31174 50176
rect 31481 50167 31539 50173
rect 31481 50164 31493 50167
rect 31168 50136 31493 50164
rect 31168 50124 31174 50136
rect 31481 50133 31493 50136
rect 31527 50133 31539 50167
rect 31481 50127 31539 50133
rect 31573 50167 31631 50173
rect 31573 50133 31585 50167
rect 31619 50164 31631 50167
rect 34422 50164 34428 50176
rect 31619 50136 34428 50164
rect 31619 50133 31631 50136
rect 31573 50127 31631 50133
rect 34422 50124 34428 50136
rect 34480 50124 34486 50176
rect 1104 50074 49864 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 27950 50074
rect 28002 50022 28014 50074
rect 28066 50022 28078 50074
rect 28130 50022 28142 50074
rect 28194 50022 28206 50074
rect 28258 50022 37950 50074
rect 38002 50022 38014 50074
rect 38066 50022 38078 50074
rect 38130 50022 38142 50074
rect 38194 50022 38206 50074
rect 38258 50022 47950 50074
rect 48002 50022 48014 50074
rect 48066 50022 48078 50074
rect 48130 50022 48142 50074
rect 48194 50022 48206 50074
rect 48258 50022 49864 50074
rect 1104 50000 49864 50022
rect 12802 49920 12808 49972
rect 12860 49960 12866 49972
rect 13265 49963 13323 49969
rect 13265 49960 13277 49963
rect 12860 49932 13277 49960
rect 12860 49920 12866 49932
rect 13265 49929 13277 49932
rect 13311 49929 13323 49963
rect 13265 49923 13323 49929
rect 13538 49920 13544 49972
rect 13596 49960 13602 49972
rect 14093 49963 14151 49969
rect 14093 49960 14105 49963
rect 13596 49932 14105 49960
rect 13596 49920 13602 49932
rect 14093 49929 14105 49932
rect 14139 49929 14151 49963
rect 16114 49960 16120 49972
rect 14093 49923 14151 49929
rect 14844 49932 16120 49960
rect 1765 49827 1823 49833
rect 1765 49793 1777 49827
rect 1811 49824 1823 49827
rect 5718 49824 5724 49836
rect 1811 49796 5724 49824
rect 1811 49793 1823 49796
rect 1765 49787 1823 49793
rect 5718 49784 5724 49796
rect 5776 49784 5782 49836
rect 13449 49827 13507 49833
rect 13449 49793 13461 49827
rect 13495 49793 13507 49827
rect 13449 49787 13507 49793
rect 14001 49827 14059 49833
rect 14001 49793 14013 49827
rect 14047 49824 14059 49827
rect 14844 49824 14872 49932
rect 16114 49920 16120 49932
rect 16172 49920 16178 49972
rect 16206 49920 16212 49972
rect 16264 49920 16270 49972
rect 22094 49920 22100 49972
rect 22152 49960 22158 49972
rect 22189 49963 22247 49969
rect 22189 49960 22201 49963
rect 22152 49932 22201 49960
rect 22152 49920 22158 49932
rect 22189 49929 22201 49932
rect 22235 49929 22247 49963
rect 22189 49923 22247 49929
rect 26326 49920 26332 49972
rect 26384 49960 26390 49972
rect 29825 49963 29883 49969
rect 29825 49960 29837 49963
rect 26384 49932 29837 49960
rect 26384 49920 26390 49932
rect 29825 49929 29837 49932
rect 29871 49929 29883 49963
rect 31021 49963 31079 49969
rect 31021 49960 31033 49963
rect 29825 49923 29883 49929
rect 29932 49932 31033 49960
rect 15102 49852 15108 49904
rect 15160 49852 15166 49904
rect 21453 49895 21511 49901
rect 21453 49892 21465 49895
rect 15212 49864 21465 49892
rect 14047 49796 14872 49824
rect 14921 49827 14979 49833
rect 14047 49793 14059 49796
rect 14001 49787 14059 49793
rect 14921 49793 14933 49827
rect 14967 49793 14979 49827
rect 14921 49787 14979 49793
rect 1302 49716 1308 49768
rect 1360 49756 1366 49768
rect 2041 49759 2099 49765
rect 2041 49756 2053 49759
rect 1360 49728 2053 49756
rect 1360 49716 1366 49728
rect 2041 49725 2053 49728
rect 2087 49725 2099 49759
rect 13464 49756 13492 49787
rect 13464 49728 14872 49756
rect 2041 49719 2099 49725
rect 14844 49620 14872 49728
rect 14936 49688 14964 49787
rect 15010 49784 15016 49836
rect 15068 49824 15074 49836
rect 15212 49824 15240 49864
rect 21453 49861 21465 49864
rect 21499 49861 21511 49895
rect 21453 49855 21511 49861
rect 15068 49796 15240 49824
rect 16117 49827 16175 49833
rect 15068 49784 15074 49796
rect 16117 49793 16129 49827
rect 16163 49824 16175 49827
rect 18966 49824 18972 49836
rect 16163 49796 18972 49824
rect 16163 49793 16175 49796
rect 16117 49787 16175 49793
rect 18966 49784 18972 49796
rect 19024 49784 19030 49836
rect 21269 49827 21327 49833
rect 21269 49793 21281 49827
rect 21315 49824 21327 49827
rect 21910 49824 21916 49836
rect 21315 49796 21916 49824
rect 21315 49793 21327 49796
rect 21269 49787 21327 49793
rect 21910 49784 21916 49796
rect 21968 49784 21974 49836
rect 22097 49827 22155 49833
rect 22097 49793 22109 49827
rect 22143 49824 22155 49827
rect 26602 49824 26608 49836
rect 22143 49796 26608 49824
rect 22143 49793 22155 49796
rect 22097 49787 22155 49793
rect 26602 49784 26608 49796
rect 26660 49784 26666 49836
rect 28994 49784 29000 49836
rect 29052 49784 29058 49836
rect 27614 49716 27620 49768
rect 27672 49716 27678 49768
rect 29932 49756 29960 49932
rect 31021 49929 31033 49932
rect 31067 49929 31079 49963
rect 31021 49923 31079 49929
rect 31481 49963 31539 49969
rect 31481 49929 31493 49963
rect 31527 49960 31539 49963
rect 31662 49960 31668 49972
rect 31527 49932 31668 49960
rect 31527 49929 31539 49932
rect 31481 49923 31539 49929
rect 31662 49920 31668 49932
rect 31720 49920 31726 49972
rect 32582 49920 32588 49972
rect 32640 49960 32646 49972
rect 32677 49963 32735 49969
rect 32677 49960 32689 49963
rect 32640 49932 32689 49960
rect 32640 49920 32646 49932
rect 32677 49929 32689 49932
rect 32723 49960 32735 49963
rect 32766 49960 32772 49972
rect 32723 49932 32772 49960
rect 32723 49929 32735 49932
rect 32677 49923 32735 49929
rect 32766 49920 32772 49932
rect 32824 49920 32830 49972
rect 32858 49920 32864 49972
rect 32916 49960 32922 49972
rect 33505 49963 33563 49969
rect 33505 49960 33517 49963
rect 32916 49932 33517 49960
rect 32916 49920 32922 49932
rect 33505 49929 33517 49932
rect 33551 49929 33563 49963
rect 33505 49923 33563 49929
rect 33965 49963 34023 49969
rect 33965 49929 33977 49963
rect 34011 49960 34023 49963
rect 34514 49960 34520 49972
rect 34011 49932 34520 49960
rect 34011 49929 34023 49932
rect 33965 49923 34023 49929
rect 34514 49920 34520 49932
rect 34572 49920 34578 49972
rect 34701 49963 34759 49969
rect 34701 49929 34713 49963
rect 34747 49929 34759 49963
rect 34701 49923 34759 49929
rect 30193 49895 30251 49901
rect 30193 49861 30205 49895
rect 30239 49892 30251 49895
rect 30466 49892 30472 49904
rect 30239 49864 30472 49892
rect 30239 49861 30251 49864
rect 30193 49855 30251 49861
rect 30466 49852 30472 49864
rect 30524 49892 30530 49904
rect 30742 49892 30748 49904
rect 30524 49864 30748 49892
rect 30524 49852 30530 49864
rect 30742 49852 30748 49864
rect 30800 49852 30806 49904
rect 31389 49895 31447 49901
rect 31389 49861 31401 49895
rect 31435 49892 31447 49895
rect 33594 49892 33600 49904
rect 31435 49864 33600 49892
rect 31435 49861 31447 49864
rect 31389 49855 31447 49861
rect 33594 49852 33600 49864
rect 33652 49892 33658 49904
rect 33873 49895 33931 49901
rect 33873 49892 33885 49895
rect 33652 49864 33885 49892
rect 33652 49852 33658 49864
rect 33873 49861 33885 49864
rect 33919 49861 33931 49895
rect 34716 49892 34744 49923
rect 35158 49920 35164 49972
rect 35216 49960 35222 49972
rect 39022 49960 39028 49972
rect 35216 49932 39028 49960
rect 35216 49920 35222 49932
rect 39022 49920 39028 49932
rect 39080 49920 39086 49972
rect 36998 49892 37004 49904
rect 34716 49864 37004 49892
rect 33873 49855 33931 49861
rect 36998 49852 37004 49864
rect 37056 49852 37062 49904
rect 30285 49827 30343 49833
rect 30285 49793 30297 49827
rect 30331 49824 30343 49827
rect 31938 49824 31944 49836
rect 30331 49796 31944 49824
rect 30331 49793 30343 49796
rect 30285 49787 30343 49793
rect 31938 49784 31944 49796
rect 31996 49824 32002 49836
rect 32582 49824 32588 49836
rect 31996 49796 32588 49824
rect 31996 49784 32002 49796
rect 32582 49784 32588 49796
rect 32640 49784 32646 49836
rect 32674 49784 32680 49836
rect 32732 49824 32738 49836
rect 32732 49796 32904 49824
rect 32732 49784 32738 49796
rect 27724 49728 29960 49756
rect 16666 49688 16672 49700
rect 14936 49660 16672 49688
rect 16666 49648 16672 49660
rect 16724 49648 16730 49700
rect 27338 49648 27344 49700
rect 27396 49688 27402 49700
rect 27724 49688 27752 49728
rect 30190 49716 30196 49768
rect 30248 49756 30254 49768
rect 30377 49759 30435 49765
rect 30377 49756 30389 49759
rect 30248 49728 30389 49756
rect 30248 49716 30254 49728
rect 30377 49725 30389 49728
rect 30423 49725 30435 49759
rect 30377 49719 30435 49725
rect 31570 49716 31576 49768
rect 31628 49716 31634 49768
rect 31662 49716 31668 49768
rect 31720 49756 31726 49768
rect 32876 49765 32904 49796
rect 32950 49784 32956 49836
rect 33008 49824 33014 49836
rect 35069 49827 35127 49833
rect 35069 49824 35081 49827
rect 33008 49796 35081 49824
rect 33008 49784 33014 49796
rect 35069 49793 35081 49796
rect 35115 49793 35127 49827
rect 37090 49824 37096 49836
rect 35069 49787 35127 49793
rect 35268 49796 37096 49824
rect 32769 49759 32827 49765
rect 31720 49728 32352 49756
rect 31720 49716 31726 49728
rect 32324 49697 32352 49728
rect 32769 49725 32781 49759
rect 32815 49725 32827 49759
rect 32769 49719 32827 49725
rect 32861 49759 32919 49765
rect 32861 49725 32873 49759
rect 32907 49725 32919 49759
rect 34054 49756 34060 49768
rect 32861 49719 32919 49725
rect 32968 49728 34060 49756
rect 27396 49660 27752 49688
rect 32309 49691 32367 49697
rect 27396 49648 27402 49660
rect 32309 49657 32321 49691
rect 32355 49657 32367 49691
rect 32784 49688 32812 49719
rect 32968 49688 32996 49728
rect 34054 49716 34060 49728
rect 34112 49716 34118 49768
rect 34149 49759 34207 49765
rect 34149 49725 34161 49759
rect 34195 49725 34207 49759
rect 34149 49719 34207 49725
rect 32784 49660 32996 49688
rect 32309 49651 32367 49657
rect 15194 49620 15200 49632
rect 14844 49592 15200 49620
rect 15194 49580 15200 49592
rect 15252 49580 15258 49632
rect 27154 49580 27160 49632
rect 27212 49620 27218 49632
rect 27880 49623 27938 49629
rect 27880 49620 27892 49623
rect 27212 49592 27892 49620
rect 27212 49580 27218 49592
rect 27880 49589 27892 49592
rect 27926 49620 27938 49623
rect 29086 49620 29092 49632
rect 27926 49592 29092 49620
rect 27926 49589 27938 49592
rect 27880 49583 27938 49589
rect 29086 49580 29092 49592
rect 29144 49580 29150 49632
rect 29362 49580 29368 49632
rect 29420 49580 29426 49632
rect 32490 49580 32496 49632
rect 32548 49620 32554 49632
rect 34164 49620 34192 49719
rect 34238 49716 34244 49768
rect 34296 49756 34302 49768
rect 35268 49756 35296 49796
rect 37090 49784 37096 49796
rect 37148 49784 37154 49836
rect 49326 49784 49332 49836
rect 49384 49784 49390 49836
rect 34296 49728 35296 49756
rect 35345 49759 35403 49765
rect 34296 49716 34302 49728
rect 35345 49725 35357 49759
rect 35391 49756 35403 49759
rect 36630 49756 36636 49768
rect 35391 49728 36636 49756
rect 35391 49725 35403 49728
rect 35345 49719 35403 49725
rect 36630 49716 36636 49728
rect 36688 49716 36694 49768
rect 43438 49716 43444 49768
rect 43496 49756 43502 49768
rect 43496 49728 49188 49756
rect 43496 49716 43502 49728
rect 49160 49697 49188 49728
rect 49145 49691 49203 49697
rect 49145 49657 49157 49691
rect 49191 49657 49203 49691
rect 49145 49651 49203 49657
rect 32548 49592 34192 49620
rect 32548 49580 32554 49592
rect 1104 49530 49864 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 32950 49530
rect 33002 49478 33014 49530
rect 33066 49478 33078 49530
rect 33130 49478 33142 49530
rect 33194 49478 33206 49530
rect 33258 49478 42950 49530
rect 43002 49478 43014 49530
rect 43066 49478 43078 49530
rect 43130 49478 43142 49530
rect 43194 49478 43206 49530
rect 43258 49478 49864 49530
rect 1104 49456 49864 49478
rect 8478 49376 8484 49428
rect 8536 49416 8542 49428
rect 10045 49419 10103 49425
rect 10045 49416 10057 49419
rect 8536 49388 10057 49416
rect 8536 49376 8542 49388
rect 10045 49385 10057 49388
rect 10091 49385 10103 49419
rect 13449 49419 13507 49425
rect 13449 49416 13461 49419
rect 10045 49379 10103 49385
rect 12406 49388 13461 49416
rect 9766 49308 9772 49360
rect 9824 49348 9830 49360
rect 12406 49348 12434 49388
rect 13449 49385 13461 49388
rect 13495 49385 13507 49419
rect 13449 49379 13507 49385
rect 15286 49376 15292 49428
rect 15344 49416 15350 49428
rect 19981 49419 20039 49425
rect 19981 49416 19993 49419
rect 15344 49388 19993 49416
rect 15344 49376 15350 49388
rect 19981 49385 19993 49388
rect 20027 49385 20039 49419
rect 19981 49379 20039 49385
rect 24946 49376 24952 49428
rect 25004 49416 25010 49428
rect 28813 49419 28871 49425
rect 28813 49416 28825 49419
rect 25004 49388 28825 49416
rect 25004 49376 25010 49388
rect 28813 49385 28825 49388
rect 28859 49385 28871 49419
rect 28813 49379 28871 49385
rect 30098 49376 30104 49428
rect 30156 49416 30162 49428
rect 30156 49388 33456 49416
rect 30156 49376 30162 49388
rect 9824 49320 12434 49348
rect 9824 49308 9830 49320
rect 27154 49308 27160 49360
rect 27212 49308 27218 49360
rect 29454 49348 29460 49360
rect 28092 49320 29460 49348
rect 1302 49240 1308 49292
rect 1360 49280 1366 49292
rect 28092 49289 28120 49320
rect 29454 49308 29460 49320
rect 29512 49308 29518 49360
rect 33318 49348 33324 49360
rect 33060 49320 33324 49348
rect 2041 49283 2099 49289
rect 2041 49280 2053 49283
rect 1360 49252 2053 49280
rect 1360 49240 1366 49252
rect 2041 49249 2053 49252
rect 2087 49249 2099 49283
rect 2041 49243 2099 49249
rect 28077 49283 28135 49289
rect 28077 49249 28089 49283
rect 28123 49249 28135 49283
rect 28077 49243 28135 49249
rect 28169 49283 28227 49289
rect 28169 49249 28181 49283
rect 28215 49249 28227 49283
rect 28169 49243 28227 49249
rect 1765 49215 1823 49221
rect 1765 49181 1777 49215
rect 1811 49212 1823 49215
rect 5810 49212 5816 49224
rect 1811 49184 5816 49212
rect 1811 49181 1823 49184
rect 1765 49175 1823 49181
rect 5810 49172 5816 49184
rect 5868 49172 5874 49224
rect 25406 49172 25412 49224
rect 25464 49172 25470 49224
rect 26786 49172 26792 49224
rect 26844 49172 26850 49224
rect 26970 49172 26976 49224
rect 27028 49212 27034 49224
rect 28184 49212 28212 49243
rect 29362 49240 29368 49292
rect 29420 49280 29426 49292
rect 30285 49283 30343 49289
rect 30285 49280 30297 49283
rect 29420 49252 30297 49280
rect 29420 49240 29426 49252
rect 30285 49249 30297 49252
rect 30331 49249 30343 49283
rect 33060 49280 33088 49320
rect 33318 49308 33324 49320
rect 33376 49308 33382 49360
rect 33428 49348 33456 49388
rect 33502 49376 33508 49428
rect 33560 49376 33566 49428
rect 34422 49376 34428 49428
rect 34480 49416 34486 49428
rect 34885 49419 34943 49425
rect 34885 49416 34897 49419
rect 34480 49388 34897 49416
rect 34480 49376 34486 49388
rect 34885 49385 34897 49388
rect 34931 49385 34943 49419
rect 34885 49379 34943 49385
rect 36538 49348 36544 49360
rect 33428 49320 36544 49348
rect 36538 49308 36544 49320
rect 36596 49308 36602 49360
rect 30285 49243 30343 49249
rect 30392 49252 33088 49280
rect 27028 49184 28212 49212
rect 28997 49215 29055 49221
rect 27028 49172 27034 49184
rect 28997 49181 29009 49215
rect 29043 49212 29055 49215
rect 30392 49212 30420 49252
rect 34146 49240 34152 49292
rect 34204 49280 34210 49292
rect 35437 49283 35495 49289
rect 35437 49280 35449 49283
rect 34204 49252 35449 49280
rect 34204 49240 34210 49252
rect 35437 49249 35449 49252
rect 35483 49249 35495 49283
rect 35437 49243 35495 49249
rect 29043 49184 30420 49212
rect 29043 49181 29055 49184
rect 28997 49175 29055 49181
rect 31754 49172 31760 49224
rect 31812 49172 31818 49224
rect 33318 49172 33324 49224
rect 33376 49212 33382 49224
rect 33594 49212 33600 49224
rect 33376 49184 33600 49212
rect 33376 49172 33382 49184
rect 33594 49172 33600 49184
rect 33652 49172 33658 49224
rect 34698 49172 34704 49224
rect 34756 49212 34762 49224
rect 34756 49184 41414 49212
rect 34756 49172 34762 49184
rect 9953 49147 10011 49153
rect 9953 49113 9965 49147
rect 9999 49144 10011 49147
rect 11974 49144 11980 49156
rect 9999 49116 11980 49144
rect 9999 49113 10011 49116
rect 9953 49107 10011 49113
rect 11974 49104 11980 49116
rect 12032 49104 12038 49156
rect 13357 49147 13415 49153
rect 13357 49113 13369 49147
rect 13403 49144 13415 49147
rect 16390 49144 16396 49156
rect 13403 49116 16396 49144
rect 13403 49113 13415 49116
rect 13357 49107 13415 49113
rect 16390 49104 16396 49116
rect 16448 49104 16454 49156
rect 19889 49147 19947 49153
rect 19889 49113 19901 49147
rect 19935 49144 19947 49147
rect 22738 49144 22744 49156
rect 19935 49116 22744 49144
rect 19935 49113 19947 49116
rect 19889 49107 19947 49113
rect 22738 49104 22744 49116
rect 22796 49104 22802 49156
rect 25682 49104 25688 49156
rect 25740 49104 25746 49156
rect 27985 49147 28043 49153
rect 27985 49113 27997 49147
rect 28031 49144 28043 49147
rect 29178 49144 29184 49156
rect 28031 49116 29184 49144
rect 28031 49113 28043 49116
rect 27985 49107 28043 49113
rect 29178 49104 29184 49116
rect 29236 49104 29242 49156
rect 30098 49104 30104 49156
rect 30156 49104 30162 49156
rect 30193 49147 30251 49153
rect 30193 49113 30205 49147
rect 30239 49144 30251 49147
rect 31018 49144 31024 49156
rect 30239 49116 31024 49144
rect 30239 49113 30251 49116
rect 30193 49107 30251 49113
rect 31018 49104 31024 49116
rect 31076 49104 31082 49156
rect 32030 49104 32036 49156
rect 32088 49104 32094 49156
rect 33778 49144 33784 49156
rect 33258 49116 33784 49144
rect 33778 49104 33784 49116
rect 33836 49104 33842 49156
rect 35253 49147 35311 49153
rect 35253 49113 35265 49147
rect 35299 49144 35311 49147
rect 37182 49144 37188 49156
rect 35299 49116 37188 49144
rect 35299 49113 35311 49116
rect 35253 49107 35311 49113
rect 37182 49104 37188 49116
rect 37240 49104 37246 49156
rect 41386 49144 41414 49184
rect 49050 49172 49056 49224
rect 49108 49172 49114 49224
rect 41386 49116 45554 49144
rect 27246 49036 27252 49088
rect 27304 49076 27310 49088
rect 27617 49079 27675 49085
rect 27617 49076 27629 49079
rect 27304 49048 27629 49076
rect 27304 49036 27310 49048
rect 27617 49045 27629 49048
rect 27663 49045 27675 49079
rect 27617 49039 27675 49045
rect 28994 49036 29000 49088
rect 29052 49076 29058 49088
rect 29733 49079 29791 49085
rect 29733 49076 29745 49079
rect 29052 49048 29745 49076
rect 29052 49036 29058 49048
rect 29733 49045 29745 49048
rect 29779 49045 29791 49079
rect 29733 49039 29791 49045
rect 30374 49036 30380 49088
rect 30432 49076 30438 49088
rect 33410 49076 33416 49088
rect 30432 49048 33416 49076
rect 30432 49036 30438 49048
rect 33410 49036 33416 49048
rect 33468 49036 33474 49088
rect 35342 49036 35348 49088
rect 35400 49036 35406 49088
rect 45526 49076 45554 49116
rect 49237 49079 49295 49085
rect 49237 49076 49249 49079
rect 45526 49048 49249 49076
rect 49237 49045 49249 49048
rect 49283 49045 49295 49079
rect 49237 49039 49295 49045
rect 1104 48986 49864 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 27950 48986
rect 28002 48934 28014 48986
rect 28066 48934 28078 48986
rect 28130 48934 28142 48986
rect 28194 48934 28206 48986
rect 28258 48934 37950 48986
rect 38002 48934 38014 48986
rect 38066 48934 38078 48986
rect 38130 48934 38142 48986
rect 38194 48934 38206 48986
rect 38258 48934 47950 48986
rect 48002 48934 48014 48986
rect 48066 48934 48078 48986
rect 48130 48934 48142 48986
rect 48194 48934 48206 48986
rect 48258 48934 49864 48986
rect 1104 48912 49864 48934
rect 24762 48832 24768 48884
rect 24820 48872 24826 48884
rect 25225 48875 25283 48881
rect 25225 48872 25237 48875
rect 24820 48844 25237 48872
rect 24820 48832 24826 48844
rect 25225 48841 25237 48844
rect 25271 48841 25283 48875
rect 25225 48835 25283 48841
rect 26329 48875 26387 48881
rect 26329 48841 26341 48875
rect 26375 48872 26387 48875
rect 27617 48875 27675 48881
rect 26375 48844 27568 48872
rect 26375 48841 26387 48844
rect 26329 48835 26387 48841
rect 24213 48807 24271 48813
rect 24213 48773 24225 48807
rect 24259 48804 24271 48807
rect 27246 48804 27252 48816
rect 24259 48776 27252 48804
rect 24259 48773 24271 48776
rect 24213 48767 24271 48773
rect 27246 48764 27252 48776
rect 27304 48764 27310 48816
rect 27540 48804 27568 48844
rect 27617 48841 27629 48875
rect 27663 48872 27675 48875
rect 30837 48875 30895 48881
rect 30837 48872 30849 48875
rect 27663 48844 30849 48872
rect 27663 48841 27675 48844
rect 27617 48835 27675 48841
rect 30837 48841 30849 48844
rect 30883 48872 30895 48875
rect 31846 48872 31852 48884
rect 30883 48844 31852 48872
rect 30883 48841 30895 48844
rect 30837 48835 30895 48841
rect 31846 48832 31852 48844
rect 31904 48832 31910 48884
rect 32030 48832 32036 48884
rect 32088 48872 32094 48884
rect 33042 48872 33048 48884
rect 32088 48844 33048 48872
rect 32088 48832 32094 48844
rect 33042 48832 33048 48844
rect 33100 48832 33106 48884
rect 33410 48832 33416 48884
rect 33468 48872 33474 48884
rect 34977 48875 35035 48881
rect 34977 48872 34989 48875
rect 33468 48844 34989 48872
rect 33468 48832 33474 48844
rect 34977 48841 34989 48844
rect 35023 48841 35035 48875
rect 34977 48835 35035 48841
rect 35069 48875 35127 48881
rect 35069 48841 35081 48875
rect 35115 48872 35127 48875
rect 35250 48872 35256 48884
rect 35115 48844 35256 48872
rect 35115 48841 35127 48844
rect 35069 48835 35127 48841
rect 35250 48832 35256 48844
rect 35308 48832 35314 48884
rect 29270 48804 29276 48816
rect 27540 48776 29276 48804
rect 29270 48764 29276 48776
rect 29328 48764 29334 48816
rect 29641 48807 29699 48813
rect 29641 48773 29653 48807
rect 29687 48804 29699 48807
rect 32677 48807 32735 48813
rect 32677 48804 32689 48807
rect 29687 48776 31754 48804
rect 29687 48773 29699 48776
rect 29641 48767 29699 48773
rect 24121 48739 24179 48745
rect 24121 48705 24133 48739
rect 24167 48736 24179 48739
rect 25038 48736 25044 48748
rect 24167 48708 25044 48736
rect 24167 48705 24179 48708
rect 24121 48699 24179 48705
rect 25038 48696 25044 48708
rect 25096 48696 25102 48748
rect 25409 48739 25467 48745
rect 25409 48705 25421 48739
rect 25455 48705 25467 48739
rect 25409 48699 25467 48705
rect 26237 48739 26295 48745
rect 26237 48705 26249 48739
rect 26283 48705 26295 48739
rect 26237 48699 26295 48705
rect 23474 48628 23480 48680
rect 23532 48668 23538 48680
rect 24305 48671 24363 48677
rect 24305 48668 24317 48671
rect 23532 48640 24317 48668
rect 23532 48628 23538 48640
rect 24305 48637 24317 48640
rect 24351 48637 24363 48671
rect 25424 48668 25452 48699
rect 25424 48640 26188 48668
rect 24305 48631 24363 48637
rect 20990 48560 20996 48612
rect 21048 48600 21054 48612
rect 25869 48603 25927 48609
rect 25869 48600 25881 48603
rect 21048 48572 25881 48600
rect 21048 48560 21054 48572
rect 25869 48569 25881 48572
rect 25915 48569 25927 48603
rect 25869 48563 25927 48569
rect 18874 48492 18880 48544
rect 18932 48532 18938 48544
rect 23753 48535 23811 48541
rect 23753 48532 23765 48535
rect 18932 48504 23765 48532
rect 18932 48492 18938 48504
rect 23753 48501 23765 48504
rect 23799 48501 23811 48535
rect 26160 48532 26188 48640
rect 26252 48600 26280 48699
rect 27430 48696 27436 48748
rect 27488 48736 27494 48748
rect 27525 48739 27583 48745
rect 27525 48736 27537 48739
rect 27488 48708 27537 48736
rect 27488 48696 27494 48708
rect 27525 48705 27537 48708
rect 27571 48736 27583 48739
rect 27571 48708 28580 48736
rect 27571 48705 27583 48708
rect 27525 48699 27583 48705
rect 26418 48628 26424 48680
rect 26476 48628 26482 48680
rect 26510 48628 26516 48680
rect 26568 48668 26574 48680
rect 27709 48671 27767 48677
rect 27709 48668 27721 48671
rect 26568 48640 27721 48668
rect 26568 48628 26574 48640
rect 27709 48637 27721 48640
rect 27755 48637 27767 48671
rect 28552 48668 28580 48708
rect 29546 48696 29552 48748
rect 29604 48696 29610 48748
rect 30745 48739 30803 48745
rect 30745 48736 30757 48739
rect 29656 48708 30757 48736
rect 29656 48668 29684 48708
rect 30745 48705 30757 48708
rect 30791 48705 30803 48739
rect 30745 48699 30803 48705
rect 28552 48640 29684 48668
rect 29825 48671 29883 48677
rect 27709 48631 27767 48637
rect 29825 48637 29837 48671
rect 29871 48668 29883 48671
rect 30650 48668 30656 48680
rect 29871 48640 30656 48668
rect 29871 48637 29883 48640
rect 29825 48631 29883 48637
rect 30650 48628 30656 48640
rect 30708 48628 30714 48680
rect 31021 48671 31079 48677
rect 31021 48637 31033 48671
rect 31067 48668 31079 48671
rect 31202 48668 31208 48680
rect 31067 48640 31208 48668
rect 31067 48637 31079 48640
rect 31021 48631 31079 48637
rect 31202 48628 31208 48640
rect 31260 48628 31266 48680
rect 31726 48668 31754 48776
rect 31864 48776 32689 48804
rect 31864 48748 31892 48776
rect 32677 48773 32689 48776
rect 32723 48773 32735 48807
rect 32677 48767 32735 48773
rect 31846 48696 31852 48748
rect 31904 48696 31910 48748
rect 33778 48696 33784 48748
rect 33836 48696 33842 48748
rect 32306 48668 32312 48680
rect 31726 48640 32312 48668
rect 32306 48628 32312 48640
rect 32364 48628 32370 48680
rect 32401 48671 32459 48677
rect 32401 48637 32413 48671
rect 32447 48637 32459 48671
rect 32401 48631 32459 48637
rect 28534 48600 28540 48612
rect 26252 48572 28540 48600
rect 28534 48560 28540 48572
rect 28592 48560 28598 48612
rect 28902 48560 28908 48612
rect 28960 48600 28966 48612
rect 29181 48603 29239 48609
rect 29181 48600 29193 48603
rect 28960 48572 29193 48600
rect 28960 48560 28966 48572
rect 29181 48569 29193 48572
rect 29227 48569 29239 48603
rect 29181 48563 29239 48569
rect 29270 48560 29276 48612
rect 29328 48600 29334 48612
rect 30282 48600 30288 48612
rect 29328 48572 30288 48600
rect 29328 48560 29334 48572
rect 30282 48560 30288 48572
rect 30340 48560 30346 48612
rect 27062 48532 27068 48544
rect 26160 48504 27068 48532
rect 23753 48495 23811 48501
rect 27062 48492 27068 48504
rect 27120 48492 27126 48544
rect 27154 48492 27160 48544
rect 27212 48492 27218 48544
rect 30377 48535 30435 48541
rect 30377 48501 30389 48535
rect 30423 48532 30435 48535
rect 30742 48532 30748 48544
rect 30423 48504 30748 48532
rect 30423 48501 30435 48504
rect 30377 48495 30435 48501
rect 30742 48492 30748 48504
rect 30800 48492 30806 48544
rect 32416 48532 32444 48631
rect 33042 48628 33048 48680
rect 33100 48668 33106 48680
rect 34146 48668 34152 48680
rect 33100 48640 34152 48668
rect 33100 48628 33106 48640
rect 34146 48628 34152 48640
rect 34204 48628 34210 48680
rect 34330 48628 34336 48680
rect 34388 48668 34394 48680
rect 35161 48671 35219 48677
rect 35161 48668 35173 48671
rect 34388 48640 35173 48668
rect 34388 48628 34394 48640
rect 35161 48637 35173 48640
rect 35207 48637 35219 48671
rect 35161 48631 35219 48637
rect 34514 48600 34520 48612
rect 33693 48572 34520 48600
rect 33693 48532 33721 48572
rect 34514 48560 34520 48572
rect 34572 48560 34578 48612
rect 32416 48504 33721 48532
rect 33962 48492 33968 48544
rect 34020 48532 34026 48544
rect 34609 48535 34667 48541
rect 34609 48532 34621 48535
rect 34020 48504 34621 48532
rect 34020 48492 34026 48504
rect 34609 48501 34621 48504
rect 34655 48501 34667 48535
rect 34609 48495 34667 48501
rect 1104 48442 49864 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 32950 48442
rect 33002 48390 33014 48442
rect 33066 48390 33078 48442
rect 33130 48390 33142 48442
rect 33194 48390 33206 48442
rect 33258 48390 42950 48442
rect 43002 48390 43014 48442
rect 43066 48390 43078 48442
rect 43130 48390 43142 48442
rect 43194 48390 43206 48442
rect 43258 48390 49864 48442
rect 1104 48368 49864 48390
rect 25222 48288 25228 48340
rect 25280 48328 25286 48340
rect 27154 48328 27160 48340
rect 25280 48300 27160 48328
rect 25280 48288 25286 48300
rect 27154 48288 27160 48300
rect 27212 48288 27218 48340
rect 27706 48288 27712 48340
rect 27764 48328 27770 48340
rect 27764 48300 28396 48328
rect 27764 48288 27770 48300
rect 28368 48260 28396 48300
rect 32306 48288 32312 48340
rect 32364 48328 32370 48340
rect 34790 48328 34796 48340
rect 32364 48300 34796 48328
rect 32364 48288 32370 48300
rect 34790 48288 34796 48300
rect 34848 48288 34854 48340
rect 34885 48331 34943 48337
rect 34885 48297 34897 48331
rect 34931 48328 34943 48331
rect 35342 48328 35348 48340
rect 34931 48300 35348 48328
rect 34931 48297 34943 48300
rect 34885 48291 34943 48297
rect 35342 48288 35348 48300
rect 35400 48288 35406 48340
rect 28626 48260 28632 48272
rect 28368 48232 28632 48260
rect 28626 48220 28632 48232
rect 28684 48220 28690 48272
rect 33045 48263 33103 48269
rect 33045 48229 33057 48263
rect 33091 48229 33103 48263
rect 37366 48260 37372 48272
rect 33045 48223 33103 48229
rect 33520 48232 37372 48260
rect 1302 48152 1308 48204
rect 1360 48192 1366 48204
rect 2041 48195 2099 48201
rect 2041 48192 2053 48195
rect 1360 48164 2053 48192
rect 1360 48152 1366 48164
rect 2041 48161 2053 48164
rect 2087 48161 2099 48195
rect 2041 48155 2099 48161
rect 20349 48195 20407 48201
rect 20349 48161 20361 48195
rect 20395 48192 20407 48195
rect 21450 48192 21456 48204
rect 20395 48164 21456 48192
rect 20395 48161 20407 48164
rect 20349 48155 20407 48161
rect 21450 48152 21456 48164
rect 21508 48152 21514 48204
rect 25406 48152 25412 48204
rect 25464 48192 25470 48204
rect 26050 48192 26056 48204
rect 25464 48164 26056 48192
rect 25464 48152 25470 48164
rect 26050 48152 26056 48164
rect 26108 48192 26114 48204
rect 27065 48195 27123 48201
rect 27065 48192 27077 48195
rect 26108 48164 27077 48192
rect 26108 48152 26114 48164
rect 27065 48161 27077 48164
rect 27111 48192 27123 48195
rect 27706 48192 27712 48204
rect 27111 48164 27712 48192
rect 27111 48161 27123 48164
rect 27065 48155 27123 48161
rect 27706 48152 27712 48164
rect 27764 48152 27770 48204
rect 28350 48152 28356 48204
rect 28408 48192 28414 48204
rect 28718 48192 28724 48204
rect 28408 48164 28724 48192
rect 28408 48152 28414 48164
rect 28718 48152 28724 48164
rect 28776 48152 28782 48204
rect 30650 48152 30656 48204
rect 30708 48192 30714 48204
rect 31018 48192 31024 48204
rect 30708 48164 31024 48192
rect 30708 48152 30714 48164
rect 31018 48152 31024 48164
rect 31076 48152 31082 48204
rect 31386 48152 31392 48204
rect 31444 48192 31450 48204
rect 33060 48192 33088 48223
rect 33520 48201 33548 48232
rect 37366 48220 37372 48232
rect 37424 48220 37430 48272
rect 31444 48164 33088 48192
rect 33505 48195 33563 48201
rect 31444 48152 31450 48164
rect 33505 48161 33517 48195
rect 33551 48161 33563 48195
rect 33505 48155 33563 48161
rect 33689 48195 33747 48201
rect 33689 48161 33701 48195
rect 33735 48192 33747 48195
rect 35342 48192 35348 48204
rect 33735 48164 35348 48192
rect 33735 48161 33747 48164
rect 33689 48155 33747 48161
rect 35342 48152 35348 48164
rect 35400 48152 35406 48204
rect 35437 48195 35495 48201
rect 35437 48161 35449 48195
rect 35483 48161 35495 48195
rect 35437 48155 35495 48161
rect 1765 48127 1823 48133
rect 1765 48093 1777 48127
rect 1811 48124 1823 48127
rect 11054 48124 11060 48136
rect 1811 48096 11060 48124
rect 1811 48093 1823 48096
rect 1765 48087 1823 48093
rect 11054 48084 11060 48096
rect 11112 48084 11118 48136
rect 18506 48084 18512 48136
rect 18564 48124 18570 48136
rect 21729 48127 21787 48133
rect 21729 48124 21741 48127
rect 18564 48096 21741 48124
rect 18564 48084 18570 48096
rect 21729 48093 21741 48096
rect 21775 48093 21787 48127
rect 21729 48087 21787 48093
rect 22094 48084 22100 48136
rect 22152 48124 22158 48136
rect 22281 48127 22339 48133
rect 22281 48124 22293 48127
rect 22152 48096 22293 48124
rect 22152 48084 22158 48096
rect 22281 48093 22293 48096
rect 22327 48093 22339 48127
rect 22281 48087 22339 48093
rect 24670 48084 24676 48136
rect 24728 48124 24734 48136
rect 24765 48127 24823 48133
rect 24765 48124 24777 48127
rect 24728 48096 24777 48124
rect 24728 48084 24734 48096
rect 24765 48093 24777 48096
rect 24811 48093 24823 48127
rect 24765 48087 24823 48093
rect 30006 48084 30012 48136
rect 30064 48124 30070 48136
rect 30745 48127 30803 48133
rect 30745 48124 30757 48127
rect 30064 48096 30757 48124
rect 30064 48084 30070 48096
rect 30745 48093 30757 48096
rect 30791 48093 30803 48127
rect 30745 48087 30803 48093
rect 32122 48084 32128 48136
rect 32180 48084 32186 48136
rect 35452 48124 35480 48155
rect 36814 48152 36820 48204
rect 36872 48201 36878 48204
rect 36872 48195 36921 48201
rect 36872 48161 36875 48195
rect 36909 48161 36921 48195
rect 36872 48155 36921 48161
rect 36872 48152 36878 48155
rect 35452 48096 36860 48124
rect 22554 48016 22560 48068
rect 22612 48016 22618 48068
rect 24578 48056 24584 48068
rect 23782 48028 24584 48056
rect 24578 48016 24584 48028
rect 24636 48016 24642 48068
rect 25041 48059 25099 48065
rect 25041 48025 25053 48059
rect 25087 48056 25099 48059
rect 25130 48056 25136 48068
rect 25087 48028 25136 48056
rect 25087 48025 25099 48028
rect 25041 48019 25099 48025
rect 25130 48016 25136 48028
rect 25188 48016 25194 48068
rect 25498 48016 25504 48068
rect 25556 48016 25562 48068
rect 27341 48059 27399 48065
rect 27341 48025 27353 48059
rect 27387 48056 27399 48059
rect 27430 48056 27436 48068
rect 27387 48028 27436 48056
rect 27387 48025 27399 48028
rect 27341 48019 27399 48025
rect 27430 48016 27436 48028
rect 27488 48016 27494 48068
rect 29086 48056 29092 48068
rect 28566 48028 29092 48056
rect 29086 48016 29092 48028
rect 29144 48056 29150 48068
rect 31294 48056 31300 48068
rect 29144 48028 31300 48056
rect 29144 48016 29150 48028
rect 31294 48016 31300 48028
rect 31352 48016 31358 48068
rect 32674 48056 32680 48068
rect 32324 48028 32680 48056
rect 16574 47948 16580 48000
rect 16632 47988 16638 48000
rect 19705 47991 19763 47997
rect 19705 47988 19717 47991
rect 16632 47960 19717 47988
rect 16632 47948 16638 47960
rect 19705 47957 19717 47960
rect 19751 47957 19763 47991
rect 19705 47951 19763 47957
rect 19794 47948 19800 48000
rect 19852 47988 19858 48000
rect 20073 47991 20131 47997
rect 20073 47988 20085 47991
rect 19852 47960 20085 47988
rect 19852 47948 19858 47960
rect 20073 47957 20085 47960
rect 20119 47957 20131 47991
rect 20073 47951 20131 47957
rect 20165 47991 20223 47997
rect 20165 47957 20177 47991
rect 20211 47988 20223 47991
rect 22002 47988 22008 48000
rect 20211 47960 22008 47988
rect 20211 47957 20223 47960
rect 20165 47951 20223 47957
rect 22002 47948 22008 47960
rect 22060 47948 22066 48000
rect 22646 47948 22652 48000
rect 22704 47988 22710 48000
rect 24029 47991 24087 47997
rect 24029 47988 24041 47991
rect 22704 47960 24041 47988
rect 22704 47948 22710 47960
rect 24029 47957 24041 47960
rect 24075 47957 24087 47991
rect 24029 47951 24087 47957
rect 24762 47948 24768 48000
rect 24820 47988 24826 48000
rect 26513 47991 26571 47997
rect 26513 47988 26525 47991
rect 24820 47960 26525 47988
rect 24820 47948 24826 47960
rect 26513 47957 26525 47960
rect 26559 47988 26571 47991
rect 27246 47988 27252 48000
rect 26559 47960 27252 47988
rect 26559 47957 26571 47960
rect 26513 47951 26571 47957
rect 27246 47948 27252 47960
rect 27304 47948 27310 48000
rect 27706 47948 27712 48000
rect 27764 47988 27770 48000
rect 28813 47991 28871 47997
rect 28813 47988 28825 47991
rect 27764 47960 28825 47988
rect 27764 47948 27770 47960
rect 28813 47957 28825 47960
rect 28859 47988 28871 47991
rect 32324 47988 32352 48028
rect 32674 48016 32680 48028
rect 32732 48016 32738 48068
rect 35452 48056 35480 48096
rect 32784 48028 35480 48056
rect 32784 48000 32812 48028
rect 36354 48016 36360 48068
rect 36412 48056 36418 48068
rect 36633 48059 36691 48065
rect 36633 48056 36645 48059
rect 36412 48028 36645 48056
rect 36412 48016 36418 48028
rect 36633 48025 36645 48028
rect 36679 48025 36691 48059
rect 36633 48019 36691 48025
rect 36722 48016 36728 48068
rect 36780 48016 36786 48068
rect 28859 47960 32352 47988
rect 32493 47991 32551 47997
rect 28859 47957 28871 47960
rect 28813 47951 28871 47957
rect 32493 47957 32505 47991
rect 32539 47988 32551 47991
rect 32766 47988 32772 48000
rect 32539 47960 32772 47988
rect 32539 47957 32551 47960
rect 32493 47951 32551 47957
rect 32766 47948 32772 47960
rect 32824 47948 32830 48000
rect 33410 47948 33416 48000
rect 33468 47948 33474 48000
rect 34974 47948 34980 48000
rect 35032 47988 35038 48000
rect 35253 47991 35311 47997
rect 35253 47988 35265 47991
rect 35032 47960 35265 47988
rect 35032 47948 35038 47960
rect 35253 47957 35265 47960
rect 35299 47957 35311 47991
rect 35253 47951 35311 47957
rect 35345 47991 35403 47997
rect 35345 47957 35357 47991
rect 35391 47988 35403 47991
rect 35434 47988 35440 48000
rect 35391 47960 35440 47988
rect 35391 47957 35403 47960
rect 35345 47951 35403 47957
rect 35434 47948 35440 47960
rect 35492 47948 35498 48000
rect 35710 47948 35716 48000
rect 35768 47988 35774 48000
rect 36081 47991 36139 47997
rect 36081 47988 36093 47991
rect 35768 47960 36093 47988
rect 35768 47948 35774 47960
rect 36081 47957 36093 47960
rect 36127 47957 36139 47991
rect 36081 47951 36139 47957
rect 36262 47948 36268 48000
rect 36320 47948 36326 48000
rect 36832 47988 36860 48096
rect 49326 48084 49332 48136
rect 49384 48084 49390 48136
rect 39022 47988 39028 48000
rect 36832 47960 39028 47988
rect 39022 47948 39028 47960
rect 39080 47948 39086 48000
rect 43346 47948 43352 48000
rect 43404 47988 43410 48000
rect 49145 47991 49203 47997
rect 49145 47988 49157 47991
rect 43404 47960 49157 47988
rect 43404 47948 43410 47960
rect 49145 47957 49157 47960
rect 49191 47957 49203 47991
rect 49145 47951 49203 47957
rect 1104 47898 49864 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 27950 47898
rect 28002 47846 28014 47898
rect 28066 47846 28078 47898
rect 28130 47846 28142 47898
rect 28194 47846 28206 47898
rect 28258 47846 37950 47898
rect 38002 47846 38014 47898
rect 38066 47846 38078 47898
rect 38130 47846 38142 47898
rect 38194 47846 38206 47898
rect 38258 47846 47950 47898
rect 48002 47846 48014 47898
rect 48066 47846 48078 47898
rect 48130 47846 48142 47898
rect 48194 47846 48206 47898
rect 48258 47846 49864 47898
rect 1104 47824 49864 47846
rect 10686 47744 10692 47796
rect 10744 47784 10750 47796
rect 12253 47787 12311 47793
rect 12253 47784 12265 47787
rect 10744 47756 12265 47784
rect 10744 47744 10750 47756
rect 12253 47753 12265 47756
rect 12299 47753 12311 47787
rect 12253 47747 12311 47753
rect 19996 47756 21312 47784
rect 19518 47676 19524 47728
rect 19576 47716 19582 47728
rect 19996 47725 20024 47756
rect 19981 47719 20039 47725
rect 19981 47716 19993 47719
rect 19576 47688 19993 47716
rect 19576 47676 19582 47688
rect 19981 47685 19993 47688
rect 20027 47685 20039 47719
rect 19981 47679 20039 47685
rect 1765 47651 1823 47657
rect 1765 47617 1777 47651
rect 1811 47648 1823 47651
rect 4062 47648 4068 47660
rect 1811 47620 4068 47648
rect 1811 47617 1823 47620
rect 1765 47611 1823 47617
rect 4062 47608 4068 47620
rect 4120 47608 4126 47660
rect 12437 47651 12495 47657
rect 12437 47617 12449 47651
rect 12483 47648 12495 47651
rect 15102 47648 15108 47660
rect 12483 47620 15108 47648
rect 12483 47617 12495 47620
rect 12437 47611 12495 47617
rect 15102 47608 15108 47620
rect 15160 47608 15166 47660
rect 21082 47608 21088 47660
rect 21140 47608 21146 47660
rect 1302 47540 1308 47592
rect 1360 47580 1366 47592
rect 2041 47583 2099 47589
rect 2041 47580 2053 47583
rect 1360 47552 2053 47580
rect 1360 47540 1366 47552
rect 2041 47549 2053 47552
rect 2087 47549 2099 47583
rect 2041 47543 2099 47549
rect 19702 47540 19708 47592
rect 19760 47540 19766 47592
rect 21284 47580 21312 47756
rect 21450 47744 21456 47796
rect 21508 47744 21514 47796
rect 22002 47744 22008 47796
rect 22060 47744 22066 47796
rect 22186 47744 22192 47796
rect 22244 47784 22250 47796
rect 24949 47787 25007 47793
rect 24949 47784 24961 47787
rect 22244 47756 24961 47784
rect 22244 47744 22250 47756
rect 24949 47753 24961 47756
rect 24995 47784 25007 47787
rect 25682 47784 25688 47796
rect 24995 47756 25688 47784
rect 24995 47753 25007 47756
rect 24949 47747 25007 47753
rect 25682 47744 25688 47756
rect 25740 47744 25746 47796
rect 26786 47784 26792 47796
rect 25792 47756 26792 47784
rect 22462 47676 22468 47728
rect 22520 47676 22526 47728
rect 25130 47676 25136 47728
rect 25188 47716 25194 47728
rect 25792 47716 25820 47756
rect 26786 47744 26792 47756
rect 26844 47744 26850 47796
rect 26896 47756 27739 47784
rect 25188 47688 25820 47716
rect 25869 47719 25927 47725
rect 25188 47676 25194 47688
rect 25869 47685 25881 47719
rect 25915 47716 25927 47719
rect 26896 47716 26924 47756
rect 25915 47688 26924 47716
rect 27525 47719 27583 47725
rect 25915 47685 25927 47688
rect 25869 47679 25927 47685
rect 27525 47685 27537 47719
rect 27571 47685 27583 47719
rect 27525 47679 27583 47685
rect 22373 47651 22431 47657
rect 22373 47617 22385 47651
rect 22419 47648 22431 47651
rect 22830 47648 22836 47660
rect 22419 47620 22836 47648
rect 22419 47617 22431 47620
rect 22373 47611 22431 47617
rect 22830 47608 22836 47620
rect 22888 47608 22894 47660
rect 24578 47608 24584 47660
rect 24636 47648 24642 47660
rect 25498 47648 25504 47660
rect 24636 47620 25504 47648
rect 24636 47608 24642 47620
rect 25498 47608 25504 47620
rect 25556 47648 25562 47660
rect 25682 47648 25688 47660
rect 25556 47620 25688 47648
rect 25556 47608 25562 47620
rect 25682 47608 25688 47620
rect 25740 47608 25746 47660
rect 25777 47651 25835 47657
rect 25777 47617 25789 47651
rect 25823 47648 25835 47651
rect 26234 47648 26240 47660
rect 25823 47620 26240 47648
rect 25823 47617 25835 47620
rect 25777 47611 25835 47617
rect 26234 47608 26240 47620
rect 26292 47608 26298 47660
rect 27540 47648 27568 47679
rect 27614 47676 27620 47728
rect 27672 47676 27678 47728
rect 27711 47716 27739 47756
rect 28258 47744 28264 47796
rect 28316 47784 28322 47796
rect 29362 47784 29368 47796
rect 28316 47756 29368 47784
rect 28316 47744 28322 47756
rect 29362 47744 29368 47756
rect 29420 47744 29426 47796
rect 31754 47784 31760 47796
rect 29472 47756 31760 47784
rect 28994 47716 29000 47728
rect 27711 47688 29000 47716
rect 28994 47676 29000 47688
rect 29052 47676 29058 47728
rect 28350 47648 28356 47660
rect 27540 47620 28356 47648
rect 28350 47608 28356 47620
rect 28408 47608 28414 47660
rect 29472 47657 29500 47756
rect 31754 47744 31760 47756
rect 31812 47784 31818 47796
rect 31938 47784 31944 47796
rect 31812 47756 31944 47784
rect 31812 47744 31818 47756
rect 31938 47744 31944 47756
rect 31996 47784 32002 47796
rect 31996 47756 32996 47784
rect 31996 47744 32002 47756
rect 31294 47716 31300 47728
rect 30958 47688 31300 47716
rect 31294 47676 31300 47688
rect 31352 47716 31358 47728
rect 32122 47716 32128 47728
rect 31352 47688 32128 47716
rect 31352 47676 31358 47688
rect 32122 47676 32128 47688
rect 32180 47676 32186 47728
rect 32968 47657 32996 47756
rect 34790 47744 34796 47796
rect 34848 47784 34854 47796
rect 35161 47787 35219 47793
rect 35161 47784 35173 47787
rect 34848 47756 35173 47784
rect 34848 47744 34854 47756
rect 35161 47753 35173 47756
rect 35207 47753 35219 47787
rect 35161 47747 35219 47753
rect 35529 47787 35587 47793
rect 35529 47753 35541 47787
rect 35575 47784 35587 47787
rect 38289 47787 38347 47793
rect 38289 47784 38301 47787
rect 35575 47756 38301 47784
rect 35575 47753 35587 47756
rect 35529 47747 35587 47753
rect 38289 47753 38301 47756
rect 38335 47753 38347 47787
rect 38289 47747 38347 47753
rect 38657 47787 38715 47793
rect 38657 47753 38669 47787
rect 38703 47784 38715 47787
rect 42794 47784 42800 47796
rect 38703 47756 42800 47784
rect 38703 47753 38715 47756
rect 38657 47747 38715 47753
rect 42794 47744 42800 47756
rect 42852 47744 42858 47796
rect 33229 47719 33287 47725
rect 33229 47685 33241 47719
rect 33275 47716 33287 47719
rect 33502 47716 33508 47728
rect 33275 47688 33508 47716
rect 33275 47685 33287 47688
rect 33229 47679 33287 47685
rect 33502 47676 33508 47688
rect 33560 47676 33566 47728
rect 33778 47676 33784 47728
rect 33836 47676 33842 47728
rect 40126 47676 40132 47728
rect 40184 47716 40190 47728
rect 48866 47716 48872 47728
rect 40184 47688 48872 47716
rect 40184 47676 40190 47688
rect 48866 47676 48872 47688
rect 48924 47676 48930 47728
rect 29457 47651 29515 47657
rect 29457 47617 29469 47651
rect 29503 47617 29515 47651
rect 29457 47611 29515 47617
rect 32953 47651 33011 47657
rect 32953 47617 32965 47651
rect 32999 47617 33011 47651
rect 32953 47611 33011 47617
rect 35250 47608 35256 47660
rect 35308 47648 35314 47660
rect 37550 47648 37556 47660
rect 35308 47620 37556 47648
rect 35308 47608 35314 47620
rect 37550 47608 37556 47620
rect 37608 47608 37614 47660
rect 38749 47651 38807 47657
rect 38749 47617 38761 47651
rect 38795 47648 38807 47651
rect 39758 47648 39764 47660
rect 38795 47620 39764 47648
rect 38795 47617 38807 47620
rect 38749 47611 38807 47617
rect 39758 47608 39764 47620
rect 39816 47648 39822 47660
rect 48682 47648 48688 47660
rect 39816 47620 48688 47648
rect 39816 47608 39822 47620
rect 48682 47608 48688 47620
rect 48740 47608 48746 47660
rect 49326 47608 49332 47660
rect 49384 47608 49390 47660
rect 22646 47580 22652 47592
rect 21284 47552 22652 47580
rect 22646 47540 22652 47552
rect 22704 47540 22710 47592
rect 23201 47583 23259 47589
rect 23201 47549 23213 47583
rect 23247 47549 23259 47583
rect 23201 47543 23259 47549
rect 23477 47583 23535 47589
rect 23477 47549 23489 47583
rect 23523 47580 23535 47583
rect 23566 47580 23572 47592
rect 23523 47552 23572 47580
rect 23523 47549 23535 47552
rect 23477 47543 23535 47549
rect 22094 47472 22100 47524
rect 22152 47512 22158 47524
rect 23216 47512 23244 47543
rect 23566 47540 23572 47552
rect 23624 47580 23630 47592
rect 24762 47580 24768 47592
rect 23624 47552 24768 47580
rect 23624 47540 23630 47552
rect 24762 47540 24768 47552
rect 24820 47540 24826 47592
rect 26053 47583 26111 47589
rect 26053 47549 26065 47583
rect 26099 47580 26111 47583
rect 27430 47580 27436 47592
rect 26099 47552 27436 47580
rect 26099 47549 26111 47552
rect 26053 47543 26111 47549
rect 27430 47540 27436 47552
rect 27488 47540 27494 47592
rect 27709 47583 27767 47589
rect 27709 47549 27721 47583
rect 27755 47549 27767 47583
rect 27709 47543 27767 47549
rect 27157 47515 27215 47521
rect 27157 47512 27169 47515
rect 22152 47484 23244 47512
rect 24504 47484 27169 47512
rect 22152 47472 22158 47484
rect 21266 47404 21272 47456
rect 21324 47444 21330 47456
rect 24504 47444 24532 47484
rect 27157 47481 27169 47484
rect 27203 47481 27215 47515
rect 27157 47475 27215 47481
rect 27246 47472 27252 47524
rect 27304 47512 27310 47524
rect 27724 47512 27752 47543
rect 29362 47540 29368 47592
rect 29420 47580 29426 47592
rect 29733 47583 29791 47589
rect 29733 47580 29745 47583
rect 29420 47552 29745 47580
rect 29420 47540 29426 47552
rect 29733 47549 29745 47552
rect 29779 47580 29791 47583
rect 29779 47552 30788 47580
rect 29779 47549 29791 47552
rect 29733 47543 29791 47549
rect 27304 47484 27752 47512
rect 30760 47512 30788 47552
rect 31018 47540 31024 47592
rect 31076 47580 31082 47592
rect 31205 47583 31263 47589
rect 31205 47580 31217 47583
rect 31076 47552 31217 47580
rect 31076 47540 31082 47552
rect 31205 47549 31217 47552
rect 31251 47549 31263 47583
rect 31205 47543 31263 47549
rect 31726 47552 34284 47580
rect 31726 47524 31754 47552
rect 31726 47512 31760 47524
rect 30760 47484 31760 47512
rect 27304 47472 27310 47484
rect 31754 47472 31760 47484
rect 31812 47472 31818 47524
rect 31846 47472 31852 47524
rect 31904 47512 31910 47524
rect 32122 47512 32128 47524
rect 31904 47484 32128 47512
rect 31904 47472 31910 47484
rect 32122 47472 32128 47484
rect 32180 47512 32186 47524
rect 32766 47512 32772 47524
rect 32180 47484 32772 47512
rect 32180 47472 32186 47484
rect 32766 47472 32772 47484
rect 32824 47472 32830 47524
rect 34256 47512 34284 47552
rect 34882 47540 34888 47592
rect 34940 47580 34946 47592
rect 35621 47583 35679 47589
rect 35621 47580 35633 47583
rect 34940 47552 35633 47580
rect 34940 47540 34946 47552
rect 35621 47549 35633 47552
rect 35667 47549 35679 47583
rect 35621 47543 35679 47549
rect 35713 47583 35771 47589
rect 35713 47549 35725 47583
rect 35759 47549 35771 47583
rect 35713 47543 35771 47549
rect 35728 47512 35756 47543
rect 35802 47540 35808 47592
rect 35860 47580 35866 47592
rect 38930 47580 38936 47592
rect 35860 47552 38936 47580
rect 35860 47540 35866 47552
rect 38930 47540 38936 47552
rect 38988 47540 38994 47592
rect 34256 47484 35756 47512
rect 21324 47416 24532 47444
rect 21324 47404 21330 47416
rect 25130 47404 25136 47456
rect 25188 47444 25194 47456
rect 25409 47447 25467 47453
rect 25409 47444 25421 47447
rect 25188 47416 25421 47444
rect 25188 47404 25194 47416
rect 25409 47413 25421 47416
rect 25455 47413 25467 47447
rect 25409 47407 25467 47413
rect 25498 47404 25504 47456
rect 25556 47444 25562 47456
rect 30190 47444 30196 47456
rect 25556 47416 30196 47444
rect 25556 47404 25562 47416
rect 30190 47404 30196 47416
rect 30248 47404 30254 47456
rect 34606 47404 34612 47456
rect 34664 47444 34670 47456
rect 34701 47447 34759 47453
rect 34701 47444 34713 47447
rect 34664 47416 34713 47444
rect 34664 47404 34670 47416
rect 34701 47413 34713 47416
rect 34747 47413 34759 47447
rect 34701 47407 34759 47413
rect 34974 47404 34980 47456
rect 35032 47444 35038 47456
rect 35710 47444 35716 47456
rect 35032 47416 35716 47444
rect 35032 47404 35038 47416
rect 35710 47404 35716 47416
rect 35768 47444 35774 47456
rect 37458 47444 37464 47456
rect 35768 47416 37464 47444
rect 35768 47404 35774 47416
rect 37458 47404 37464 47416
rect 37516 47444 37522 47456
rect 37826 47444 37832 47456
rect 37516 47416 37832 47444
rect 37516 47404 37522 47416
rect 37826 47404 37832 47416
rect 37884 47404 37890 47456
rect 42794 47404 42800 47456
rect 42852 47444 42858 47456
rect 49145 47447 49203 47453
rect 49145 47444 49157 47447
rect 42852 47416 49157 47444
rect 42852 47404 42858 47416
rect 49145 47413 49157 47416
rect 49191 47413 49203 47447
rect 49145 47407 49203 47413
rect 1104 47354 49864 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 32950 47354
rect 33002 47302 33014 47354
rect 33066 47302 33078 47354
rect 33130 47302 33142 47354
rect 33194 47302 33206 47354
rect 33258 47302 42950 47354
rect 43002 47302 43014 47354
rect 43066 47302 43078 47354
rect 43130 47302 43142 47354
rect 43194 47302 43206 47354
rect 43258 47302 49864 47354
rect 1104 47280 49864 47302
rect 15194 47200 15200 47252
rect 15252 47240 15258 47252
rect 18141 47243 18199 47249
rect 18141 47240 18153 47243
rect 15252 47212 18153 47240
rect 15252 47200 15258 47212
rect 18141 47209 18153 47212
rect 18187 47209 18199 47243
rect 18141 47203 18199 47209
rect 22830 47200 22836 47252
rect 22888 47240 22894 47252
rect 24949 47243 25007 47249
rect 24949 47240 24961 47243
rect 22888 47212 24961 47240
rect 22888 47200 22894 47212
rect 24949 47209 24961 47212
rect 24995 47209 25007 47243
rect 24949 47203 25007 47209
rect 25682 47200 25688 47252
rect 25740 47240 25746 47252
rect 26878 47240 26884 47252
rect 25740 47212 26884 47240
rect 25740 47200 25746 47212
rect 26878 47200 26884 47212
rect 26936 47200 26942 47252
rect 27522 47200 27528 47252
rect 27580 47240 27586 47252
rect 27893 47243 27951 47249
rect 27893 47240 27905 47243
rect 27580 47212 27905 47240
rect 27580 47200 27586 47212
rect 27893 47209 27905 47212
rect 27939 47209 27951 47243
rect 27893 47203 27951 47209
rect 28350 47200 28356 47252
rect 28408 47200 28414 47252
rect 28626 47200 28632 47252
rect 28684 47240 28690 47252
rect 28684 47212 30880 47240
rect 28684 47200 28690 47212
rect 19150 47132 19156 47184
rect 19208 47172 19214 47184
rect 20533 47175 20591 47181
rect 20533 47172 20545 47175
rect 19208 47144 20545 47172
rect 19208 47132 19214 47144
rect 20533 47141 20545 47144
rect 20579 47141 20591 47175
rect 22186 47172 22192 47184
rect 20533 47135 20591 47141
rect 21192 47144 22192 47172
rect 18785 47107 18843 47113
rect 18785 47073 18797 47107
rect 18831 47104 18843 47107
rect 20898 47104 20904 47116
rect 18831 47076 20904 47104
rect 18831 47073 18843 47076
rect 18785 47067 18843 47073
rect 20898 47064 20904 47076
rect 20956 47064 20962 47116
rect 21192 47113 21220 47144
rect 22186 47132 22192 47144
rect 22244 47132 22250 47184
rect 23937 47175 23995 47181
rect 23937 47141 23949 47175
rect 23983 47172 23995 47175
rect 25498 47172 25504 47184
rect 23983 47144 25504 47172
rect 23983 47141 23995 47144
rect 23937 47135 23995 47141
rect 21177 47107 21235 47113
rect 21177 47073 21189 47107
rect 21223 47073 21235 47107
rect 21177 47067 21235 47073
rect 21450 47064 21456 47116
rect 21508 47104 21514 47116
rect 22465 47107 22523 47113
rect 22465 47104 22477 47107
rect 21508 47076 22477 47104
rect 21508 47064 21514 47076
rect 22465 47073 22477 47076
rect 22511 47073 22523 47107
rect 22465 47067 22523 47073
rect 18509 47039 18567 47045
rect 18509 47005 18521 47039
rect 18555 47036 18567 47039
rect 20073 47039 20131 47045
rect 20073 47036 20085 47039
rect 18555 47008 20085 47036
rect 18555 47005 18567 47008
rect 18509 46999 18567 47005
rect 20073 47005 20085 47008
rect 20119 47005 20131 47039
rect 20073 46999 20131 47005
rect 20993 47039 21051 47045
rect 20993 47005 21005 47039
rect 21039 47036 21051 47039
rect 21266 47036 21272 47048
rect 21039 47008 21272 47036
rect 21039 47005 21051 47008
rect 20993 46999 21051 47005
rect 21266 46996 21272 47008
rect 21324 46996 21330 47048
rect 22094 46996 22100 47048
rect 22152 47036 22158 47048
rect 22189 47039 22247 47045
rect 22189 47036 22201 47039
rect 22152 47008 22201 47036
rect 22152 46996 22158 47008
rect 22189 47005 22201 47008
rect 22235 47005 22247 47039
rect 24780 47036 24808 47144
rect 25498 47132 25504 47144
rect 25556 47132 25562 47184
rect 27614 47132 27620 47184
rect 27672 47172 27678 47184
rect 29086 47172 29092 47184
rect 27672 47144 29092 47172
rect 27672 47132 27678 47144
rect 29086 47132 29092 47144
rect 29144 47172 29150 47184
rect 29270 47172 29276 47184
rect 29144 47144 29276 47172
rect 29144 47132 29150 47144
rect 29270 47132 29276 47144
rect 29328 47132 29334 47184
rect 29733 47175 29791 47181
rect 29733 47141 29745 47175
rect 29779 47172 29791 47175
rect 29822 47172 29828 47184
rect 29779 47144 29828 47172
rect 29779 47141 29791 47144
rect 29733 47135 29791 47141
rect 29822 47132 29828 47144
rect 29880 47132 29886 47184
rect 30852 47172 30880 47212
rect 30926 47200 30932 47252
rect 30984 47200 30990 47252
rect 34882 47200 34888 47252
rect 34940 47200 34946 47252
rect 37182 47200 37188 47252
rect 37240 47240 37246 47252
rect 38473 47243 38531 47249
rect 38473 47240 38485 47243
rect 37240 47212 38485 47240
rect 37240 47200 37246 47212
rect 38473 47209 38485 47212
rect 38519 47209 38531 47243
rect 38473 47203 38531 47209
rect 36081 47175 36139 47181
rect 30852 47144 33824 47172
rect 24854 47064 24860 47116
rect 24912 47104 24918 47116
rect 25593 47107 25651 47113
rect 25593 47104 25605 47107
rect 24912 47076 25605 47104
rect 24912 47064 24918 47076
rect 25593 47073 25605 47076
rect 25639 47104 25651 47107
rect 25866 47104 25872 47116
rect 25639 47076 25872 47104
rect 25639 47073 25651 47076
rect 25593 47067 25651 47073
rect 25866 47064 25872 47076
rect 25924 47064 25930 47116
rect 26050 47064 26056 47116
rect 26108 47104 26114 47116
rect 26145 47107 26203 47113
rect 26145 47104 26157 47107
rect 26108 47076 26157 47104
rect 26108 47064 26114 47076
rect 26145 47073 26157 47076
rect 26191 47073 26203 47107
rect 26145 47067 26203 47073
rect 26786 47064 26792 47116
rect 26844 47104 26850 47116
rect 28905 47107 28963 47113
rect 28905 47104 28917 47107
rect 26844 47076 28917 47104
rect 26844 47064 26850 47076
rect 28905 47073 28917 47076
rect 28951 47104 28963 47107
rect 29914 47104 29920 47116
rect 28951 47076 29920 47104
rect 28951 47073 28963 47076
rect 28905 47067 28963 47073
rect 29914 47064 29920 47076
rect 29972 47064 29978 47116
rect 30190 47064 30196 47116
rect 30248 47104 30254 47116
rect 30285 47107 30343 47113
rect 30285 47104 30297 47107
rect 30248 47076 30297 47104
rect 30248 47064 30254 47076
rect 30285 47073 30297 47076
rect 30331 47073 30343 47107
rect 30285 47067 30343 47073
rect 31018 47064 31024 47116
rect 31076 47104 31082 47116
rect 31389 47107 31447 47113
rect 31389 47104 31401 47107
rect 31076 47076 31401 47104
rect 31076 47064 31082 47076
rect 31389 47073 31401 47076
rect 31435 47073 31447 47107
rect 31389 47067 31447 47073
rect 31478 47064 31484 47116
rect 31536 47064 31542 47116
rect 32582 47064 32588 47116
rect 32640 47064 32646 47116
rect 32674 47064 32680 47116
rect 32732 47064 32738 47116
rect 33796 47113 33824 47144
rect 36081 47141 36093 47175
rect 36127 47172 36139 47175
rect 37090 47172 37096 47184
rect 36127 47144 37096 47172
rect 36127 47141 36139 47144
rect 36081 47135 36139 47141
rect 37090 47132 37096 47144
rect 37148 47132 37154 47184
rect 33781 47107 33839 47113
rect 33781 47073 33793 47107
rect 33827 47073 33839 47107
rect 33781 47067 33839 47073
rect 33870 47064 33876 47116
rect 33928 47104 33934 47116
rect 33965 47107 34023 47113
rect 33965 47104 33977 47107
rect 33928 47076 33977 47104
rect 33928 47064 33934 47076
rect 33965 47073 33977 47076
rect 34011 47104 34023 47107
rect 34330 47104 34336 47116
rect 34011 47076 34336 47104
rect 34011 47073 34023 47076
rect 33965 47067 34023 47073
rect 34330 47064 34336 47076
rect 34388 47064 34394 47116
rect 34422 47064 34428 47116
rect 34480 47104 34486 47116
rect 35529 47107 35587 47113
rect 35529 47104 35541 47107
rect 34480 47076 35541 47104
rect 34480 47064 34486 47076
rect 35529 47073 35541 47076
rect 35575 47104 35587 47107
rect 35802 47104 35808 47116
rect 35575 47076 35808 47104
rect 35575 47073 35587 47076
rect 35529 47067 35587 47073
rect 35802 47064 35808 47076
rect 35860 47064 35866 47116
rect 36538 47064 36544 47116
rect 36596 47064 36602 47116
rect 36630 47064 36636 47116
rect 36688 47064 36694 47116
rect 39022 47064 39028 47116
rect 39080 47064 39086 47116
rect 24946 47036 24952 47048
rect 24780 47008 24952 47036
rect 22189 46999 22247 47005
rect 24946 46996 24952 47008
rect 25004 46996 25010 47048
rect 25314 46996 25320 47048
rect 25372 46996 25378 47048
rect 28721 47039 28779 47045
rect 28721 47005 28733 47039
rect 28767 47036 28779 47039
rect 28810 47036 28816 47048
rect 28767 47008 28816 47036
rect 28767 47005 28779 47008
rect 28721 46999 28779 47005
rect 28810 46996 28816 47008
rect 28868 46996 28874 47048
rect 30466 46996 30472 47048
rect 30524 47036 30530 47048
rect 32493 47039 32551 47045
rect 32493 47036 32505 47039
rect 30524 47008 32505 47036
rect 30524 46996 30530 47008
rect 32493 47005 32505 47008
rect 32539 47005 32551 47039
rect 32493 46999 32551 47005
rect 33686 46996 33692 47048
rect 33744 46996 33750 47048
rect 34698 46996 34704 47048
rect 34756 47036 34762 47048
rect 35250 47036 35256 47048
rect 34756 47008 35256 47036
rect 34756 46996 34762 47008
rect 35250 46996 35256 47008
rect 35308 46996 35314 47048
rect 35345 47039 35403 47045
rect 35345 47005 35357 47039
rect 35391 47036 35403 47039
rect 38286 47036 38292 47048
rect 35391 47008 38292 47036
rect 35391 47005 35403 47008
rect 35345 46999 35403 47005
rect 38286 46996 38292 47008
rect 38344 46996 38350 47048
rect 38841 47039 38899 47045
rect 38841 47005 38853 47039
rect 38887 47036 38899 47039
rect 43438 47036 43444 47048
rect 38887 47008 43444 47036
rect 38887 47005 38899 47008
rect 38841 46999 38899 47005
rect 43438 46996 43444 47008
rect 43496 46996 43502 47048
rect 18601 46971 18659 46977
rect 18601 46937 18613 46971
rect 18647 46968 18659 46971
rect 20714 46968 20720 46980
rect 18647 46940 20720 46968
rect 18647 46937 18659 46940
rect 18601 46931 18659 46937
rect 20714 46928 20720 46940
rect 20772 46928 20778 46980
rect 20901 46971 20959 46977
rect 20901 46937 20913 46971
rect 20947 46968 20959 46971
rect 22002 46968 22008 46980
rect 20947 46940 22008 46968
rect 20947 46937 20959 46940
rect 20901 46931 20959 46937
rect 22002 46928 22008 46940
rect 22060 46928 22066 46980
rect 23842 46968 23848 46980
rect 23690 46940 23848 46968
rect 23842 46928 23848 46940
rect 23900 46968 23906 46980
rect 24578 46968 24584 46980
rect 23900 46940 24584 46968
rect 23900 46928 23906 46940
rect 24578 46928 24584 46940
rect 24636 46928 24642 46980
rect 25409 46971 25467 46977
rect 25409 46937 25421 46971
rect 25455 46968 25467 46971
rect 25774 46968 25780 46980
rect 25455 46940 25780 46968
rect 25455 46937 25467 46940
rect 25409 46931 25467 46937
rect 25774 46928 25780 46940
rect 25832 46968 25838 46980
rect 26142 46968 26148 46980
rect 25832 46940 26148 46968
rect 25832 46928 25838 46940
rect 26142 46928 26148 46940
rect 26200 46928 26206 46980
rect 26421 46971 26479 46977
rect 26421 46937 26433 46971
rect 26467 46968 26479 46971
rect 26467 46940 26832 46968
rect 26467 46937 26479 46940
rect 26421 46931 26479 46937
rect 21174 46860 21180 46912
rect 21232 46900 21238 46912
rect 23474 46900 23480 46912
rect 21232 46872 23480 46900
rect 21232 46860 21238 46872
rect 23474 46860 23480 46872
rect 23532 46860 23538 46912
rect 26804 46900 26832 46940
rect 26878 46928 26884 46980
rect 26936 46928 26942 46980
rect 28350 46968 28356 46980
rect 27724 46940 28356 46968
rect 27724 46900 27752 46940
rect 28350 46928 28356 46940
rect 28408 46928 28414 46980
rect 28534 46928 28540 46980
rect 28592 46968 28598 46980
rect 30101 46971 30159 46977
rect 30101 46968 30113 46971
rect 28592 46940 30113 46968
rect 28592 46928 28598 46940
rect 30101 46937 30113 46940
rect 30147 46937 30159 46971
rect 30101 46931 30159 46937
rect 30193 46971 30251 46977
rect 30193 46937 30205 46971
rect 30239 46968 30251 46971
rect 30282 46968 30288 46980
rect 30239 46940 30288 46968
rect 30239 46937 30251 46940
rect 30193 46931 30251 46937
rect 30282 46928 30288 46940
rect 30340 46928 30346 46980
rect 30558 46928 30564 46980
rect 30616 46968 30622 46980
rect 31297 46971 31355 46977
rect 31297 46968 31309 46971
rect 30616 46940 31309 46968
rect 30616 46928 30622 46940
rect 31297 46937 31309 46940
rect 31343 46937 31355 46971
rect 36078 46968 36084 46980
rect 31297 46931 31355 46937
rect 32140 46940 36084 46968
rect 26804 46872 27752 46900
rect 28626 46860 28632 46912
rect 28684 46900 28690 46912
rect 28813 46903 28871 46909
rect 28813 46900 28825 46903
rect 28684 46872 28825 46900
rect 28684 46860 28690 46872
rect 28813 46869 28825 46872
rect 28859 46869 28871 46903
rect 28813 46863 28871 46869
rect 29086 46860 29092 46912
rect 29144 46900 29150 46912
rect 31570 46900 31576 46912
rect 29144 46872 31576 46900
rect 29144 46860 29150 46872
rect 31570 46860 31576 46872
rect 31628 46860 31634 46912
rect 32140 46909 32168 46940
rect 36078 46928 36084 46940
rect 36136 46928 36142 46980
rect 36446 46928 36452 46980
rect 36504 46928 36510 46980
rect 38933 46971 38991 46977
rect 38933 46937 38945 46971
rect 38979 46968 38991 46971
rect 40126 46968 40132 46980
rect 38979 46940 40132 46968
rect 38979 46937 38991 46940
rect 38933 46931 38991 46937
rect 40126 46928 40132 46940
rect 40184 46928 40190 46980
rect 32125 46903 32183 46909
rect 32125 46869 32137 46903
rect 32171 46869 32183 46903
rect 32125 46863 32183 46869
rect 33318 46860 33324 46912
rect 33376 46860 33382 46912
rect 1104 46810 49864 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 27950 46810
rect 28002 46758 28014 46810
rect 28066 46758 28078 46810
rect 28130 46758 28142 46810
rect 28194 46758 28206 46810
rect 28258 46758 37950 46810
rect 38002 46758 38014 46810
rect 38066 46758 38078 46810
rect 38130 46758 38142 46810
rect 38194 46758 38206 46810
rect 38258 46758 47950 46810
rect 48002 46758 48014 46810
rect 48066 46758 48078 46810
rect 48130 46758 48142 46810
rect 48194 46758 48206 46810
rect 48258 46758 49864 46810
rect 1104 46736 49864 46758
rect 10962 46656 10968 46708
rect 11020 46696 11026 46708
rect 11977 46699 12035 46705
rect 11977 46696 11989 46699
rect 11020 46668 11989 46696
rect 11020 46656 11026 46668
rect 11977 46665 11989 46668
rect 12023 46665 12035 46699
rect 11977 46659 12035 46665
rect 22554 46656 22560 46708
rect 22612 46696 22618 46708
rect 23753 46699 23811 46705
rect 23753 46696 23765 46699
rect 22612 46668 23765 46696
rect 22612 46656 22618 46668
rect 23753 46665 23765 46668
rect 23799 46696 23811 46699
rect 24762 46696 24768 46708
rect 23799 46668 24768 46696
rect 23799 46665 23811 46668
rect 23753 46659 23811 46665
rect 24762 46656 24768 46668
rect 24820 46656 24826 46708
rect 26050 46696 26056 46708
rect 24872 46668 26056 46696
rect 21634 46588 21640 46640
rect 21692 46628 21698 46640
rect 22281 46631 22339 46637
rect 22281 46628 22293 46631
rect 21692 46600 22293 46628
rect 21692 46588 21698 46600
rect 22281 46597 22293 46600
rect 22327 46597 22339 46631
rect 23842 46628 23848 46640
rect 23506 46600 23848 46628
rect 22281 46591 22339 46597
rect 23842 46588 23848 46600
rect 23900 46588 23906 46640
rect 24670 46588 24676 46640
rect 24728 46628 24734 46640
rect 24872 46628 24900 46668
rect 26050 46656 26056 46668
rect 26108 46656 26114 46708
rect 26605 46699 26663 46705
rect 26605 46665 26617 46699
rect 26651 46696 26663 46699
rect 26786 46696 26792 46708
rect 26651 46668 26792 46696
rect 26651 46665 26663 46668
rect 26605 46659 26663 46665
rect 26786 46656 26792 46668
rect 26844 46656 26850 46708
rect 27985 46699 28043 46705
rect 27985 46665 27997 46699
rect 28031 46696 28043 46699
rect 28902 46696 28908 46708
rect 28031 46668 28908 46696
rect 28031 46665 28043 46668
rect 27985 46659 28043 46665
rect 28902 46656 28908 46668
rect 28960 46656 28966 46708
rect 29178 46656 29184 46708
rect 29236 46656 29242 46708
rect 29273 46699 29331 46705
rect 29273 46665 29285 46699
rect 29319 46696 29331 46699
rect 29454 46696 29460 46708
rect 29319 46668 29460 46696
rect 29319 46665 29331 46668
rect 29273 46659 29331 46665
rect 29454 46656 29460 46668
rect 29512 46656 29518 46708
rect 32582 46696 32588 46708
rect 30300 46668 32588 46696
rect 24728 46600 24900 46628
rect 24728 46588 24734 46600
rect 24872 46572 24900 46600
rect 25682 46588 25688 46640
rect 25740 46588 25746 46640
rect 27890 46588 27896 46640
rect 27948 46628 27954 46640
rect 28534 46628 28540 46640
rect 27948 46600 28540 46628
rect 27948 46588 27954 46600
rect 28534 46588 28540 46600
rect 28592 46588 28598 46640
rect 28626 46588 28632 46640
rect 28684 46628 28690 46640
rect 30300 46637 30328 46668
rect 32582 46656 32588 46668
rect 32640 46656 32646 46708
rect 32677 46699 32735 46705
rect 32677 46665 32689 46699
rect 32723 46696 32735 46699
rect 33686 46696 33692 46708
rect 32723 46668 33692 46696
rect 32723 46665 32735 46668
rect 32677 46659 32735 46665
rect 30285 46631 30343 46637
rect 30285 46628 30297 46631
rect 28684 46600 30297 46628
rect 28684 46588 28690 46600
rect 30285 46597 30297 46600
rect 30331 46597 30343 46631
rect 30285 46591 30343 46597
rect 31294 46588 31300 46640
rect 31352 46588 31358 46640
rect 31662 46588 31668 46640
rect 31720 46628 31726 46640
rect 32692 46628 32720 46659
rect 33686 46656 33692 46668
rect 33744 46656 33750 46708
rect 36538 46628 36544 46640
rect 31720 46600 32720 46628
rect 36018 46600 36544 46628
rect 31720 46588 31726 46600
rect 36538 46588 36544 46600
rect 36596 46628 36602 46640
rect 39298 46628 39304 46640
rect 36596 46600 39304 46628
rect 36596 46588 36602 46600
rect 39298 46588 39304 46600
rect 39356 46588 39362 46640
rect 1765 46563 1823 46569
rect 1765 46529 1777 46563
rect 1811 46560 1823 46563
rect 8662 46560 8668 46572
rect 1811 46532 8668 46560
rect 1811 46529 1823 46532
rect 1765 46523 1823 46529
rect 8662 46520 8668 46532
rect 8720 46520 8726 46572
rect 12161 46563 12219 46569
rect 12161 46529 12173 46563
rect 12207 46560 12219 46563
rect 13722 46560 13728 46572
rect 12207 46532 13728 46560
rect 12207 46529 12219 46532
rect 12161 46523 12219 46529
rect 13722 46520 13728 46532
rect 13780 46520 13786 46572
rect 21082 46520 21088 46572
rect 21140 46520 21146 46572
rect 24854 46520 24860 46572
rect 24912 46520 24918 46572
rect 26436 46532 29684 46560
rect 1302 46452 1308 46504
rect 1360 46492 1366 46504
rect 2041 46495 2099 46501
rect 2041 46492 2053 46495
rect 1360 46464 2053 46492
rect 1360 46452 1366 46464
rect 2041 46461 2053 46464
rect 2087 46461 2099 46495
rect 2041 46455 2099 46461
rect 19702 46452 19708 46504
rect 19760 46452 19766 46504
rect 19981 46495 20039 46501
rect 19981 46461 19993 46495
rect 20027 46492 20039 46495
rect 21174 46492 21180 46504
rect 20027 46464 21180 46492
rect 20027 46461 20039 46464
rect 19981 46455 20039 46461
rect 21174 46452 21180 46464
rect 21232 46452 21238 46504
rect 22005 46495 22063 46501
rect 22005 46461 22017 46495
rect 22051 46492 22063 46495
rect 22051 46464 22140 46492
rect 22051 46461 22063 46464
rect 22005 46455 22063 46461
rect 22112 46368 22140 46464
rect 22830 46452 22836 46504
rect 22888 46492 22894 46504
rect 25133 46495 25191 46501
rect 25133 46492 25145 46495
rect 22888 46464 25145 46492
rect 22888 46452 22894 46464
rect 25133 46461 25145 46464
rect 25179 46492 25191 46495
rect 25866 46492 25872 46504
rect 25179 46464 25872 46492
rect 25179 46461 25191 46464
rect 25133 46455 25191 46461
rect 25866 46452 25872 46464
rect 25924 46452 25930 46504
rect 26142 46452 26148 46504
rect 26200 46492 26206 46504
rect 26436 46492 26464 46532
rect 26200 46464 26464 46492
rect 28169 46495 28227 46501
rect 26200 46452 26206 46464
rect 28169 46461 28181 46495
rect 28215 46492 28227 46495
rect 29086 46492 29092 46504
rect 28215 46464 29092 46492
rect 28215 46461 28227 46464
rect 28169 46455 28227 46461
rect 27522 46384 27528 46436
rect 27580 46384 27586 46436
rect 21453 46359 21511 46365
rect 21453 46325 21465 46359
rect 21499 46356 21511 46359
rect 21634 46356 21640 46368
rect 21499 46328 21640 46356
rect 21499 46325 21511 46328
rect 21453 46319 21511 46325
rect 21634 46316 21640 46328
rect 21692 46316 21698 46368
rect 22094 46316 22100 46368
rect 22152 46316 22158 46368
rect 22646 46316 22652 46368
rect 22704 46356 22710 46368
rect 25222 46356 25228 46368
rect 22704 46328 25228 46356
rect 22704 46316 22710 46328
rect 25222 46316 25228 46328
rect 25280 46316 25286 46368
rect 25314 46316 25320 46368
rect 25372 46356 25378 46368
rect 28184 46356 28212 46455
rect 29086 46452 29092 46464
rect 29144 46452 29150 46504
rect 29457 46495 29515 46501
rect 29457 46461 29469 46495
rect 29503 46492 29515 46495
rect 29656 46492 29684 46532
rect 30006 46520 30012 46572
rect 30064 46520 30070 46572
rect 31846 46520 31852 46572
rect 31904 46560 31910 46572
rect 32490 46560 32496 46572
rect 31904 46532 32496 46560
rect 31904 46520 31910 46532
rect 32490 46520 32496 46532
rect 32548 46560 32554 46572
rect 32548 46532 32904 46560
rect 32548 46520 32554 46532
rect 30834 46492 30840 46504
rect 29503 46464 29592 46492
rect 29656 46464 30840 46492
rect 29503 46461 29515 46464
rect 29457 46455 29515 46461
rect 25372 46328 28212 46356
rect 28813 46359 28871 46365
rect 25372 46316 25378 46328
rect 28813 46325 28825 46359
rect 28859 46356 28871 46359
rect 28902 46356 28908 46368
rect 28859 46328 28908 46356
rect 28859 46325 28871 46328
rect 28813 46319 28871 46325
rect 28902 46316 28908 46328
rect 28960 46316 28966 46368
rect 29564 46356 29592 46464
rect 30834 46452 30840 46464
rect 30892 46452 30898 46504
rect 31754 46452 31760 46504
rect 31812 46452 31818 46504
rect 32766 46452 32772 46504
rect 32824 46452 32830 46504
rect 32876 46501 32904 46532
rect 34514 46520 34520 46572
rect 34572 46520 34578 46572
rect 49050 46520 49056 46572
rect 49108 46520 49114 46572
rect 32861 46495 32919 46501
rect 32861 46461 32873 46495
rect 32907 46461 32919 46495
rect 32861 46455 32919 46461
rect 34790 46452 34796 46504
rect 34848 46452 34854 46504
rect 35342 46452 35348 46504
rect 35400 46492 35406 46504
rect 36265 46495 36323 46501
rect 36265 46492 36277 46495
rect 35400 46464 36277 46492
rect 35400 46452 35406 46464
rect 36265 46461 36277 46464
rect 36311 46461 36323 46495
rect 36265 46455 36323 46461
rect 49237 46427 49295 46433
rect 49237 46424 49249 46427
rect 31726 46396 34652 46424
rect 30282 46356 30288 46368
rect 29564 46328 30288 46356
rect 30282 46316 30288 46328
rect 30340 46316 30346 46368
rect 30466 46316 30472 46368
rect 30524 46356 30530 46368
rect 31726 46356 31754 46396
rect 30524 46328 31754 46356
rect 30524 46316 30530 46328
rect 32306 46316 32312 46368
rect 32364 46316 32370 46368
rect 32582 46316 32588 46368
rect 32640 46356 32646 46368
rect 34422 46356 34428 46368
rect 32640 46328 34428 46356
rect 32640 46316 32646 46328
rect 34422 46316 34428 46328
rect 34480 46316 34486 46368
rect 34624 46356 34652 46396
rect 35820 46396 49249 46424
rect 35820 46356 35848 46396
rect 49237 46393 49249 46396
rect 49283 46393 49295 46427
rect 49237 46387 49295 46393
rect 34624 46328 35848 46356
rect 1104 46266 49864 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 32950 46266
rect 33002 46214 33014 46266
rect 33066 46214 33078 46266
rect 33130 46214 33142 46266
rect 33194 46214 33206 46266
rect 33258 46214 42950 46266
rect 43002 46214 43014 46266
rect 43066 46214 43078 46266
rect 43130 46214 43142 46266
rect 43194 46214 43206 46266
rect 43258 46214 49864 46266
rect 1104 46192 49864 46214
rect 11054 46112 11060 46164
rect 11112 46112 11118 46164
rect 19242 46112 19248 46164
rect 19300 46152 19306 46164
rect 19429 46155 19487 46161
rect 19429 46152 19441 46155
rect 19300 46124 19441 46152
rect 19300 46112 19306 46124
rect 19429 46121 19441 46124
rect 19475 46121 19487 46155
rect 19429 46115 19487 46121
rect 21726 46112 21732 46164
rect 21784 46152 21790 46164
rect 21986 46155 22044 46161
rect 21986 46152 21998 46155
rect 21784 46124 21998 46152
rect 21784 46112 21790 46124
rect 21986 46121 21998 46124
rect 22032 46152 22044 46155
rect 22032 46124 23428 46152
rect 22032 46121 22044 46124
rect 21986 46115 22044 46121
rect 1302 45976 1308 46028
rect 1360 46016 1366 46028
rect 2041 46019 2099 46025
rect 2041 46016 2053 46019
rect 1360 45988 2053 46016
rect 1360 45976 1366 45988
rect 2041 45985 2053 45988
rect 2087 45985 2099 46019
rect 2041 45979 2099 45985
rect 20990 45976 20996 46028
rect 21048 45976 21054 46028
rect 21177 46019 21235 46025
rect 21177 45985 21189 46019
rect 21223 46016 21235 46019
rect 21358 46016 21364 46028
rect 21223 45988 21364 46016
rect 21223 45985 21235 45988
rect 21177 45979 21235 45985
rect 21358 45976 21364 45988
rect 21416 45976 21422 46028
rect 21729 46019 21787 46025
rect 21729 45985 21741 46019
rect 21775 46016 21787 46019
rect 22094 46016 22100 46028
rect 21775 45988 22100 46016
rect 21775 45985 21787 45988
rect 21729 45979 21787 45985
rect 1765 45951 1823 45957
rect 1765 45917 1777 45951
rect 1811 45948 1823 45951
rect 12250 45948 12256 45960
rect 1811 45920 12256 45948
rect 1811 45917 1823 45920
rect 1765 45911 1823 45917
rect 12250 45908 12256 45920
rect 12308 45908 12314 45960
rect 19610 45908 19616 45960
rect 19668 45908 19674 45960
rect 19702 45908 19708 45960
rect 19760 45948 19766 45960
rect 21744 45948 21772 45979
rect 22094 45976 22100 45988
rect 22152 46016 22158 46028
rect 23290 46016 23296 46028
rect 22152 45988 23296 46016
rect 22152 45976 22158 45988
rect 23290 45976 23296 45988
rect 23348 45976 23354 46028
rect 23400 46016 23428 46124
rect 23474 46112 23480 46164
rect 23532 46112 23538 46164
rect 25038 46112 25044 46164
rect 25096 46112 25102 46164
rect 25406 46112 25412 46164
rect 25464 46152 25470 46164
rect 29914 46152 29920 46164
rect 25464 46124 29920 46152
rect 25464 46112 25470 46124
rect 29914 46112 29920 46124
rect 29972 46112 29978 46164
rect 30009 46155 30067 46161
rect 30009 46121 30021 46155
rect 30055 46152 30067 46155
rect 30650 46152 30656 46164
rect 30055 46124 30656 46152
rect 30055 46121 30067 46124
rect 30009 46115 30067 46121
rect 30650 46112 30656 46124
rect 30708 46112 30714 46164
rect 32766 46152 32772 46164
rect 30760 46124 32772 46152
rect 24302 46044 24308 46096
rect 24360 46084 24366 46096
rect 26237 46087 26295 46093
rect 26237 46084 26249 46087
rect 24360 46056 26249 46084
rect 24360 46044 24366 46056
rect 26237 46053 26249 46056
rect 26283 46053 26295 46087
rect 26970 46084 26976 46096
rect 26237 46047 26295 46053
rect 26344 46056 26976 46084
rect 25685 46019 25743 46025
rect 25685 46016 25697 46019
rect 23400 45988 25697 46016
rect 25685 45985 25697 45988
rect 25731 46016 25743 46019
rect 26344 46016 26372 46056
rect 26970 46044 26976 46056
rect 27028 46044 27034 46096
rect 28994 46044 29000 46096
rect 29052 46084 29058 46096
rect 30760 46084 30788 46124
rect 32766 46112 32772 46124
rect 32824 46112 32830 46164
rect 35434 46112 35440 46164
rect 35492 46152 35498 46164
rect 35492 46124 38148 46152
rect 35492 46112 35498 46124
rect 29052 46056 30788 46084
rect 29052 46044 29058 46056
rect 31018 46044 31024 46096
rect 31076 46044 31082 46096
rect 33428 46056 35296 46084
rect 25731 45988 26372 46016
rect 25731 45985 25743 45988
rect 25685 45979 25743 45985
rect 26694 45976 26700 46028
rect 26752 45976 26758 46028
rect 26786 45976 26792 46028
rect 26844 45976 26850 46028
rect 27433 46019 27491 46025
rect 27433 45985 27445 46019
rect 27479 46016 27491 46019
rect 29454 46016 29460 46028
rect 27479 45988 29460 46016
rect 27479 45985 27491 45988
rect 27433 45979 27491 45985
rect 29454 45976 29460 45988
rect 29512 46016 29518 46028
rect 30006 46016 30012 46028
rect 29512 45988 30012 46016
rect 29512 45976 29518 45988
rect 30006 45976 30012 45988
rect 30064 45976 30070 46028
rect 30190 45976 30196 46028
rect 30248 46016 30254 46028
rect 30561 46019 30619 46025
rect 30561 46016 30573 46019
rect 30248 45988 30573 46016
rect 30248 45976 30254 45988
rect 30561 45985 30573 45988
rect 30607 45985 30619 46019
rect 30561 45979 30619 45985
rect 30834 45976 30840 46028
rect 30892 46016 30898 46028
rect 31481 46019 31539 46025
rect 31481 46016 31493 46019
rect 30892 45988 31493 46016
rect 30892 45976 30898 45988
rect 31481 45985 31493 45988
rect 31527 45985 31539 46019
rect 31481 45979 31539 45985
rect 31570 45976 31576 46028
rect 31628 45976 31634 46028
rect 33428 46025 33456 46056
rect 33413 46019 33471 46025
rect 33413 45985 33425 46019
rect 33459 45985 33471 46019
rect 33413 45979 33471 45985
rect 34514 45976 34520 46028
rect 34572 46016 34578 46028
rect 34882 46016 34888 46028
rect 34572 45988 34888 46016
rect 34572 45976 34578 45988
rect 34882 45976 34888 45988
rect 34940 46016 34946 46028
rect 35161 46019 35219 46025
rect 35161 46016 35173 46019
rect 34940 45988 35173 46016
rect 34940 45976 34946 45988
rect 35161 45985 35173 45988
rect 35207 45985 35219 46019
rect 35268 46016 35296 46056
rect 35434 46016 35440 46028
rect 35268 45988 35440 46016
rect 35161 45979 35219 45985
rect 35434 45976 35440 45988
rect 35492 46016 35498 46028
rect 36814 46016 36820 46028
rect 35492 45988 36820 46016
rect 35492 45976 35498 45988
rect 36814 45976 36820 45988
rect 36872 45976 36878 46028
rect 38013 46019 38071 46025
rect 38013 45985 38025 46019
rect 38059 45985 38071 46019
rect 38013 45979 38071 45985
rect 19760 45920 21772 45948
rect 25409 45951 25467 45957
rect 19760 45908 19766 45920
rect 25409 45917 25421 45951
rect 25455 45948 25467 45951
rect 25498 45948 25504 45960
rect 25455 45920 25504 45948
rect 25455 45917 25467 45920
rect 25409 45911 25467 45917
rect 25498 45908 25504 45920
rect 25556 45908 25562 45960
rect 25958 45908 25964 45960
rect 26016 45948 26022 45960
rect 26605 45951 26663 45957
rect 26605 45948 26617 45951
rect 26016 45920 26617 45948
rect 26016 45908 26022 45920
rect 26605 45917 26617 45920
rect 26651 45948 26663 45951
rect 27338 45948 27344 45960
rect 26651 45920 27344 45948
rect 26651 45917 26663 45920
rect 26605 45911 26663 45917
rect 27338 45908 27344 45920
rect 27396 45908 27402 45960
rect 29178 45908 29184 45960
rect 29236 45908 29242 45960
rect 29914 45908 29920 45960
rect 29972 45948 29978 45960
rect 30469 45951 30527 45957
rect 30469 45948 30481 45951
rect 29972 45920 30481 45948
rect 29972 45908 29978 45920
rect 30469 45917 30481 45920
rect 30515 45917 30527 45951
rect 30469 45911 30527 45917
rect 31389 45951 31447 45957
rect 31389 45917 31401 45951
rect 31435 45948 31447 45951
rect 31662 45948 31668 45960
rect 31435 45920 31668 45948
rect 31435 45917 31447 45920
rect 31389 45911 31447 45917
rect 31662 45908 31668 45920
rect 31720 45908 31726 45960
rect 32309 45951 32367 45957
rect 32309 45917 32321 45951
rect 32355 45948 32367 45951
rect 32490 45948 32496 45960
rect 32355 45920 32496 45948
rect 32355 45917 32367 45920
rect 32309 45911 32367 45917
rect 32490 45908 32496 45920
rect 32548 45948 32554 45960
rect 33137 45951 33195 45957
rect 33137 45948 33149 45951
rect 32548 45920 33149 45948
rect 32548 45908 32554 45920
rect 33137 45917 33149 45920
rect 33183 45948 33195 45951
rect 33183 45920 33548 45948
rect 33183 45917 33195 45920
rect 33137 45911 33195 45917
rect 10965 45883 11023 45889
rect 10965 45849 10977 45883
rect 11011 45880 11023 45883
rect 12526 45880 12532 45892
rect 11011 45852 12532 45880
rect 11011 45849 11023 45852
rect 10965 45843 11023 45849
rect 12526 45840 12532 45852
rect 12584 45880 12590 45892
rect 13630 45880 13636 45892
rect 12584 45852 13636 45880
rect 12584 45840 12590 45852
rect 13630 45840 13636 45852
rect 13688 45840 13694 45892
rect 20901 45883 20959 45889
rect 20901 45849 20913 45883
rect 20947 45880 20959 45883
rect 23842 45880 23848 45892
rect 20947 45852 21496 45880
rect 23230 45852 23848 45880
rect 20947 45849 20959 45852
rect 20901 45843 20959 45849
rect 18598 45772 18604 45824
rect 18656 45812 18662 45824
rect 20533 45815 20591 45821
rect 20533 45812 20545 45815
rect 18656 45784 20545 45812
rect 18656 45772 18662 45784
rect 20533 45781 20545 45784
rect 20579 45781 20591 45815
rect 21468 45812 21496 45852
rect 23842 45840 23848 45852
rect 23900 45840 23906 45892
rect 27706 45840 27712 45892
rect 27764 45840 27770 45892
rect 29196 45880 29224 45908
rect 28934 45852 29224 45880
rect 30377 45883 30435 45889
rect 30377 45849 30389 45883
rect 30423 45880 30435 45883
rect 31294 45880 31300 45892
rect 30423 45852 31300 45880
rect 30423 45849 30435 45852
rect 30377 45843 30435 45849
rect 31294 45840 31300 45852
rect 31352 45840 31358 45892
rect 32950 45880 32956 45892
rect 31588 45852 32956 45880
rect 23382 45812 23388 45824
rect 21468 45784 23388 45812
rect 20533 45775 20591 45781
rect 23382 45772 23388 45784
rect 23440 45772 23446 45824
rect 23474 45772 23480 45824
rect 23532 45812 23538 45824
rect 25501 45815 25559 45821
rect 25501 45812 25513 45815
rect 23532 45784 25513 45812
rect 23532 45772 23538 45784
rect 25501 45781 25513 45784
rect 25547 45812 25559 45815
rect 26694 45812 26700 45824
rect 25547 45784 26700 45812
rect 25547 45781 25559 45784
rect 25501 45775 25559 45781
rect 26694 45772 26700 45784
rect 26752 45772 26758 45824
rect 26786 45772 26792 45824
rect 26844 45812 26850 45824
rect 29181 45815 29239 45821
rect 29181 45812 29193 45815
rect 26844 45784 29193 45812
rect 26844 45772 26850 45784
rect 29181 45781 29193 45784
rect 29227 45781 29239 45815
rect 29181 45775 29239 45781
rect 29270 45772 29276 45824
rect 29328 45812 29334 45824
rect 31588 45812 31616 45852
rect 32950 45840 32956 45852
rect 33008 45840 33014 45892
rect 33226 45840 33232 45892
rect 33284 45840 33290 45892
rect 33520 45880 33548 45920
rect 34146 45908 34152 45960
rect 34204 45908 34210 45960
rect 36538 45908 36544 45960
rect 36596 45908 36602 45960
rect 37826 45908 37832 45960
rect 37884 45908 37890 45960
rect 34238 45880 34244 45892
rect 33520 45852 34244 45880
rect 34238 45840 34244 45852
rect 34296 45840 34302 45892
rect 35342 45840 35348 45892
rect 35400 45880 35406 45892
rect 35437 45883 35495 45889
rect 35437 45880 35449 45883
rect 35400 45852 35449 45880
rect 35400 45840 35406 45852
rect 35437 45849 35449 45852
rect 35483 45849 35495 45883
rect 38028 45880 38056 45979
rect 35437 45843 35495 45849
rect 37200 45852 38056 45880
rect 37200 45824 37228 45852
rect 29328 45784 31616 45812
rect 32769 45815 32827 45821
rect 29328 45772 29334 45784
rect 32769 45781 32781 45815
rect 32815 45812 32827 45815
rect 35526 45812 35532 45824
rect 32815 45784 35532 45812
rect 32815 45781 32827 45784
rect 32769 45775 32827 45781
rect 35526 45772 35532 45784
rect 35584 45772 35590 45824
rect 36909 45815 36967 45821
rect 36909 45781 36921 45815
rect 36955 45812 36967 45815
rect 37182 45812 37188 45824
rect 36955 45784 37188 45812
rect 36955 45781 36967 45784
rect 36909 45775 36967 45781
rect 37182 45772 37188 45784
rect 37240 45772 37246 45824
rect 37461 45815 37519 45821
rect 37461 45781 37473 45815
rect 37507 45812 37519 45815
rect 37734 45812 37740 45824
rect 37507 45784 37740 45812
rect 37507 45781 37519 45784
rect 37461 45775 37519 45781
rect 37734 45772 37740 45784
rect 37792 45772 37798 45824
rect 37921 45815 37979 45821
rect 37921 45781 37933 45815
rect 37967 45812 37979 45815
rect 38120 45812 38148 46124
rect 49050 45908 49056 45960
rect 49108 45908 49114 45960
rect 39114 45812 39120 45824
rect 37967 45784 39120 45812
rect 37967 45781 37979 45784
rect 37921 45775 37979 45781
rect 39114 45772 39120 45784
rect 39172 45772 39178 45824
rect 48590 45772 48596 45824
rect 48648 45812 48654 45824
rect 49237 45815 49295 45821
rect 49237 45812 49249 45815
rect 48648 45784 49249 45812
rect 48648 45772 48654 45784
rect 49237 45781 49249 45784
rect 49283 45781 49295 45815
rect 49237 45775 49295 45781
rect 1104 45722 49864 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 27950 45722
rect 28002 45670 28014 45722
rect 28066 45670 28078 45722
rect 28130 45670 28142 45722
rect 28194 45670 28206 45722
rect 28258 45670 37950 45722
rect 38002 45670 38014 45722
rect 38066 45670 38078 45722
rect 38130 45670 38142 45722
rect 38194 45670 38206 45722
rect 38258 45670 47950 45722
rect 48002 45670 48014 45722
rect 48066 45670 48078 45722
rect 48130 45670 48142 45722
rect 48194 45670 48206 45722
rect 48258 45670 49864 45722
rect 1104 45648 49864 45670
rect 20806 45608 20812 45620
rect 20364 45580 20812 45608
rect 7558 45500 7564 45552
rect 7616 45540 7622 45552
rect 7653 45543 7711 45549
rect 7653 45540 7665 45543
rect 7616 45512 7665 45540
rect 7616 45500 7622 45512
rect 7653 45509 7665 45512
rect 7699 45509 7711 45543
rect 20364 45540 20392 45580
rect 20806 45568 20812 45580
rect 20864 45568 20870 45620
rect 22741 45611 22799 45617
rect 22741 45577 22753 45611
rect 22787 45608 22799 45611
rect 25133 45611 25191 45617
rect 22787 45580 24348 45608
rect 22787 45577 22799 45580
rect 22741 45571 22799 45577
rect 7653 45503 7711 45509
rect 18248 45512 20392 45540
rect 22649 45543 22707 45549
rect 7469 45475 7527 45481
rect 7469 45441 7481 45475
rect 7515 45441 7527 45475
rect 7469 45435 7527 45441
rect 12161 45475 12219 45481
rect 12161 45441 12173 45475
rect 12207 45472 12219 45475
rect 12802 45472 12808 45484
rect 12207 45444 12808 45472
rect 12207 45441 12219 45444
rect 12161 45435 12219 45441
rect 7484 45404 7512 45435
rect 12802 45432 12808 45444
rect 12860 45432 12866 45484
rect 13357 45475 13415 45481
rect 13357 45441 13369 45475
rect 13403 45472 13415 45475
rect 16574 45472 16580 45484
rect 13403 45444 16580 45472
rect 13403 45441 13415 45444
rect 13357 45435 13415 45441
rect 16574 45432 16580 45444
rect 16632 45432 16638 45484
rect 18248 45481 18276 45512
rect 22649 45509 22661 45543
rect 22695 45540 22707 45543
rect 23750 45540 23756 45552
rect 22695 45512 23756 45540
rect 22695 45509 22707 45512
rect 22649 45503 22707 45509
rect 23750 45500 23756 45512
rect 23808 45500 23814 45552
rect 23934 45500 23940 45552
rect 23992 45500 23998 45552
rect 24320 45540 24348 45580
rect 25133 45577 25145 45611
rect 25179 45608 25191 45611
rect 25406 45608 25412 45620
rect 25179 45580 25412 45608
rect 25179 45577 25191 45580
rect 25133 45571 25191 45577
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 25869 45611 25927 45617
rect 25869 45577 25881 45611
rect 25915 45577 25927 45611
rect 26418 45608 26424 45620
rect 25869 45571 25927 45577
rect 25976 45580 26424 45608
rect 25884 45540 25912 45571
rect 24320 45512 25912 45540
rect 18233 45475 18291 45481
rect 18233 45441 18245 45475
rect 18279 45441 18291 45475
rect 18233 45435 18291 45441
rect 19702 45432 19708 45484
rect 19760 45432 19766 45484
rect 21082 45432 21088 45484
rect 21140 45432 21146 45484
rect 23842 45432 23848 45484
rect 23900 45432 23906 45484
rect 25038 45432 25044 45484
rect 25096 45432 25102 45484
rect 13814 45404 13820 45416
rect 7484 45376 13820 45404
rect 13814 45364 13820 45376
rect 13872 45364 13878 45416
rect 19978 45364 19984 45416
rect 20036 45364 20042 45416
rect 20714 45364 20720 45416
rect 20772 45404 20778 45416
rect 20772 45376 22094 45404
rect 20772 45364 20778 45376
rect 9950 45296 9956 45348
rect 10008 45336 10014 45348
rect 11977 45339 12035 45345
rect 11977 45336 11989 45339
rect 10008 45308 11989 45336
rect 10008 45296 10014 45308
rect 11977 45305 11989 45308
rect 12023 45305 12035 45339
rect 11977 45299 12035 45305
rect 18049 45339 18107 45345
rect 18049 45305 18061 45339
rect 18095 45336 18107 45339
rect 18322 45336 18328 45348
rect 18095 45308 18328 45336
rect 18095 45305 18107 45308
rect 18049 45299 18107 45305
rect 18322 45296 18328 45308
rect 18380 45296 18386 45348
rect 20990 45296 20996 45348
rect 21048 45336 21054 45348
rect 21453 45339 21511 45345
rect 21453 45336 21465 45339
rect 21048 45308 21465 45336
rect 21048 45296 21054 45308
rect 21453 45305 21465 45308
rect 21499 45336 21511 45339
rect 21542 45336 21548 45348
rect 21499 45308 21548 45336
rect 21499 45305 21511 45308
rect 21453 45299 21511 45305
rect 21542 45296 21548 45308
rect 21600 45296 21606 45348
rect 22066 45336 22094 45376
rect 22830 45364 22836 45416
rect 22888 45364 22894 45416
rect 24026 45364 24032 45416
rect 24084 45364 24090 45416
rect 24118 45364 24124 45416
rect 24176 45404 24182 45416
rect 25317 45407 25375 45413
rect 25317 45404 25329 45407
rect 24176 45376 25329 45404
rect 24176 45364 24182 45376
rect 25317 45373 25329 45376
rect 25363 45404 25375 45407
rect 25976 45404 26004 45580
rect 26418 45568 26424 45580
rect 26476 45568 26482 45620
rect 26694 45568 26700 45620
rect 26752 45608 26758 45620
rect 28166 45608 28172 45620
rect 26752 45580 28172 45608
rect 26752 45568 26758 45580
rect 28166 45568 28172 45580
rect 28224 45568 28230 45620
rect 28258 45568 28264 45620
rect 28316 45608 28322 45620
rect 28626 45608 28632 45620
rect 28316 45580 28632 45608
rect 28316 45568 28322 45580
rect 28626 45568 28632 45580
rect 28684 45568 28690 45620
rect 32306 45568 32312 45620
rect 32364 45608 32370 45620
rect 32953 45611 33011 45617
rect 32953 45608 32965 45611
rect 32364 45580 32965 45608
rect 32364 45568 32370 45580
rect 32953 45577 32965 45580
rect 32999 45577 33011 45611
rect 32953 45571 33011 45577
rect 33410 45568 33416 45620
rect 33468 45608 33474 45620
rect 33781 45611 33839 45617
rect 33781 45608 33793 45611
rect 33468 45580 33793 45608
rect 33468 45568 33474 45580
rect 33781 45577 33793 45580
rect 33827 45577 33839 45611
rect 33781 45571 33839 45577
rect 34146 45568 34152 45620
rect 34204 45568 34210 45620
rect 34238 45568 34244 45620
rect 34296 45608 34302 45620
rect 38654 45608 38660 45620
rect 34296 45580 38660 45608
rect 34296 45568 34302 45580
rect 38654 45568 38660 45580
rect 38712 45568 38718 45620
rect 26326 45500 26332 45552
rect 26384 45500 26390 45552
rect 27525 45543 27583 45549
rect 27525 45509 27537 45543
rect 27571 45540 27583 45543
rect 27706 45540 27712 45552
rect 27571 45512 27712 45540
rect 27571 45509 27583 45512
rect 27525 45503 27583 45509
rect 27706 45500 27712 45512
rect 27764 45540 27770 45552
rect 28442 45540 28448 45552
rect 27764 45512 28448 45540
rect 27764 45500 27770 45512
rect 28442 45500 28448 45512
rect 28500 45500 28506 45552
rect 29638 45540 29644 45552
rect 28552 45512 29644 45540
rect 26237 45475 26295 45481
rect 26237 45441 26249 45475
rect 26283 45441 26295 45475
rect 26237 45435 26295 45441
rect 27617 45475 27675 45481
rect 27617 45441 27629 45475
rect 27663 45472 27675 45475
rect 28552 45472 28580 45512
rect 29638 45500 29644 45512
rect 29696 45500 29702 45552
rect 30101 45543 30159 45549
rect 30101 45509 30113 45543
rect 30147 45540 30159 45543
rect 32490 45540 32496 45552
rect 30147 45512 32496 45540
rect 30147 45509 30159 45512
rect 30101 45503 30159 45509
rect 32490 45500 32496 45512
rect 32548 45500 32554 45552
rect 32858 45500 32864 45552
rect 32916 45540 32922 45552
rect 33045 45543 33103 45549
rect 33045 45540 33057 45543
rect 32916 45512 33057 45540
rect 32916 45500 32922 45512
rect 33045 45509 33057 45512
rect 33091 45509 33103 45543
rect 33045 45503 33103 45509
rect 33226 45500 33232 45552
rect 33284 45540 33290 45552
rect 34330 45540 34336 45552
rect 33284 45512 34336 45540
rect 33284 45500 33290 45512
rect 34330 45500 34336 45512
rect 34388 45540 34394 45552
rect 39669 45543 39727 45549
rect 34388 45512 35756 45540
rect 34388 45500 34394 45512
rect 27663 45444 28580 45472
rect 27663 45441 27675 45444
rect 27617 45435 27675 45441
rect 25363 45376 26004 45404
rect 25363 45373 25375 45376
rect 25317 45367 25375 45373
rect 23477 45339 23535 45345
rect 23477 45336 23489 45339
rect 22066 45308 23489 45336
rect 23477 45305 23489 45308
rect 23523 45305 23535 45339
rect 26252 45336 26280 45435
rect 28626 45432 28632 45484
rect 28684 45472 28690 45484
rect 28721 45475 28779 45481
rect 28721 45472 28733 45475
rect 28684 45444 28733 45472
rect 28684 45432 28690 45444
rect 28721 45441 28733 45444
rect 28767 45441 28779 45475
rect 28721 45435 28779 45441
rect 28994 45432 29000 45484
rect 29052 45472 29058 45484
rect 29730 45472 29736 45484
rect 29052 45444 29736 45472
rect 29052 45432 29058 45444
rect 29730 45432 29736 45444
rect 29788 45472 29794 45484
rect 30558 45472 30564 45484
rect 29788 45444 30564 45472
rect 29788 45432 29794 45444
rect 30558 45432 30564 45444
rect 30616 45432 30622 45484
rect 31389 45475 31447 45481
rect 31389 45441 31401 45475
rect 31435 45472 31447 45475
rect 34054 45472 34060 45484
rect 31435 45444 34060 45472
rect 31435 45441 31447 45444
rect 31389 45435 31447 45441
rect 34054 45432 34060 45444
rect 34112 45432 34118 45484
rect 35728 45481 35756 45512
rect 39669 45509 39681 45543
rect 39715 45540 39727 45543
rect 39758 45540 39764 45552
rect 39715 45512 39764 45540
rect 39715 45509 39727 45512
rect 39669 45503 39727 45509
rect 39758 45500 39764 45512
rect 39816 45500 39822 45552
rect 35713 45475 35771 45481
rect 35713 45441 35725 45475
rect 35759 45472 35771 45475
rect 36541 45475 36599 45481
rect 36541 45472 36553 45475
rect 35759 45444 36553 45472
rect 35759 45441 35771 45444
rect 35713 45435 35771 45441
rect 36541 45441 36553 45444
rect 36587 45472 36599 45475
rect 37829 45475 37887 45481
rect 36587 45444 36860 45472
rect 36587 45441 36599 45444
rect 36541 45435 36599 45441
rect 26513 45407 26571 45413
rect 26513 45373 26525 45407
rect 26559 45404 26571 45407
rect 26602 45404 26608 45416
rect 26559 45376 26608 45404
rect 26559 45373 26571 45376
rect 26513 45367 26571 45373
rect 26602 45364 26608 45376
rect 26660 45364 26666 45416
rect 26970 45364 26976 45416
rect 27028 45404 27034 45416
rect 27709 45407 27767 45413
rect 27709 45404 27721 45407
rect 27028 45376 27721 45404
rect 27028 45364 27034 45376
rect 27709 45373 27721 45376
rect 27755 45373 27767 45407
rect 27709 45367 27767 45373
rect 28813 45407 28871 45413
rect 28813 45373 28825 45407
rect 28859 45373 28871 45407
rect 28813 45367 28871 45373
rect 28905 45407 28963 45413
rect 28905 45373 28917 45407
rect 28951 45373 28963 45407
rect 28905 45367 28963 45373
rect 28353 45339 28411 45345
rect 28353 45336 28365 45339
rect 26252 45308 28365 45336
rect 23477 45299 23535 45305
rect 28353 45305 28365 45308
rect 28399 45305 28411 45339
rect 28353 45299 28411 45305
rect 28718 45296 28724 45348
rect 28776 45336 28782 45348
rect 28828 45336 28856 45367
rect 28776 45308 28856 45336
rect 28920 45336 28948 45367
rect 29270 45364 29276 45416
rect 29328 45404 29334 45416
rect 30193 45407 30251 45413
rect 30193 45404 30205 45407
rect 29328 45376 30205 45404
rect 29328 45364 29334 45376
rect 30193 45373 30205 45376
rect 30239 45373 30251 45407
rect 30193 45367 30251 45373
rect 30282 45364 30288 45416
rect 30340 45364 30346 45416
rect 30374 45364 30380 45416
rect 30432 45404 30438 45416
rect 31481 45407 31539 45413
rect 31481 45404 31493 45407
rect 30432 45376 31493 45404
rect 30432 45364 30438 45376
rect 31481 45373 31493 45376
rect 31527 45373 31539 45407
rect 31481 45367 31539 45373
rect 31665 45407 31723 45413
rect 31665 45373 31677 45407
rect 31711 45404 31723 45407
rect 32030 45404 32036 45416
rect 31711 45376 32036 45404
rect 31711 45373 31723 45376
rect 31665 45367 31723 45373
rect 32030 45364 32036 45376
rect 32088 45364 32094 45416
rect 32766 45364 32772 45416
rect 32824 45404 32830 45416
rect 33137 45407 33195 45413
rect 33137 45404 33149 45407
rect 32824 45376 33149 45404
rect 32824 45364 32830 45376
rect 33137 45373 33149 45376
rect 33183 45373 33195 45407
rect 33137 45367 33195 45373
rect 33502 45364 33508 45416
rect 33560 45404 33566 45416
rect 34241 45407 34299 45413
rect 34241 45404 34253 45407
rect 33560 45376 34253 45404
rect 33560 45364 33566 45376
rect 34241 45373 34253 45376
rect 34287 45373 34299 45407
rect 34241 45367 34299 45373
rect 34425 45407 34483 45413
rect 34425 45373 34437 45407
rect 34471 45404 34483 45407
rect 34790 45404 34796 45416
rect 34471 45376 34796 45404
rect 34471 45373 34483 45376
rect 34425 45367 34483 45373
rect 34790 45364 34796 45376
rect 34848 45364 34854 45416
rect 36446 45364 36452 45416
rect 36504 45404 36510 45416
rect 36633 45407 36691 45413
rect 36633 45404 36645 45407
rect 36504 45376 36645 45404
rect 36504 45364 36510 45376
rect 36633 45373 36645 45376
rect 36679 45373 36691 45407
rect 36633 45367 36691 45373
rect 36725 45407 36783 45413
rect 36725 45373 36737 45407
rect 36771 45373 36783 45407
rect 36725 45367 36783 45373
rect 30098 45336 30104 45348
rect 28920 45308 30104 45336
rect 28776 45296 28782 45308
rect 30098 45296 30104 45308
rect 30156 45296 30162 45348
rect 31021 45339 31079 45345
rect 31021 45305 31033 45339
rect 31067 45336 31079 45339
rect 31110 45336 31116 45348
rect 31067 45308 31116 45336
rect 31067 45305 31079 45308
rect 31021 45299 31079 45305
rect 31110 45296 31116 45308
rect 31168 45296 31174 45348
rect 31294 45296 31300 45348
rect 31352 45336 31358 45348
rect 33226 45336 33232 45348
rect 31352 45308 33232 45336
rect 31352 45296 31358 45308
rect 33226 45296 33232 45308
rect 33284 45296 33290 45348
rect 34146 45296 34152 45348
rect 34204 45336 34210 45348
rect 36740 45336 36768 45367
rect 34204 45308 36768 45336
rect 36832 45336 36860 45444
rect 37829 45441 37841 45475
rect 37875 45472 37887 45475
rect 39577 45475 39635 45481
rect 37875 45444 39252 45472
rect 37875 45441 37887 45444
rect 37829 45435 37887 45441
rect 37458 45364 37464 45416
rect 37516 45404 37522 45416
rect 37921 45407 37979 45413
rect 37921 45404 37933 45407
rect 37516 45376 37933 45404
rect 37516 45364 37522 45376
rect 37921 45373 37933 45376
rect 37967 45373 37979 45407
rect 37921 45367 37979 45373
rect 38010 45364 38016 45416
rect 38068 45364 38074 45416
rect 39224 45345 39252 45444
rect 39577 45441 39589 45475
rect 39623 45472 39635 45475
rect 42794 45472 42800 45484
rect 39623 45444 42800 45472
rect 39623 45441 39635 45444
rect 39577 45435 39635 45441
rect 42794 45432 42800 45444
rect 42852 45432 42858 45484
rect 39482 45364 39488 45416
rect 39540 45404 39546 45416
rect 39761 45407 39819 45413
rect 39761 45404 39773 45407
rect 39540 45376 39773 45404
rect 39540 45364 39546 45376
rect 39761 45373 39773 45376
rect 39807 45373 39819 45407
rect 39761 45367 39819 45373
rect 39209 45339 39267 45345
rect 36832 45308 37596 45336
rect 34204 45296 34210 45308
rect 6822 45228 6828 45280
rect 6880 45268 6886 45280
rect 13173 45271 13231 45277
rect 13173 45268 13185 45271
rect 6880 45240 13185 45268
rect 6880 45228 6886 45240
rect 13173 45237 13185 45240
rect 13219 45237 13231 45271
rect 13173 45231 13231 45237
rect 18877 45271 18935 45277
rect 18877 45237 18889 45271
rect 18923 45268 18935 45271
rect 20438 45268 20444 45280
rect 18923 45240 20444 45268
rect 18923 45237 18935 45240
rect 18877 45231 18935 45237
rect 20438 45228 20444 45240
rect 20496 45228 20502 45280
rect 22186 45228 22192 45280
rect 22244 45268 22250 45280
rect 22281 45271 22339 45277
rect 22281 45268 22293 45271
rect 22244 45240 22293 45268
rect 22244 45228 22250 45240
rect 22281 45237 22293 45240
rect 22327 45237 22339 45271
rect 22281 45231 22339 45237
rect 23382 45228 23388 45280
rect 23440 45268 23446 45280
rect 24673 45271 24731 45277
rect 24673 45268 24685 45271
rect 23440 45240 24685 45268
rect 23440 45228 23446 45240
rect 24673 45237 24685 45240
rect 24719 45237 24731 45271
rect 24673 45231 24731 45237
rect 24762 45228 24768 45280
rect 24820 45268 24826 45280
rect 27157 45271 27215 45277
rect 27157 45268 27169 45271
rect 24820 45240 27169 45268
rect 24820 45228 24826 45240
rect 27157 45237 27169 45240
rect 27203 45237 27215 45271
rect 27157 45231 27215 45237
rect 28166 45228 28172 45280
rect 28224 45268 28230 45280
rect 29270 45268 29276 45280
rect 28224 45240 29276 45268
rect 28224 45228 28230 45240
rect 29270 45228 29276 45240
rect 29328 45228 29334 45280
rect 29730 45228 29736 45280
rect 29788 45228 29794 45280
rect 32585 45271 32643 45277
rect 32585 45237 32597 45271
rect 32631 45268 32643 45271
rect 35250 45268 35256 45280
rect 32631 45240 35256 45268
rect 32631 45237 32643 45240
rect 32585 45231 32643 45237
rect 35250 45228 35256 45240
rect 35308 45228 35314 45280
rect 36170 45228 36176 45280
rect 36228 45228 36234 45280
rect 37366 45228 37372 45280
rect 37424 45268 37430 45280
rect 37461 45271 37519 45277
rect 37461 45268 37473 45271
rect 37424 45240 37473 45268
rect 37424 45228 37430 45240
rect 37461 45237 37473 45240
rect 37507 45237 37519 45271
rect 37568 45268 37596 45308
rect 39209 45305 39221 45339
rect 39255 45305 39267 45339
rect 39209 45299 39267 45305
rect 46198 45268 46204 45280
rect 37568 45240 46204 45268
rect 37461 45231 37519 45237
rect 46198 45228 46204 45240
rect 46256 45228 46262 45280
rect 1104 45178 49864 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 32950 45178
rect 33002 45126 33014 45178
rect 33066 45126 33078 45178
rect 33130 45126 33142 45178
rect 33194 45126 33206 45178
rect 33258 45126 42950 45178
rect 43002 45126 43014 45178
rect 43066 45126 43078 45178
rect 43130 45126 43142 45178
rect 43194 45126 43206 45178
rect 43258 45126 49864 45178
rect 1104 45104 49864 45126
rect 5626 45024 5632 45076
rect 5684 45064 5690 45076
rect 7285 45067 7343 45073
rect 7285 45064 7297 45067
rect 5684 45036 7297 45064
rect 5684 45024 5690 45036
rect 7285 45033 7297 45036
rect 7331 45033 7343 45067
rect 7285 45027 7343 45033
rect 11606 45024 11612 45076
rect 11664 45064 11670 45076
rect 12713 45067 12771 45073
rect 12713 45064 12725 45067
rect 11664 45036 12725 45064
rect 11664 45024 11670 45036
rect 12713 45033 12725 45036
rect 12759 45033 12771 45067
rect 12713 45027 12771 45033
rect 18141 45067 18199 45073
rect 18141 45033 18153 45067
rect 18187 45064 18199 45067
rect 19794 45064 19800 45076
rect 18187 45036 19800 45064
rect 18187 45033 18199 45036
rect 18141 45027 18199 45033
rect 19794 45024 19800 45036
rect 19852 45024 19858 45076
rect 21818 45064 21824 45076
rect 19904 45036 21824 45064
rect 18690 44956 18696 45008
rect 18748 44996 18754 45008
rect 19904 44996 19932 45036
rect 21818 45024 21824 45036
rect 21876 45024 21882 45076
rect 26789 45067 26847 45073
rect 26789 45064 26801 45067
rect 23768 45036 26801 45064
rect 18748 44968 19932 44996
rect 18748 44956 18754 44968
rect 1302 44888 1308 44940
rect 1360 44928 1366 44940
rect 2041 44931 2099 44937
rect 2041 44928 2053 44931
rect 1360 44900 2053 44928
rect 1360 44888 1366 44900
rect 2041 44897 2053 44900
rect 2087 44897 2099 44931
rect 2041 44891 2099 44897
rect 18785 44931 18843 44937
rect 18785 44897 18797 44931
rect 18831 44928 18843 44931
rect 19518 44928 19524 44940
rect 18831 44900 19524 44928
rect 18831 44897 18843 44900
rect 18785 44891 18843 44897
rect 19518 44888 19524 44900
rect 19576 44888 19582 44940
rect 20162 44888 20168 44940
rect 20220 44928 20226 44940
rect 23768 44937 23796 45036
rect 26789 45033 26801 45036
rect 26835 45033 26847 45067
rect 26789 45027 26847 45033
rect 27062 45024 27068 45076
rect 27120 45064 27126 45076
rect 29733 45067 29791 45073
rect 29733 45064 29745 45067
rect 27120 45036 29745 45064
rect 27120 45024 27126 45036
rect 29733 45033 29745 45036
rect 29779 45033 29791 45067
rect 29733 45027 29791 45033
rect 31202 45024 31208 45076
rect 31260 45064 31266 45076
rect 34146 45064 34152 45076
rect 31260 45036 34152 45064
rect 31260 45024 31266 45036
rect 34146 45024 34152 45036
rect 34204 45024 34210 45076
rect 34790 45024 34796 45076
rect 34848 45064 34854 45076
rect 36633 45067 36691 45073
rect 36633 45064 36645 45067
rect 34848 45036 36645 45064
rect 34848 45024 34854 45036
rect 36633 45033 36645 45036
rect 36679 45064 36691 45067
rect 38010 45064 38016 45076
rect 36679 45036 38016 45064
rect 36679 45033 36691 45036
rect 36633 45027 36691 45033
rect 38010 45024 38016 45036
rect 38068 45024 38074 45076
rect 25866 44956 25872 45008
rect 25924 44996 25930 45008
rect 26329 44999 26387 45005
rect 26329 44996 26341 44999
rect 25924 44968 26341 44996
rect 25924 44956 25930 44968
rect 26329 44965 26341 44968
rect 26375 44965 26387 44999
rect 27985 44999 28043 45005
rect 27985 44996 27997 44999
rect 26329 44959 26387 44965
rect 26436 44968 27997 44996
rect 23753 44931 23811 44937
rect 20220 44900 23060 44928
rect 20220 44888 20226 44900
rect 1765 44863 1823 44869
rect 1765 44829 1777 44863
rect 1811 44860 1823 44863
rect 11054 44860 11060 44872
rect 1811 44832 11060 44860
rect 1811 44829 1823 44832
rect 1765 44823 1823 44829
rect 11054 44820 11060 44832
rect 11112 44820 11118 44872
rect 12897 44863 12955 44869
rect 12897 44829 12909 44863
rect 12943 44860 12955 44863
rect 15010 44860 15016 44872
rect 12943 44832 15016 44860
rect 12943 44829 12955 44832
rect 12897 44823 12955 44829
rect 15010 44820 15016 44832
rect 15068 44820 15074 44872
rect 18506 44820 18512 44872
rect 18564 44820 18570 44872
rect 19702 44820 19708 44872
rect 19760 44860 19766 44872
rect 19889 44863 19947 44869
rect 19889 44860 19901 44863
rect 19760 44832 19901 44860
rect 19760 44820 19766 44832
rect 19889 44829 19901 44832
rect 19935 44829 19947 44863
rect 19889 44823 19947 44829
rect 21450 44820 21456 44872
rect 21508 44860 21514 44872
rect 22373 44863 22431 44869
rect 22373 44860 22385 44863
rect 21508 44832 22385 44860
rect 21508 44820 21514 44832
rect 22373 44829 22385 44832
rect 22419 44829 22431 44863
rect 23032 44860 23060 44900
rect 23753 44897 23765 44931
rect 23799 44897 23811 44931
rect 23753 44891 23811 44897
rect 23934 44888 23940 44940
rect 23992 44888 23998 44940
rect 25590 44888 25596 44940
rect 25648 44928 25654 44940
rect 26436 44928 26464 44968
rect 27985 44965 27997 44968
rect 28031 44965 28043 44999
rect 27985 44959 28043 44965
rect 28718 44956 28724 45008
rect 28776 44956 28782 45008
rect 29270 44956 29276 45008
rect 29328 44996 29334 45008
rect 31220 44996 31248 45024
rect 29328 44968 31248 44996
rect 29328 44956 29334 44968
rect 33594 44956 33600 45008
rect 33652 44996 33658 45008
rect 36725 44999 36783 45005
rect 33652 44968 35020 44996
rect 33652 44956 33658 44968
rect 25648 44900 26464 44928
rect 25648 44888 25654 44900
rect 27246 44888 27252 44940
rect 27304 44888 27310 44940
rect 27338 44888 27344 44940
rect 27396 44888 27402 44940
rect 28736 44928 28764 44956
rect 30377 44931 30435 44937
rect 28736 44900 28994 44928
rect 24026 44860 24032 44872
rect 23032 44832 24032 44860
rect 22373 44823 22431 44829
rect 24026 44820 24032 44832
rect 24084 44820 24090 44872
rect 24581 44863 24639 44869
rect 24581 44829 24593 44863
rect 24627 44829 24639 44863
rect 24581 44823 24639 44829
rect 27157 44863 27215 44869
rect 27157 44829 27169 44863
rect 27203 44860 27215 44863
rect 27522 44860 27528 44872
rect 27203 44832 27528 44860
rect 27203 44829 27215 44832
rect 27157 44823 27215 44829
rect 7193 44795 7251 44801
rect 7193 44761 7205 44795
rect 7239 44792 7251 44795
rect 13538 44792 13544 44804
rect 7239 44764 13544 44792
rect 7239 44761 7251 44764
rect 7193 44755 7251 44761
rect 13538 44752 13544 44764
rect 13596 44752 13602 44804
rect 16298 44752 16304 44804
rect 16356 44792 16362 44804
rect 16356 44764 19932 44792
rect 16356 44752 16362 44764
rect 19904 44736 19932 44764
rect 20162 44752 20168 44804
rect 20220 44752 20226 44804
rect 21174 44752 21180 44804
rect 21232 44752 21238 44804
rect 21818 44752 21824 44804
rect 21876 44792 21882 44804
rect 24596 44792 24624 44823
rect 27522 44820 27528 44832
rect 27580 44820 27586 44872
rect 28169 44863 28227 44869
rect 28169 44829 28181 44863
rect 28215 44860 28227 44863
rect 28442 44860 28448 44872
rect 28215 44832 28448 44860
rect 28215 44829 28227 44832
rect 28169 44823 28227 44829
rect 28442 44820 28448 44832
rect 28500 44820 28506 44872
rect 28718 44820 28724 44872
rect 28776 44860 28782 44872
rect 28813 44863 28871 44869
rect 28813 44860 28825 44863
rect 28776 44832 28825 44860
rect 28776 44820 28782 44832
rect 28813 44829 28825 44832
rect 28859 44829 28871 44863
rect 28966 44860 28994 44900
rect 30377 44897 30389 44931
rect 30423 44928 30435 44931
rect 31570 44928 31576 44940
rect 30423 44900 31576 44928
rect 30423 44897 30435 44900
rect 30377 44891 30435 44897
rect 31570 44888 31576 44900
rect 31628 44888 31634 44940
rect 31665 44931 31723 44937
rect 31665 44897 31677 44931
rect 31711 44928 31723 44931
rect 31754 44928 31760 44940
rect 31711 44900 31760 44928
rect 31711 44897 31723 44900
rect 31665 44891 31723 44897
rect 31754 44888 31760 44900
rect 31812 44928 31818 44940
rect 32674 44928 32680 44940
rect 31812 44900 32680 44928
rect 31812 44888 31818 44900
rect 32674 44888 32680 44900
rect 32732 44888 32738 44940
rect 33134 44888 33140 44940
rect 33192 44888 33198 44940
rect 33410 44888 33416 44940
rect 33468 44888 33474 44940
rect 34054 44888 34060 44940
rect 34112 44928 34118 44940
rect 34149 44931 34207 44937
rect 34149 44928 34161 44931
rect 34112 44900 34161 44928
rect 34112 44888 34118 44900
rect 34149 44897 34161 44900
rect 34195 44897 34207 44931
rect 34149 44891 34207 44897
rect 34882 44888 34888 44940
rect 34940 44888 34946 44940
rect 34992 44928 35020 44968
rect 36725 44965 36737 44999
rect 36771 44996 36783 44999
rect 37366 44996 37372 45008
rect 36771 44968 37372 44996
rect 36771 44965 36783 44968
rect 36725 44959 36783 44965
rect 37366 44956 37372 44968
rect 37424 44956 37430 45008
rect 47394 44956 47400 45008
rect 47452 44996 47458 45008
rect 49237 44999 49295 45005
rect 49237 44996 49249 44999
rect 47452 44968 49249 44996
rect 47452 44956 47458 44968
rect 49237 44965 49249 44968
rect 49283 44965 49295 44999
rect 49237 44959 49295 44965
rect 35894 44928 35900 44940
rect 34992 44900 35900 44928
rect 35894 44888 35900 44900
rect 35952 44888 35958 44940
rect 36906 44888 36912 44940
rect 36964 44928 36970 44940
rect 37277 44931 37335 44937
rect 37277 44928 37289 44931
rect 36964 44900 37289 44928
rect 36964 44888 36970 44900
rect 37277 44897 37289 44900
rect 37323 44897 37335 44931
rect 37277 44891 37335 44897
rect 37734 44888 37740 44940
rect 37792 44928 37798 44940
rect 38013 44931 38071 44937
rect 38013 44928 38025 44931
rect 37792 44900 38025 44928
rect 37792 44888 37798 44900
rect 38013 44897 38025 44900
rect 38059 44897 38071 44931
rect 38013 44891 38071 44897
rect 38197 44931 38255 44937
rect 38197 44897 38209 44931
rect 38243 44928 38255 44931
rect 38654 44928 38660 44940
rect 38243 44900 38660 44928
rect 38243 44897 38255 44900
rect 38197 44891 38255 44897
rect 38654 44888 38660 44900
rect 38712 44888 38718 44940
rect 38933 44931 38991 44937
rect 38933 44928 38945 44931
rect 38764 44900 38945 44928
rect 31389 44863 31447 44869
rect 28966 44832 30236 44860
rect 28813 44823 28871 44829
rect 24762 44792 24768 44804
rect 21876 44764 22094 44792
rect 24596 44764 24768 44792
rect 21876 44752 21882 44764
rect 18601 44727 18659 44733
rect 18601 44693 18613 44727
rect 18647 44724 18659 44727
rect 19058 44724 19064 44736
rect 18647 44696 19064 44724
rect 18647 44693 18659 44696
rect 18601 44687 18659 44693
rect 19058 44684 19064 44696
rect 19116 44684 19122 44736
rect 19886 44684 19892 44736
rect 19944 44684 19950 44736
rect 21637 44727 21695 44733
rect 21637 44693 21649 44727
rect 21683 44724 21695 44727
rect 21726 44724 21732 44736
rect 21683 44696 21732 44724
rect 21683 44693 21695 44696
rect 21637 44687 21695 44693
rect 21726 44684 21732 44696
rect 21784 44684 21790 44736
rect 22066 44724 22094 44764
rect 24762 44752 24768 44764
rect 24820 44752 24826 44804
rect 24857 44795 24915 44801
rect 24857 44761 24869 44795
rect 24903 44792 24915 44795
rect 24903 44764 25268 44792
rect 24903 44761 24915 44764
rect 24857 44755 24915 44761
rect 23293 44727 23351 44733
rect 23293 44724 23305 44727
rect 22066 44696 23305 44724
rect 23293 44693 23305 44696
rect 23339 44693 23351 44727
rect 23293 44687 23351 44693
rect 23658 44684 23664 44736
rect 23716 44684 23722 44736
rect 24394 44684 24400 44736
rect 24452 44724 24458 44736
rect 25038 44724 25044 44736
rect 24452 44696 25044 44724
rect 24452 44684 24458 44696
rect 25038 44684 25044 44696
rect 25096 44684 25102 44736
rect 25240 44724 25268 44764
rect 25590 44752 25596 44804
rect 25648 44752 25654 44804
rect 29086 44752 29092 44804
rect 29144 44792 29150 44804
rect 30101 44795 30159 44801
rect 30101 44792 30113 44795
rect 29144 44764 30113 44792
rect 29144 44752 29150 44764
rect 30101 44761 30113 44764
rect 30147 44761 30159 44795
rect 30208 44792 30236 44832
rect 31389 44829 31401 44863
rect 31435 44860 31447 44863
rect 33152 44860 33180 44888
rect 31435 44832 33180 44860
rect 33229 44863 33287 44869
rect 31435 44829 31447 44832
rect 31389 44823 31447 44829
rect 33229 44829 33241 44863
rect 33275 44860 33287 44863
rect 33962 44860 33968 44872
rect 33275 44832 33968 44860
rect 33275 44829 33287 44832
rect 33229 44823 33287 44829
rect 33962 44820 33968 44832
rect 34020 44820 34026 44872
rect 37090 44820 37096 44872
rect 37148 44820 37154 44872
rect 38764 44860 38792 44900
rect 38933 44897 38945 44900
rect 38979 44897 38991 44931
rect 38933 44891 38991 44897
rect 37292 44832 38792 44860
rect 38841 44863 38899 44869
rect 31481 44795 31539 44801
rect 31481 44792 31493 44795
rect 30208 44764 31493 44792
rect 30101 44755 30159 44761
rect 31481 44761 31493 44764
rect 31527 44761 31539 44795
rect 31481 44755 31539 44761
rect 33137 44795 33195 44801
rect 33137 44761 33149 44795
rect 33183 44792 33195 44795
rect 33318 44792 33324 44804
rect 33183 44764 33324 44792
rect 33183 44761 33195 44764
rect 33137 44755 33195 44761
rect 33318 44752 33324 44764
rect 33376 44752 33382 44804
rect 35158 44752 35164 44804
rect 35216 44752 35222 44804
rect 36538 44792 36544 44804
rect 36386 44764 36544 44792
rect 36538 44752 36544 44764
rect 36596 44752 36602 44804
rect 36998 44752 37004 44804
rect 37056 44792 37062 44804
rect 37185 44795 37243 44801
rect 37185 44792 37197 44795
rect 37056 44764 37197 44792
rect 37056 44752 37062 44764
rect 37185 44761 37197 44764
rect 37231 44761 37243 44795
rect 37185 44755 37243 44761
rect 26602 44724 26608 44736
rect 25240 44696 26608 44724
rect 26602 44684 26608 44696
rect 26660 44684 26666 44736
rect 30193 44727 30251 44733
rect 30193 44693 30205 44727
rect 30239 44724 30251 44727
rect 30834 44724 30840 44736
rect 30239 44696 30840 44724
rect 30239 44693 30251 44696
rect 30193 44687 30251 44693
rect 30834 44684 30840 44696
rect 30892 44684 30898 44736
rect 31021 44727 31079 44733
rect 31021 44693 31033 44727
rect 31067 44724 31079 44727
rect 31202 44724 31208 44736
rect 31067 44696 31208 44724
rect 31067 44693 31079 44696
rect 31021 44687 31079 44693
rect 31202 44684 31208 44696
rect 31260 44684 31266 44736
rect 32490 44684 32496 44736
rect 32548 44724 32554 44736
rect 32769 44727 32827 44733
rect 32769 44724 32781 44727
rect 32548 44696 32781 44724
rect 32548 44684 32554 44696
rect 32769 44693 32781 44696
rect 32815 44693 32827 44727
rect 32769 44687 32827 44693
rect 35802 44684 35808 44736
rect 35860 44724 35866 44736
rect 37292 44724 37320 44832
rect 38841 44829 38853 44863
rect 38887 44860 38899 44863
rect 43346 44860 43352 44872
rect 38887 44832 43352 44860
rect 38887 44829 38899 44832
rect 38841 44823 38899 44829
rect 43346 44820 43352 44832
rect 43404 44820 43410 44872
rect 49050 44820 49056 44872
rect 49108 44820 49114 44872
rect 37921 44795 37979 44801
rect 37921 44761 37933 44795
rect 37967 44792 37979 44795
rect 39666 44792 39672 44804
rect 37967 44764 39672 44792
rect 37967 44761 37979 44764
rect 37921 44755 37979 44761
rect 39666 44752 39672 44764
rect 39724 44752 39730 44804
rect 35860 44696 37320 44724
rect 35860 44684 35866 44696
rect 37550 44684 37556 44736
rect 37608 44684 37614 44736
rect 38378 44684 38384 44736
rect 38436 44684 38442 44736
rect 38746 44684 38752 44736
rect 38804 44724 38810 44736
rect 48590 44724 48596 44736
rect 38804 44696 48596 44724
rect 38804 44684 38810 44696
rect 48590 44684 48596 44696
rect 48648 44684 48654 44736
rect 1104 44634 49864 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 27950 44634
rect 28002 44582 28014 44634
rect 28066 44582 28078 44634
rect 28130 44582 28142 44634
rect 28194 44582 28206 44634
rect 28258 44582 37950 44634
rect 38002 44582 38014 44634
rect 38066 44582 38078 44634
rect 38130 44582 38142 44634
rect 38194 44582 38206 44634
rect 38258 44582 47950 44634
rect 48002 44582 48014 44634
rect 48066 44582 48078 44634
rect 48130 44582 48142 44634
rect 48194 44582 48206 44634
rect 48258 44582 49864 44634
rect 1104 44560 49864 44582
rect 2038 44480 2044 44532
rect 2096 44520 2102 44532
rect 3881 44523 3939 44529
rect 3881 44520 3893 44523
rect 2096 44492 3893 44520
rect 2096 44480 2102 44492
rect 3881 44489 3893 44492
rect 3927 44489 3939 44523
rect 3881 44483 3939 44489
rect 9582 44480 9588 44532
rect 9640 44520 9646 44532
rect 10229 44523 10287 44529
rect 10229 44520 10241 44523
rect 9640 44492 10241 44520
rect 9640 44480 9646 44492
rect 10229 44489 10241 44492
rect 10275 44489 10287 44523
rect 10229 44483 10287 44489
rect 14918 44480 14924 44532
rect 14976 44520 14982 44532
rect 15473 44523 15531 44529
rect 15473 44520 15485 44523
rect 14976 44492 15485 44520
rect 14976 44480 14982 44492
rect 15473 44489 15485 44492
rect 15519 44489 15531 44523
rect 15473 44483 15531 44489
rect 17494 44480 17500 44532
rect 17552 44520 17558 44532
rect 17773 44523 17831 44529
rect 17773 44520 17785 44523
rect 17552 44492 17785 44520
rect 17552 44480 17558 44492
rect 17773 44489 17785 44492
rect 17819 44489 17831 44523
rect 20070 44520 20076 44532
rect 17773 44483 17831 44489
rect 18340 44492 20076 44520
rect 5534 44412 5540 44464
rect 5592 44412 5598 44464
rect 6822 44412 6828 44464
rect 6880 44412 6886 44464
rect 1765 44387 1823 44393
rect 1765 44353 1777 44387
rect 1811 44353 1823 44387
rect 1765 44347 1823 44353
rect 1780 44248 1808 44347
rect 3418 44344 3424 44396
rect 3476 44384 3482 44396
rect 3789 44387 3847 44393
rect 3789 44384 3801 44387
rect 3476 44356 3801 44384
rect 3476 44344 3482 44356
rect 3789 44353 3801 44356
rect 3835 44353 3847 44387
rect 3789 44347 3847 44353
rect 5350 44344 5356 44396
rect 5408 44344 5414 44396
rect 10413 44387 10471 44393
rect 10413 44353 10425 44387
rect 10459 44384 10471 44387
rect 12434 44384 12440 44396
rect 10459 44356 12440 44384
rect 10459 44353 10471 44356
rect 10413 44347 10471 44353
rect 12434 44344 12440 44356
rect 12492 44344 12498 44396
rect 15657 44387 15715 44393
rect 15657 44353 15669 44387
rect 15703 44353 15715 44387
rect 15657 44347 15715 44353
rect 2038 44276 2044 44328
rect 2096 44276 2102 44328
rect 15672 44316 15700 44347
rect 16298 44344 16304 44396
rect 16356 44344 16362 44396
rect 17957 44387 18015 44393
rect 17957 44353 17969 44387
rect 18003 44384 18015 44387
rect 18340 44384 18368 44492
rect 20070 44480 20076 44492
rect 20128 44480 20134 44532
rect 21085 44523 21143 44529
rect 21085 44489 21097 44523
rect 21131 44520 21143 44523
rect 21450 44520 21456 44532
rect 21131 44492 21456 44520
rect 21131 44489 21143 44492
rect 21085 44483 21143 44489
rect 21450 44480 21456 44492
rect 21508 44480 21514 44532
rect 22002 44480 22008 44532
rect 22060 44480 22066 44532
rect 24486 44480 24492 44532
rect 24544 44520 24550 44532
rect 25593 44523 25651 44529
rect 25593 44520 25605 44523
rect 24544 44492 25605 44520
rect 24544 44480 24550 44492
rect 25593 44489 25605 44492
rect 25639 44489 25651 44523
rect 25593 44483 25651 44489
rect 27614 44480 27620 44532
rect 27672 44520 27678 44532
rect 28353 44523 28411 44529
rect 28353 44520 28365 44523
rect 27672 44492 28365 44520
rect 27672 44480 27678 44492
rect 28353 44489 28365 44492
rect 28399 44489 28411 44523
rect 28353 44483 28411 44489
rect 28718 44480 28724 44532
rect 28776 44480 28782 44532
rect 29733 44523 29791 44529
rect 29733 44489 29745 44523
rect 29779 44520 29791 44523
rect 30374 44520 30380 44532
rect 29779 44492 30380 44520
rect 29779 44489 29791 44492
rect 29733 44483 29791 44489
rect 30374 44480 30380 44492
rect 30432 44480 30438 44532
rect 30742 44480 30748 44532
rect 30800 44520 30806 44532
rect 31389 44523 31447 44529
rect 31389 44520 31401 44523
rect 30800 44492 31401 44520
rect 30800 44480 30806 44492
rect 31389 44489 31401 44492
rect 31435 44489 31447 44523
rect 31389 44483 31447 44489
rect 32585 44523 32643 44529
rect 32585 44489 32597 44523
rect 32631 44520 32643 44523
rect 34241 44523 34299 44529
rect 34241 44520 34253 44523
rect 32631 44492 34253 44520
rect 32631 44489 32643 44492
rect 32585 44483 32643 44489
rect 34241 44489 34253 44492
rect 34287 44489 34299 44523
rect 34241 44483 34299 44489
rect 34977 44523 35035 44529
rect 34977 44489 34989 44523
rect 35023 44520 35035 44523
rect 36173 44523 36231 44529
rect 36173 44520 36185 44523
rect 35023 44492 36185 44520
rect 35023 44489 35035 44492
rect 34977 44483 35035 44489
rect 36173 44489 36185 44492
rect 36219 44489 36231 44523
rect 36173 44483 36231 44489
rect 36265 44523 36323 44529
rect 36265 44489 36277 44523
rect 36311 44520 36323 44523
rect 37550 44520 37556 44532
rect 36311 44492 37556 44520
rect 36311 44489 36323 44492
rect 36265 44483 36323 44489
rect 37550 44480 37556 44492
rect 37608 44480 37614 44532
rect 37642 44480 37648 44532
rect 37700 44520 37706 44532
rect 37921 44523 37979 44529
rect 37921 44520 37933 44523
rect 37700 44492 37933 44520
rect 37700 44480 37706 44492
rect 37921 44489 37933 44492
rect 37967 44520 37979 44523
rect 38286 44520 38292 44532
rect 37967 44492 38292 44520
rect 37967 44489 37979 44492
rect 37921 44483 37979 44489
rect 38286 44480 38292 44492
rect 38344 44480 38350 44532
rect 39666 44480 39672 44532
rect 39724 44480 39730 44532
rect 49145 44523 49203 44529
rect 49145 44520 49157 44523
rect 45526 44492 49157 44520
rect 20438 44412 20444 44464
rect 20496 44452 20502 44464
rect 22373 44455 22431 44461
rect 22373 44452 22385 44455
rect 20496 44424 22385 44452
rect 20496 44412 20502 44424
rect 22373 44421 22385 44424
rect 22419 44421 22431 44455
rect 23566 44452 23572 44464
rect 22373 44415 22431 44421
rect 22664 44424 23572 44452
rect 21082 44384 21088 44396
rect 18003 44356 18368 44384
rect 19826 44356 21088 44384
rect 18003 44353 18015 44356
rect 17957 44347 18015 44353
rect 21082 44344 21088 44356
rect 21140 44344 21146 44396
rect 21177 44387 21235 44393
rect 21177 44353 21189 44387
rect 21223 44384 21235 44387
rect 22278 44384 22284 44396
rect 21223 44356 22284 44384
rect 21223 44353 21235 44356
rect 21177 44347 21235 44353
rect 22278 44344 22284 44356
rect 22336 44344 22342 44396
rect 18417 44319 18475 44325
rect 18417 44316 18429 44319
rect 15672 44288 17908 44316
rect 11882 44248 11888 44260
rect 1780 44220 11888 44248
rect 11882 44208 11888 44220
rect 11940 44208 11946 44260
rect 14826 44208 14832 44260
rect 14884 44248 14890 44260
rect 16117 44251 16175 44257
rect 16117 44248 16129 44251
rect 14884 44220 16129 44248
rect 14884 44208 14890 44220
rect 16117 44217 16129 44220
rect 16163 44217 16175 44251
rect 16117 44211 16175 44217
rect 6914 44140 6920 44192
rect 6972 44140 6978 44192
rect 17880 44180 17908 44288
rect 17972 44288 18429 44316
rect 17972 44260 18000 44288
rect 18417 44285 18429 44288
rect 18463 44285 18475 44319
rect 18417 44279 18475 44285
rect 18693 44319 18751 44325
rect 18693 44285 18705 44319
rect 18739 44316 18751 44319
rect 19334 44316 19340 44328
rect 18739 44288 19340 44316
rect 18739 44285 18751 44288
rect 18693 44279 18751 44285
rect 17954 44208 17960 44260
rect 18012 44208 18018 44260
rect 18322 44180 18328 44192
rect 17880 44152 18328 44180
rect 18322 44140 18328 44152
rect 18380 44140 18386 44192
rect 18432 44180 18460 44279
rect 19334 44276 19340 44288
rect 19392 44276 19398 44328
rect 21266 44276 21272 44328
rect 21324 44276 21330 44328
rect 22370 44276 22376 44328
rect 22428 44316 22434 44328
rect 22664 44325 22692 44424
rect 23566 44412 23572 44424
rect 23624 44412 23630 44464
rect 27430 44412 27436 44464
rect 27488 44452 27494 44464
rect 27525 44455 27583 44461
rect 27525 44452 27537 44455
rect 27488 44424 27537 44452
rect 27488 44412 27494 44424
rect 27525 44421 27537 44424
rect 27571 44452 27583 44455
rect 27798 44452 27804 44464
rect 27571 44424 27804 44452
rect 27571 44421 27583 44424
rect 27525 44415 27583 44421
rect 27798 44412 27804 44424
rect 27856 44412 27862 44464
rect 28534 44412 28540 44464
rect 28592 44452 28598 44464
rect 30466 44452 30472 44464
rect 28592 44424 28948 44452
rect 28592 44412 28598 44424
rect 25590 44384 25596 44396
rect 24702 44356 25596 44384
rect 25590 44344 25596 44356
rect 25648 44344 25654 44396
rect 25777 44387 25835 44393
rect 25777 44353 25789 44387
rect 25823 44384 25835 44387
rect 26326 44384 26332 44396
rect 25823 44356 26332 44384
rect 25823 44353 25835 44356
rect 25777 44347 25835 44353
rect 26326 44344 26332 44356
rect 26384 44344 26390 44396
rect 27617 44387 27675 44393
rect 27617 44353 27629 44387
rect 27663 44384 27675 44387
rect 27663 44356 27844 44384
rect 27663 44353 27675 44356
rect 27617 44347 27675 44353
rect 22465 44319 22523 44325
rect 22465 44316 22477 44319
rect 22428 44288 22477 44316
rect 22428 44276 22434 44288
rect 22465 44285 22477 44288
rect 22511 44285 22523 44319
rect 22465 44279 22523 44285
rect 22649 44319 22707 44325
rect 22649 44285 22661 44319
rect 22695 44285 22707 44319
rect 22649 44279 22707 44285
rect 23290 44276 23296 44328
rect 23348 44276 23354 44328
rect 23569 44319 23627 44325
rect 23569 44316 23581 44319
rect 23400 44288 23581 44316
rect 20070 44208 20076 44260
rect 20128 44248 20134 44260
rect 20128 44220 20852 44248
rect 20128 44208 20134 44220
rect 19702 44180 19708 44192
rect 18432 44152 19708 44180
rect 19702 44140 19708 44152
rect 19760 44140 19766 44192
rect 20162 44140 20168 44192
rect 20220 44140 20226 44192
rect 20254 44140 20260 44192
rect 20312 44180 20318 44192
rect 20717 44183 20775 44189
rect 20717 44180 20729 44183
rect 20312 44152 20729 44180
rect 20312 44140 20318 44152
rect 20717 44149 20729 44152
rect 20763 44149 20775 44183
rect 20824 44180 20852 44220
rect 21542 44208 21548 44260
rect 21600 44248 21606 44260
rect 23400 44248 23428 44288
rect 23569 44285 23581 44288
rect 23615 44285 23627 44319
rect 23569 44279 23627 44285
rect 23934 44276 23940 44328
rect 23992 44316 23998 44328
rect 24946 44316 24952 44328
rect 23992 44288 24952 44316
rect 23992 44276 23998 44288
rect 24946 44276 24952 44288
rect 25004 44276 25010 44328
rect 25041 44319 25099 44325
rect 25041 44285 25053 44319
rect 25087 44316 25099 44319
rect 26142 44316 26148 44328
rect 25087 44288 26148 44316
rect 25087 44285 25099 44288
rect 25041 44279 25099 44285
rect 26142 44276 26148 44288
rect 26200 44316 26206 44328
rect 27522 44316 27528 44328
rect 26200 44288 27528 44316
rect 26200 44276 26206 44288
rect 27522 44276 27528 44288
rect 27580 44276 27586 44328
rect 27709 44319 27767 44325
rect 27709 44285 27721 44319
rect 27755 44285 27767 44319
rect 27709 44279 27767 44285
rect 21600 44220 23428 44248
rect 21600 44208 21606 44220
rect 25866 44208 25872 44260
rect 25924 44248 25930 44260
rect 27724 44248 27752 44279
rect 25924 44220 27752 44248
rect 27816 44248 27844 44356
rect 28534 44276 28540 44328
rect 28592 44316 28598 44328
rect 28920 44325 28948 44424
rect 30208 44424 30472 44452
rect 30098 44344 30104 44396
rect 30156 44344 30162 44396
rect 28813 44319 28871 44325
rect 28813 44316 28825 44319
rect 28592 44288 28825 44316
rect 28592 44276 28598 44288
rect 28813 44285 28825 44288
rect 28859 44285 28871 44319
rect 28813 44279 28871 44285
rect 28905 44319 28963 44325
rect 28905 44285 28917 44319
rect 28951 44285 28963 44319
rect 28905 44279 28963 44285
rect 30006 44276 30012 44328
rect 30064 44316 30070 44328
rect 30208 44325 30236 44424
rect 30466 44412 30472 44424
rect 30524 44412 30530 44464
rect 31297 44455 31355 44461
rect 31297 44421 31309 44455
rect 31343 44452 31355 44455
rect 34149 44455 34207 44461
rect 31343 44424 34008 44452
rect 31343 44421 31355 44424
rect 31297 44415 31355 44421
rect 32122 44384 32128 44396
rect 30300 44356 32128 44384
rect 30300 44325 30328 44356
rect 32122 44344 32128 44356
rect 32180 44344 32186 44396
rect 32214 44344 32220 44396
rect 32272 44384 32278 44396
rect 32674 44384 32680 44396
rect 32272 44356 32680 44384
rect 32272 44344 32278 44356
rect 32674 44344 32680 44356
rect 32732 44384 32738 44396
rect 32953 44387 33011 44393
rect 32953 44384 32965 44387
rect 32732 44356 32965 44384
rect 32732 44344 32738 44356
rect 32953 44353 32965 44356
rect 32999 44353 33011 44387
rect 32953 44347 33011 44353
rect 33244 44356 33916 44384
rect 30193 44319 30251 44325
rect 30193 44316 30205 44319
rect 30064 44288 30205 44316
rect 30064 44276 30070 44288
rect 30193 44285 30205 44288
rect 30239 44285 30251 44319
rect 30193 44279 30251 44285
rect 30285 44319 30343 44325
rect 30285 44285 30297 44319
rect 30331 44285 30343 44319
rect 31481 44319 31539 44325
rect 31481 44316 31493 44319
rect 30285 44279 30343 44285
rect 30392 44288 31493 44316
rect 28994 44248 29000 44260
rect 27816 44220 29000 44248
rect 25924 44208 25930 44220
rect 28994 44208 29000 44220
rect 29052 44208 29058 44260
rect 29178 44208 29184 44260
rect 29236 44248 29242 44260
rect 30392 44248 30420 44288
rect 31481 44285 31493 44288
rect 31527 44285 31539 44319
rect 31481 44279 31539 44285
rect 32398 44276 32404 44328
rect 32456 44316 32462 44328
rect 32582 44316 32588 44328
rect 32456 44288 32588 44316
rect 32456 44276 32462 44288
rect 32582 44276 32588 44288
rect 32640 44316 32646 44328
rect 33244 44325 33272 44356
rect 33045 44319 33103 44325
rect 33045 44316 33057 44319
rect 32640 44288 33057 44316
rect 32640 44276 32646 44288
rect 33045 44285 33057 44288
rect 33091 44285 33103 44319
rect 33045 44279 33103 44285
rect 33229 44319 33287 44325
rect 33229 44285 33241 44319
rect 33275 44285 33287 44319
rect 33229 44279 33287 44285
rect 33318 44276 33324 44328
rect 33376 44316 33382 44328
rect 33502 44316 33508 44328
rect 33376 44288 33508 44316
rect 33376 44276 33382 44288
rect 33502 44276 33508 44288
rect 33560 44276 33566 44328
rect 29236 44220 30420 44248
rect 29236 44208 29242 44220
rect 30834 44208 30840 44260
rect 30892 44248 30898 44260
rect 33781 44251 33839 44257
rect 33781 44248 33793 44251
rect 30892 44220 33793 44248
rect 30892 44208 30898 44220
rect 33781 44217 33793 44220
rect 33827 44217 33839 44251
rect 33781 44211 33839 44217
rect 23382 44180 23388 44192
rect 20824 44152 23388 44180
rect 20717 44143 20775 44149
rect 23382 44140 23388 44152
rect 23440 44140 23446 44192
rect 26510 44140 26516 44192
rect 26568 44180 26574 44192
rect 27157 44183 27215 44189
rect 27157 44180 27169 44183
rect 26568 44152 27169 44180
rect 26568 44140 26574 44152
rect 27157 44149 27169 44152
rect 27203 44149 27215 44183
rect 27157 44143 27215 44149
rect 28718 44140 28724 44192
rect 28776 44180 28782 44192
rect 30282 44180 30288 44192
rect 28776 44152 30288 44180
rect 28776 44140 28782 44152
rect 30282 44140 30288 44152
rect 30340 44140 30346 44192
rect 30929 44183 30987 44189
rect 30929 44149 30941 44183
rect 30975 44180 30987 44183
rect 33594 44180 33600 44192
rect 30975 44152 33600 44180
rect 30975 44149 30987 44152
rect 30929 44143 30987 44149
rect 33594 44140 33600 44152
rect 33652 44140 33658 44192
rect 33686 44140 33692 44192
rect 33744 44180 33750 44192
rect 33888 44180 33916 44356
rect 33980 44248 34008 44424
rect 34149 44421 34161 44455
rect 34195 44452 34207 44455
rect 38378 44452 38384 44464
rect 34195 44424 35664 44452
rect 34195 44421 34207 44424
rect 34149 44415 34207 44421
rect 35342 44344 35348 44396
rect 35400 44344 35406 44396
rect 35636 44384 35664 44424
rect 36280 44424 38384 44452
rect 36280 44384 36308 44424
rect 38378 44412 38384 44424
rect 38436 44412 38442 44464
rect 35636 44356 36308 44384
rect 37734 44344 37740 44396
rect 37792 44384 37798 44396
rect 37829 44387 37887 44393
rect 37829 44384 37841 44387
rect 37792 44356 37841 44384
rect 37792 44344 37798 44356
rect 37829 44353 37841 44356
rect 37875 44353 37887 44387
rect 37829 44347 37887 44353
rect 40037 44387 40095 44393
rect 40037 44353 40049 44387
rect 40083 44384 40095 44387
rect 45526 44384 45554 44492
rect 49145 44489 49157 44492
rect 49191 44489 49203 44523
rect 49145 44483 49203 44489
rect 40083 44356 45554 44384
rect 40083 44353 40095 44356
rect 40037 44347 40095 44353
rect 49326 44344 49332 44396
rect 49384 44344 49390 44396
rect 34330 44276 34336 44328
rect 34388 44276 34394 44328
rect 34422 44276 34428 44328
rect 34480 44316 34486 44328
rect 35437 44319 35495 44325
rect 35437 44316 35449 44319
rect 34480 44288 35449 44316
rect 34480 44276 34486 44288
rect 35437 44285 35449 44288
rect 35483 44285 35495 44319
rect 35437 44279 35495 44285
rect 35621 44319 35679 44325
rect 35621 44285 35633 44319
rect 35667 44316 35679 44319
rect 35710 44316 35716 44328
rect 35667 44288 35716 44316
rect 35667 44285 35679 44288
rect 35621 44279 35679 44285
rect 35710 44276 35716 44288
rect 35768 44316 35774 44328
rect 36449 44319 36507 44325
rect 35768 44288 36400 44316
rect 35768 44276 35774 44288
rect 36170 44248 36176 44260
rect 33980 44220 36176 44248
rect 36170 44208 36176 44220
rect 36228 44208 36234 44260
rect 34606 44180 34612 44192
rect 33744 44152 34612 44180
rect 33744 44140 33750 44152
rect 34606 44140 34612 44152
rect 34664 44180 34670 44192
rect 35618 44180 35624 44192
rect 34664 44152 35624 44180
rect 34664 44140 34670 44152
rect 35618 44140 35624 44152
rect 35676 44140 35682 44192
rect 35802 44140 35808 44192
rect 35860 44140 35866 44192
rect 36372 44180 36400 44288
rect 36449 44285 36461 44319
rect 36495 44316 36507 44319
rect 36814 44316 36820 44328
rect 36495 44288 36820 44316
rect 36495 44285 36507 44288
rect 36449 44279 36507 44285
rect 36814 44276 36820 44288
rect 36872 44276 36878 44328
rect 37182 44276 37188 44328
rect 37240 44316 37246 44328
rect 37240 44288 37596 44316
rect 37240 44276 37246 44288
rect 37568 44260 37596 44288
rect 38010 44276 38016 44328
rect 38068 44316 38074 44328
rect 39482 44316 39488 44328
rect 38068 44288 39488 44316
rect 38068 44276 38074 44288
rect 39482 44276 39488 44288
rect 39540 44276 39546 44328
rect 40126 44276 40132 44328
rect 40184 44276 40190 44328
rect 40221 44319 40279 44325
rect 40221 44285 40233 44319
rect 40267 44285 40279 44319
rect 40221 44279 40279 44285
rect 37458 44208 37464 44260
rect 37516 44208 37522 44260
rect 37550 44208 37556 44260
rect 37608 44248 37614 44260
rect 40236 44248 40264 44279
rect 37608 44220 40264 44248
rect 37608 44208 37614 44220
rect 38654 44180 38660 44192
rect 36372 44152 38660 44180
rect 38654 44140 38660 44152
rect 38712 44140 38718 44192
rect 1104 44090 49864 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 32950 44090
rect 33002 44038 33014 44090
rect 33066 44038 33078 44090
rect 33130 44038 33142 44090
rect 33194 44038 33206 44090
rect 33258 44038 42950 44090
rect 43002 44038 43014 44090
rect 43066 44038 43078 44090
rect 43130 44038 43142 44090
rect 43194 44038 43206 44090
rect 43258 44038 49864 44090
rect 1104 44016 49864 44038
rect 5810 43936 5816 43988
rect 5868 43976 5874 43988
rect 7837 43979 7895 43985
rect 7837 43976 7849 43979
rect 5868 43948 7849 43976
rect 5868 43936 5874 43948
rect 7837 43945 7849 43948
rect 7883 43945 7895 43979
rect 7837 43939 7895 43945
rect 11054 43936 11060 43988
rect 11112 43976 11118 43988
rect 12897 43979 12955 43985
rect 12897 43976 12909 43979
rect 11112 43948 12909 43976
rect 11112 43936 11118 43948
rect 12897 43945 12909 43948
rect 12943 43945 12955 43979
rect 12897 43939 12955 43945
rect 16114 43936 16120 43988
rect 16172 43936 16178 43988
rect 18877 43979 18935 43985
rect 17236 43948 18828 43976
rect 4706 43868 4712 43920
rect 4764 43868 4770 43920
rect 5718 43868 5724 43920
rect 5776 43868 5782 43920
rect 12250 43868 12256 43920
rect 12308 43868 12314 43920
rect 17236 43908 17264 43948
rect 12406 43880 17264 43908
rect 18800 43908 18828 43948
rect 18877 43945 18889 43979
rect 18923 43976 18935 43979
rect 19978 43976 19984 43988
rect 18923 43948 19984 43976
rect 18923 43945 18935 43948
rect 18877 43939 18935 43945
rect 19978 43936 19984 43948
rect 20036 43936 20042 43988
rect 20070 43936 20076 43988
rect 20128 43976 20134 43988
rect 24118 43976 24124 43988
rect 20128 43948 24124 43976
rect 20128 43936 20134 43948
rect 24118 43936 24124 43948
rect 24176 43936 24182 43988
rect 26602 43936 26608 43988
rect 26660 43936 26666 43988
rect 27985 43979 28043 43985
rect 27985 43945 27997 43979
rect 28031 43976 28043 43979
rect 29546 43976 29552 43988
rect 28031 43948 29552 43976
rect 28031 43945 28043 43948
rect 27985 43939 28043 43945
rect 29546 43936 29552 43948
rect 29604 43936 29610 43988
rect 31294 43936 31300 43988
rect 31352 43976 31358 43988
rect 49234 43976 49240 43988
rect 31352 43948 49240 43976
rect 31352 43936 31358 43948
rect 49234 43936 49240 43948
rect 49292 43936 49298 43988
rect 19242 43908 19248 43920
rect 18800 43880 19248 43908
rect 5537 43775 5595 43781
rect 5537 43741 5549 43775
rect 5583 43772 5595 43775
rect 9582 43772 9588 43784
rect 5583 43744 9588 43772
rect 5583 43741 5595 43744
rect 5537 43735 5595 43741
rect 9582 43732 9588 43744
rect 9640 43732 9646 43784
rect 12069 43775 12127 43781
rect 12069 43741 12081 43775
rect 12115 43772 12127 43775
rect 12406 43772 12434 43880
rect 19242 43868 19248 43880
rect 19300 43868 19306 43920
rect 32674 43868 32680 43920
rect 32732 43908 32738 43920
rect 33962 43908 33968 43920
rect 32732 43880 33968 43908
rect 32732 43868 32738 43880
rect 33962 43868 33968 43880
rect 34020 43868 34026 43920
rect 38654 43868 38660 43920
rect 38712 43908 38718 43920
rect 39025 43911 39083 43917
rect 39025 43908 39037 43911
rect 38712 43880 39037 43908
rect 38712 43868 38718 43880
rect 39025 43877 39037 43880
rect 39071 43877 39083 43911
rect 39025 43871 39083 43877
rect 16850 43800 16856 43852
rect 16908 43840 16914 43852
rect 17129 43843 17187 43849
rect 17129 43840 17141 43843
rect 16908 43812 17141 43840
rect 16908 43800 16914 43812
rect 17129 43809 17141 43812
rect 17175 43840 17187 43843
rect 17862 43840 17868 43852
rect 17175 43812 17868 43840
rect 17175 43809 17187 43812
rect 17129 43803 17187 43809
rect 17862 43800 17868 43812
rect 17920 43800 17926 43852
rect 18414 43800 18420 43852
rect 18472 43840 18478 43852
rect 18690 43840 18696 43852
rect 18472 43812 18696 43840
rect 18472 43800 18478 43812
rect 18690 43800 18696 43812
rect 18748 43800 18754 43852
rect 19334 43800 19340 43852
rect 19392 43840 19398 43852
rect 20165 43843 20223 43849
rect 20165 43840 20177 43843
rect 19392 43812 20177 43840
rect 19392 43800 19398 43812
rect 20165 43809 20177 43812
rect 20211 43840 20223 43843
rect 21358 43840 21364 43852
rect 20211 43812 21364 43840
rect 20211 43809 20223 43812
rect 20165 43803 20223 43809
rect 21358 43800 21364 43812
rect 21416 43800 21422 43852
rect 22281 43843 22339 43849
rect 22281 43809 22293 43843
rect 22327 43840 22339 43843
rect 22462 43840 22468 43852
rect 22327 43812 22468 43840
rect 22327 43809 22339 43812
rect 22281 43803 22339 43809
rect 22462 43800 22468 43812
rect 22520 43800 22526 43852
rect 23382 43800 23388 43852
rect 23440 43800 23446 43852
rect 24857 43843 24915 43849
rect 24857 43809 24869 43843
rect 24903 43840 24915 43843
rect 27430 43840 27436 43852
rect 24903 43812 27436 43840
rect 24903 43809 24915 43812
rect 24857 43803 24915 43809
rect 27430 43800 27436 43812
rect 27488 43800 27494 43852
rect 28629 43843 28687 43849
rect 28629 43809 28641 43843
rect 28675 43840 28687 43843
rect 29362 43840 29368 43852
rect 28675 43812 29368 43840
rect 28675 43809 28687 43812
rect 28629 43803 28687 43809
rect 29362 43800 29368 43812
rect 29420 43800 29426 43852
rect 30006 43800 30012 43852
rect 30064 43840 30070 43852
rect 30285 43843 30343 43849
rect 30285 43840 30297 43843
rect 30064 43812 30297 43840
rect 30064 43800 30070 43812
rect 30285 43809 30297 43812
rect 30331 43809 30343 43843
rect 30285 43803 30343 43809
rect 31297 43843 31355 43849
rect 31297 43809 31309 43843
rect 31343 43840 31355 43843
rect 31938 43840 31944 43852
rect 31343 43812 31944 43840
rect 31343 43809 31355 43812
rect 31297 43803 31355 43809
rect 31938 43800 31944 43812
rect 31996 43800 32002 43852
rect 32214 43800 32220 43852
rect 32272 43840 32278 43852
rect 32582 43840 32588 43852
rect 32272 43812 32588 43840
rect 32272 43800 32278 43812
rect 32582 43800 32588 43812
rect 32640 43840 32646 43852
rect 32640 43812 32996 43840
rect 32640 43800 32646 43812
rect 12115 43744 12434 43772
rect 15657 43775 15715 43781
rect 12115 43741 12127 43744
rect 12069 43735 12127 43741
rect 15657 43741 15669 43775
rect 15703 43772 15715 43775
rect 15930 43772 15936 43784
rect 15703 43744 15936 43772
rect 15703 43741 15715 43744
rect 15657 43735 15715 43741
rect 15930 43732 15936 43744
rect 15988 43732 15994 43784
rect 16301 43775 16359 43781
rect 16301 43741 16313 43775
rect 16347 43772 16359 43775
rect 16482 43772 16488 43784
rect 16347 43744 16488 43772
rect 16347 43741 16359 43744
rect 16301 43735 16359 43741
rect 16482 43732 16488 43744
rect 16540 43732 16546 43784
rect 22097 43775 22155 43781
rect 22097 43741 22109 43775
rect 22143 43772 22155 43775
rect 22646 43772 22652 43784
rect 22143 43744 22652 43772
rect 22143 43741 22155 43744
rect 22097 43735 22155 43741
rect 22646 43732 22652 43744
rect 22704 43732 22710 43784
rect 23293 43775 23351 43781
rect 23293 43741 23305 43775
rect 23339 43772 23351 43775
rect 24578 43772 24584 43784
rect 23339 43744 24584 43772
rect 23339 43741 23351 43744
rect 23293 43735 23351 43741
rect 24578 43732 24584 43744
rect 24636 43732 24642 43784
rect 30193 43775 30251 43781
rect 30193 43741 30205 43775
rect 30239 43772 30251 43775
rect 30926 43772 30932 43784
rect 30239 43744 30932 43772
rect 30239 43741 30251 43744
rect 30193 43735 30251 43741
rect 30926 43732 30932 43744
rect 30984 43732 30990 43784
rect 32968 43772 32996 43812
rect 33042 43800 33048 43852
rect 33100 43840 33106 43852
rect 33686 43840 33692 43852
rect 33100 43812 33692 43840
rect 33100 43800 33106 43812
rect 33686 43800 33692 43812
rect 33744 43800 33750 43852
rect 33778 43800 33784 43852
rect 33836 43840 33842 43852
rect 34149 43843 34207 43849
rect 34149 43840 34161 43843
rect 33836 43812 34161 43840
rect 33836 43800 33842 43812
rect 34149 43809 34161 43812
rect 34195 43809 34207 43843
rect 34149 43803 34207 43809
rect 34882 43800 34888 43852
rect 34940 43840 34946 43852
rect 35069 43843 35127 43849
rect 35069 43840 35081 43843
rect 34940 43812 35081 43840
rect 34940 43800 34946 43812
rect 35069 43809 35081 43812
rect 35115 43809 35127 43843
rect 35069 43803 35127 43809
rect 35345 43843 35403 43849
rect 35345 43809 35357 43843
rect 35391 43840 35403 43843
rect 35710 43840 35716 43852
rect 35391 43812 35716 43840
rect 35391 43809 35403 43812
rect 35345 43803 35403 43809
rect 35710 43800 35716 43812
rect 35768 43800 35774 43852
rect 36538 43840 36544 43852
rect 36464 43812 36544 43840
rect 34057 43775 34115 43781
rect 34057 43772 34069 43775
rect 32968 43744 34069 43772
rect 34057 43741 34069 43744
rect 34103 43741 34115 43775
rect 36464 43758 36492 43812
rect 36538 43800 36544 43812
rect 36596 43840 36602 43852
rect 36596 43812 36676 43840
rect 36596 43800 36602 43812
rect 34057 43735 34115 43741
rect 4525 43707 4583 43713
rect 4525 43673 4537 43707
rect 4571 43704 4583 43707
rect 4798 43704 4804 43716
rect 4571 43676 4804 43704
rect 4571 43673 4583 43676
rect 4525 43667 4583 43673
rect 4798 43664 4804 43676
rect 4856 43664 4862 43716
rect 7745 43707 7803 43713
rect 7745 43673 7757 43707
rect 7791 43704 7803 43707
rect 12805 43707 12863 43713
rect 7791 43676 12434 43704
rect 7791 43673 7803 43676
rect 7745 43667 7803 43673
rect 12406 43636 12434 43676
rect 12805 43673 12817 43707
rect 12851 43704 12863 43707
rect 13630 43704 13636 43716
rect 12851 43676 13636 43704
rect 12851 43673 12863 43676
rect 12805 43667 12863 43673
rect 13630 43664 13636 43676
rect 13688 43664 13694 43716
rect 17405 43707 17463 43713
rect 17405 43673 17417 43707
rect 17451 43673 17463 43707
rect 17405 43667 17463 43673
rect 14550 43636 14556 43648
rect 12406 43608 14556 43636
rect 14550 43596 14556 43608
rect 14608 43596 14614 43648
rect 17420 43636 17448 43667
rect 18414 43664 18420 43716
rect 18472 43664 18478 43716
rect 19334 43664 19340 43716
rect 19392 43704 19398 43716
rect 22005 43707 22063 43713
rect 19392 43676 21772 43704
rect 19392 43664 19398 43676
rect 18322 43636 18328 43648
rect 17420 43608 18328 43636
rect 18322 43596 18328 43608
rect 18380 43596 18386 43648
rect 19518 43596 19524 43648
rect 19576 43596 19582 43648
rect 19886 43596 19892 43648
rect 19944 43596 19950 43648
rect 19981 43639 20039 43645
rect 19981 43605 19993 43639
rect 20027 43636 20039 43639
rect 20714 43636 20720 43648
rect 20027 43608 20720 43636
rect 20027 43605 20039 43608
rect 19981 43599 20039 43605
rect 20714 43596 20720 43608
rect 20772 43596 20778 43648
rect 21266 43596 21272 43648
rect 21324 43636 21330 43648
rect 21637 43639 21695 43645
rect 21637 43636 21649 43639
rect 21324 43608 21649 43636
rect 21324 43596 21330 43608
rect 21637 43605 21649 43608
rect 21683 43605 21695 43639
rect 21744 43636 21772 43676
rect 22005 43673 22017 43707
rect 22051 43704 22063 43707
rect 24486 43704 24492 43716
rect 22051 43676 24492 43704
rect 22051 43673 22063 43676
rect 22005 43667 22063 43673
rect 24486 43664 24492 43676
rect 24544 43664 24550 43716
rect 24670 43664 24676 43716
rect 24728 43704 24734 43716
rect 24728 43676 24992 43704
rect 24728 43664 24734 43676
rect 22833 43639 22891 43645
rect 22833 43636 22845 43639
rect 21744 43608 22845 43636
rect 21637 43599 21695 43605
rect 22833 43605 22845 43608
rect 22879 43605 22891 43639
rect 22833 43599 22891 43605
rect 23201 43639 23259 43645
rect 23201 43605 23213 43639
rect 23247 43636 23259 43639
rect 24854 43636 24860 43648
rect 23247 43608 24860 43636
rect 23247 43605 23259 43608
rect 23201 43599 23259 43605
rect 24854 43596 24860 43608
rect 24912 43596 24918 43648
rect 24964 43636 24992 43676
rect 25038 43664 25044 43716
rect 25096 43704 25102 43716
rect 25133 43707 25191 43713
rect 25133 43704 25145 43707
rect 25096 43676 25145 43704
rect 25096 43664 25102 43676
rect 25133 43673 25145 43676
rect 25179 43704 25191 43707
rect 25222 43704 25228 43716
rect 25179 43676 25228 43704
rect 25179 43673 25191 43676
rect 25133 43667 25191 43673
rect 25222 43664 25228 43676
rect 25280 43664 25286 43716
rect 25590 43664 25596 43716
rect 25648 43664 25654 43716
rect 27706 43664 27712 43716
rect 27764 43704 27770 43716
rect 28353 43707 28411 43713
rect 28353 43704 28365 43707
rect 27764 43676 28365 43704
rect 27764 43664 27770 43676
rect 28353 43673 28365 43676
rect 28399 43673 28411 43707
rect 28353 43667 28411 43673
rect 30101 43707 30159 43713
rect 30101 43673 30113 43707
rect 30147 43704 30159 43707
rect 31018 43704 31024 43716
rect 30147 43676 31024 43704
rect 30147 43673 30159 43676
rect 30101 43667 30159 43673
rect 31018 43664 31024 43676
rect 31076 43664 31082 43716
rect 31570 43664 31576 43716
rect 31628 43664 31634 43716
rect 32858 43704 32864 43716
rect 32798 43676 32864 43704
rect 32858 43664 32864 43676
rect 32916 43704 32922 43716
rect 33226 43704 33232 43716
rect 32916 43676 33232 43704
rect 32916 43664 32922 43676
rect 33226 43664 33232 43676
rect 33284 43664 33290 43716
rect 36648 43704 36676 43812
rect 37274 43800 37280 43852
rect 37332 43800 37338 43852
rect 33612 43676 35756 43704
rect 36648 43676 37504 43704
rect 28445 43639 28503 43645
rect 28445 43636 28457 43639
rect 24964 43608 28457 43636
rect 28445 43605 28457 43608
rect 28491 43605 28503 43639
rect 28445 43599 28503 43605
rect 29733 43639 29791 43645
rect 29733 43605 29745 43639
rect 29779 43636 29791 43639
rect 30742 43636 30748 43648
rect 29779 43608 30748 43636
rect 29779 43605 29791 43608
rect 29733 43599 29791 43605
rect 30742 43596 30748 43608
rect 30800 43596 30806 43648
rect 32582 43596 32588 43648
rect 32640 43636 32646 43648
rect 33045 43639 33103 43645
rect 33045 43636 33057 43639
rect 32640 43608 33057 43636
rect 32640 43596 32646 43608
rect 33045 43605 33057 43608
rect 33091 43636 33103 43639
rect 33502 43636 33508 43648
rect 33091 43608 33508 43636
rect 33091 43605 33103 43608
rect 33045 43599 33103 43605
rect 33502 43596 33508 43608
rect 33560 43596 33566 43648
rect 33612 43645 33640 43676
rect 33597 43639 33655 43645
rect 33597 43605 33609 43639
rect 33643 43605 33655 43639
rect 33597 43599 33655 43605
rect 33962 43596 33968 43648
rect 34020 43596 34026 43648
rect 35728 43636 35756 43676
rect 36354 43636 36360 43648
rect 35728 43608 36360 43636
rect 36354 43596 36360 43608
rect 36412 43596 36418 43648
rect 36814 43596 36820 43648
rect 36872 43596 36878 43648
rect 37476 43636 37504 43676
rect 37550 43664 37556 43716
rect 37608 43664 37614 43716
rect 37660 43676 38042 43704
rect 37660 43636 37688 43676
rect 37476 43608 37688 43636
rect 37936 43636 37964 43676
rect 38838 43636 38844 43648
rect 37936 43608 38844 43636
rect 38838 43596 38844 43608
rect 38896 43596 38902 43648
rect 1104 43546 49864 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 27950 43546
rect 28002 43494 28014 43546
rect 28066 43494 28078 43546
rect 28130 43494 28142 43546
rect 28194 43494 28206 43546
rect 28258 43494 37950 43546
rect 38002 43494 38014 43546
rect 38066 43494 38078 43546
rect 38130 43494 38142 43546
rect 38194 43494 38206 43546
rect 38258 43494 47950 43546
rect 48002 43494 48014 43546
rect 48066 43494 48078 43546
rect 48130 43494 48142 43546
rect 48194 43494 48206 43546
rect 48258 43494 49864 43546
rect 1104 43472 49864 43494
rect 4062 43392 4068 43444
rect 4120 43432 4126 43444
rect 5629 43435 5687 43441
rect 5629 43432 5641 43435
rect 4120 43404 5641 43432
rect 4120 43392 4126 43404
rect 5629 43401 5641 43404
rect 5675 43401 5687 43435
rect 5629 43395 5687 43401
rect 8662 43392 8668 43444
rect 8720 43392 8726 43444
rect 15102 43392 15108 43444
rect 15160 43432 15166 43444
rect 15565 43435 15623 43441
rect 15565 43432 15577 43435
rect 15160 43404 15577 43432
rect 15160 43392 15166 43404
rect 15565 43401 15577 43404
rect 15611 43401 15623 43435
rect 15565 43395 15623 43401
rect 15930 43392 15936 43444
rect 15988 43392 15994 43444
rect 18877 43435 18935 43441
rect 18877 43401 18889 43435
rect 18923 43432 18935 43435
rect 20254 43432 20260 43444
rect 18923 43404 20260 43432
rect 18923 43401 18935 43404
rect 18877 43395 18935 43401
rect 20254 43392 20260 43404
rect 20312 43392 20318 43444
rect 21358 43392 21364 43444
rect 21416 43432 21422 43444
rect 21453 43435 21511 43441
rect 21453 43432 21465 43435
rect 21416 43404 21465 43432
rect 21416 43392 21422 43404
rect 21453 43401 21465 43404
rect 21499 43401 21511 43435
rect 26418 43432 26424 43444
rect 21453 43395 21511 43401
rect 22756 43404 26424 43432
rect 6914 43364 6920 43376
rect 1780 43336 6920 43364
rect 1780 43305 1808 43336
rect 6914 43324 6920 43336
rect 6972 43324 6978 43376
rect 19981 43367 20039 43373
rect 19981 43333 19993 43367
rect 20027 43364 20039 43367
rect 20070 43364 20076 43376
rect 20027 43336 20076 43364
rect 20027 43333 20039 43336
rect 19981 43327 20039 43333
rect 20070 43324 20076 43336
rect 20128 43324 20134 43376
rect 22462 43364 22468 43376
rect 22388 43336 22468 43364
rect 1765 43299 1823 43305
rect 1765 43265 1777 43299
rect 1811 43265 1823 43299
rect 1765 43259 1823 43265
rect 5537 43299 5595 43305
rect 5537 43265 5549 43299
rect 5583 43265 5595 43299
rect 5537 43259 5595 43265
rect 8573 43299 8631 43305
rect 8573 43265 8585 43299
rect 8619 43296 8631 43299
rect 16025 43299 16083 43305
rect 8619 43268 12434 43296
rect 8619 43265 8631 43268
rect 8573 43259 8631 43265
rect 1302 43188 1308 43240
rect 1360 43228 1366 43240
rect 2041 43231 2099 43237
rect 2041 43228 2053 43231
rect 1360 43200 2053 43228
rect 1360 43188 1366 43200
rect 2041 43197 2053 43200
rect 2087 43197 2099 43231
rect 5552 43228 5580 43259
rect 9490 43228 9496 43240
rect 5552 43200 9496 43228
rect 2041 43191 2099 43197
rect 9490 43188 9496 43200
rect 9548 43188 9554 43240
rect 12406 43160 12434 43268
rect 16025 43265 16037 43299
rect 16071 43296 16083 43299
rect 17770 43296 17776 43308
rect 16071 43268 17776 43296
rect 16071 43265 16083 43268
rect 16025 43259 16083 43265
rect 17770 43256 17776 43268
rect 17828 43256 17834 43308
rect 18874 43256 18880 43308
rect 18932 43296 18938 43308
rect 18969 43299 19027 43305
rect 18969 43296 18981 43299
rect 18932 43268 18981 43296
rect 18932 43256 18938 43268
rect 18969 43265 18981 43268
rect 19015 43265 19027 43299
rect 18969 43259 19027 43265
rect 19702 43256 19708 43308
rect 19760 43256 19766 43308
rect 21082 43256 21088 43308
rect 21140 43256 21146 43308
rect 16209 43231 16267 43237
rect 16209 43197 16221 43231
rect 16255 43228 16267 43231
rect 18322 43228 18328 43240
rect 16255 43200 18328 43228
rect 16255 43197 16267 43200
rect 16209 43191 16267 43197
rect 18322 43188 18328 43200
rect 18380 43188 18386 43240
rect 19153 43231 19211 43237
rect 19153 43197 19165 43231
rect 19199 43197 19211 43231
rect 19153 43191 19211 43197
rect 17034 43160 17040 43172
rect 12406 43132 17040 43160
rect 17034 43120 17040 43132
rect 17092 43120 17098 43172
rect 18506 43052 18512 43104
rect 18564 43052 18570 43104
rect 19168 43092 19196 43191
rect 20622 43188 20628 43240
rect 20680 43228 20686 43240
rect 22388 43228 22416 43336
rect 22462 43324 22468 43336
rect 22520 43324 22526 43376
rect 22756 43373 22784 43404
rect 26418 43392 26424 43404
rect 26476 43392 26482 43444
rect 26694 43392 26700 43444
rect 26752 43432 26758 43444
rect 27157 43435 27215 43441
rect 27157 43432 27169 43435
rect 26752 43404 27169 43432
rect 26752 43392 26758 43404
rect 27157 43401 27169 43404
rect 27203 43401 27215 43435
rect 27157 43395 27215 43401
rect 27522 43392 27528 43444
rect 27580 43432 27586 43444
rect 28258 43432 28264 43444
rect 27580 43404 28264 43432
rect 27580 43392 27586 43404
rect 28258 43392 28264 43404
rect 28316 43392 28322 43444
rect 31205 43435 31263 43441
rect 31205 43401 31217 43435
rect 31251 43432 31263 43435
rect 31570 43432 31576 43444
rect 31251 43404 31576 43432
rect 31251 43401 31263 43404
rect 31205 43395 31263 43401
rect 31570 43392 31576 43404
rect 31628 43392 31634 43444
rect 33226 43392 33232 43444
rect 33284 43432 33290 43444
rect 33284 43404 33916 43432
rect 33284 43392 33290 43404
rect 22741 43367 22799 43373
rect 22741 43333 22753 43367
rect 22787 43333 22799 43367
rect 22741 43327 22799 43333
rect 22830 43324 22836 43376
rect 22888 43364 22894 43376
rect 22888 43336 23230 43364
rect 22888 43324 22894 43336
rect 24946 43324 24952 43376
rect 25004 43324 25010 43376
rect 25590 43324 25596 43376
rect 25648 43324 25654 43376
rect 32858 43364 32864 43376
rect 30958 43336 32864 43364
rect 32858 43324 32864 43336
rect 32916 43324 32922 43376
rect 33888 43364 33916 43404
rect 35526 43392 35532 43444
rect 35584 43432 35590 43444
rect 35897 43435 35955 43441
rect 35897 43432 35909 43435
rect 35584 43404 35909 43432
rect 35584 43392 35590 43404
rect 35897 43401 35909 43404
rect 35943 43401 35955 43435
rect 35897 43395 35955 43401
rect 35989 43435 36047 43441
rect 35989 43401 36001 43435
rect 36035 43432 36047 43435
rect 36262 43432 36268 43444
rect 36035 43404 36268 43432
rect 36035 43401 36047 43404
rect 35989 43395 36047 43401
rect 36262 43392 36268 43404
rect 36320 43392 36326 43444
rect 49234 43392 49240 43444
rect 49292 43392 49298 43444
rect 35158 43364 35164 43376
rect 33810 43336 35164 43364
rect 35158 43324 35164 43336
rect 35216 43324 35222 43376
rect 27246 43256 27252 43308
rect 27304 43296 27310 43308
rect 27341 43299 27399 43305
rect 27341 43296 27353 43299
rect 27304 43268 27353 43296
rect 27304 43256 27310 43268
rect 27341 43265 27353 43268
rect 27387 43265 27399 43299
rect 27341 43259 27399 43265
rect 29454 43256 29460 43308
rect 29512 43256 29518 43308
rect 31938 43256 31944 43308
rect 31996 43296 32002 43308
rect 32309 43299 32367 43305
rect 32309 43296 32321 43299
rect 31996 43268 32321 43296
rect 31996 43256 32002 43268
rect 32309 43265 32321 43268
rect 32355 43265 32367 43299
rect 32309 43259 32367 43265
rect 35069 43299 35127 43305
rect 35069 43265 35081 43299
rect 35115 43296 35127 43299
rect 35342 43296 35348 43308
rect 35115 43268 35348 43296
rect 35115 43265 35127 43268
rect 35069 43259 35127 43265
rect 35342 43256 35348 43268
rect 35400 43256 35406 43308
rect 49142 43256 49148 43308
rect 49200 43256 49206 43308
rect 20680 43200 22416 43228
rect 20680 43188 20686 43200
rect 21634 43092 21640 43104
rect 19168 43064 21640 43092
rect 21634 43052 21640 43064
rect 21692 43052 21698 43104
rect 22066 43092 22094 43200
rect 22462 43188 22468 43240
rect 22520 43228 22526 43240
rect 23290 43228 23296 43240
rect 22520 43200 23296 43228
rect 22520 43188 22526 43200
rect 23290 43188 23296 43200
rect 23348 43228 23354 43240
rect 24673 43231 24731 43237
rect 24673 43228 24685 43231
rect 23348 43200 24685 43228
rect 23348 43188 23354 43200
rect 24673 43197 24685 43200
rect 24719 43197 24731 43231
rect 24673 43191 24731 43197
rect 29362 43188 29368 43240
rect 29420 43228 29426 43240
rect 29733 43231 29791 43237
rect 29733 43228 29745 43231
rect 29420 43200 29745 43228
rect 29420 43188 29426 43200
rect 29733 43197 29745 43200
rect 29779 43228 29791 43231
rect 32585 43231 32643 43237
rect 29779 43200 31754 43228
rect 29779 43197 29791 43200
rect 29733 43191 29791 43197
rect 24213 43095 24271 43101
rect 24213 43092 24225 43095
rect 22066 43064 24225 43092
rect 24213 43061 24225 43064
rect 24259 43061 24271 43095
rect 24213 43055 24271 43061
rect 24394 43052 24400 43104
rect 24452 43092 24458 43104
rect 31110 43092 31116 43104
rect 24452 43064 31116 43092
rect 24452 43052 24458 43064
rect 31110 43052 31116 43064
rect 31168 43092 31174 43104
rect 31294 43092 31300 43104
rect 31168 43064 31300 43092
rect 31168 43052 31174 43064
rect 31294 43052 31300 43064
rect 31352 43052 31358 43104
rect 31726 43092 31754 43200
rect 32585 43197 32597 43231
rect 32631 43228 32643 43231
rect 33042 43228 33048 43240
rect 32631 43200 33048 43228
rect 32631 43197 32643 43200
rect 32585 43191 32643 43197
rect 33042 43188 33048 43200
rect 33100 43188 33106 43240
rect 36170 43188 36176 43240
rect 36228 43188 36234 43240
rect 34057 43095 34115 43101
rect 34057 43092 34069 43095
rect 31726 43064 34069 43092
rect 34057 43061 34069 43064
rect 34103 43092 34115 43095
rect 34330 43092 34336 43104
rect 34103 43064 34336 43092
rect 34103 43061 34115 43064
rect 34057 43055 34115 43061
rect 34330 43052 34336 43064
rect 34388 43052 34394 43104
rect 35529 43095 35587 43101
rect 35529 43061 35541 43095
rect 35575 43092 35587 43095
rect 36998 43092 37004 43104
rect 35575 43064 37004 43092
rect 35575 43061 35587 43064
rect 35529 43055 35587 43061
rect 36998 43052 37004 43064
rect 37056 43052 37062 43104
rect 1104 43002 49864 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 32950 43002
rect 33002 42950 33014 43002
rect 33066 42950 33078 43002
rect 33130 42950 33142 43002
rect 33194 42950 33206 43002
rect 33258 42950 42950 43002
rect 43002 42950 43014 43002
rect 43066 42950 43078 43002
rect 43130 42950 43142 43002
rect 43194 42950 43206 43002
rect 43258 42950 49864 43002
rect 1104 42928 49864 42950
rect 21634 42848 21640 42900
rect 21692 42888 21698 42900
rect 21692 42860 23520 42888
rect 21692 42848 21698 42860
rect 13354 42780 13360 42832
rect 13412 42820 13418 42832
rect 18141 42823 18199 42829
rect 18141 42820 18153 42823
rect 13412 42792 18153 42820
rect 13412 42780 13418 42792
rect 18141 42789 18153 42792
rect 18187 42789 18199 42823
rect 20162 42820 20168 42832
rect 18141 42783 18199 42789
rect 18800 42792 20168 42820
rect 1302 42712 1308 42764
rect 1360 42752 1366 42764
rect 2041 42755 2099 42761
rect 2041 42752 2053 42755
rect 1360 42724 2053 42752
rect 1360 42712 1366 42724
rect 2041 42721 2053 42724
rect 2087 42721 2099 42755
rect 2041 42715 2099 42721
rect 17052 42724 18460 42752
rect 17052 42693 17080 42724
rect 1765 42687 1823 42693
rect 1765 42653 1777 42687
rect 1811 42684 1823 42687
rect 15289 42687 15347 42693
rect 15289 42684 15301 42687
rect 1811 42656 15301 42684
rect 1811 42653 1823 42656
rect 1765 42647 1823 42653
rect 15289 42653 15301 42656
rect 15335 42653 15347 42687
rect 15289 42647 15347 42653
rect 17037 42687 17095 42693
rect 17037 42653 17049 42687
rect 17083 42653 17095 42687
rect 17037 42647 17095 42653
rect 17494 42644 17500 42696
rect 17552 42684 17558 42696
rect 17681 42687 17739 42693
rect 17681 42684 17693 42687
rect 17552 42656 17693 42684
rect 17552 42644 17558 42656
rect 17681 42653 17693 42656
rect 17727 42653 17739 42687
rect 17681 42647 17739 42653
rect 15102 42576 15108 42628
rect 15160 42576 15166 42628
rect 16666 42576 16672 42628
rect 16724 42616 16730 42628
rect 18432 42616 18460 42724
rect 18598 42712 18604 42764
rect 18656 42712 18662 42764
rect 18800 42761 18828 42792
rect 20162 42780 20168 42792
rect 20220 42780 20226 42832
rect 23492 42820 23520 42860
rect 25038 42848 25044 42900
rect 25096 42888 25102 42900
rect 25961 42891 26019 42897
rect 25961 42888 25973 42891
rect 25096 42860 25973 42888
rect 25096 42848 25102 42860
rect 25961 42857 25973 42860
rect 26007 42857 26019 42891
rect 25961 42851 26019 42857
rect 26694 42848 26700 42900
rect 26752 42848 26758 42900
rect 27522 42848 27528 42900
rect 27580 42888 27586 42900
rect 27696 42891 27754 42897
rect 27696 42888 27708 42891
rect 27580 42860 27708 42888
rect 27580 42848 27586 42860
rect 27696 42857 27708 42860
rect 27742 42888 27754 42891
rect 29270 42888 29276 42900
rect 27742 42860 29276 42888
rect 27742 42857 27754 42860
rect 27696 42851 27754 42857
rect 29270 42848 29276 42860
rect 29328 42848 29334 42900
rect 30558 42848 30564 42900
rect 30616 42888 30622 42900
rect 30834 42888 30840 42900
rect 30616 42860 30840 42888
rect 30616 42848 30622 42860
rect 30834 42848 30840 42860
rect 30892 42848 30898 42900
rect 31478 42848 31484 42900
rect 31536 42888 31542 42900
rect 35424 42891 35482 42897
rect 31536 42860 33916 42888
rect 31536 42848 31542 42860
rect 25130 42820 25136 42832
rect 23492 42792 25136 42820
rect 25130 42780 25136 42792
rect 25188 42780 25194 42832
rect 26602 42820 26608 42832
rect 25240 42792 26608 42820
rect 18785 42755 18843 42761
rect 18785 42721 18797 42755
rect 18831 42721 18843 42755
rect 18785 42715 18843 42721
rect 19426 42712 19432 42764
rect 19484 42752 19490 42764
rect 19702 42752 19708 42764
rect 19484 42724 19708 42752
rect 19484 42712 19490 42724
rect 19702 42712 19708 42724
rect 19760 42752 19766 42764
rect 20257 42755 20315 42761
rect 20257 42752 20269 42755
rect 19760 42724 20269 42752
rect 19760 42712 19766 42724
rect 20257 42721 20269 42724
rect 20303 42752 20315 42755
rect 20530 42752 20536 42764
rect 20303 42724 20536 42752
rect 20303 42721 20315 42724
rect 20257 42715 20315 42721
rect 20530 42712 20536 42724
rect 20588 42712 20594 42764
rect 22554 42712 22560 42764
rect 22612 42752 22618 42764
rect 22830 42752 22836 42764
rect 22612 42724 22836 42752
rect 22612 42712 22618 42724
rect 22830 42712 22836 42724
rect 22888 42712 22894 42764
rect 23290 42712 23296 42764
rect 23348 42712 23354 42764
rect 25240 42761 25268 42792
rect 26602 42780 26608 42792
rect 26660 42780 26666 42832
rect 25225 42755 25283 42761
rect 25225 42721 25237 42755
rect 25271 42721 25283 42755
rect 25225 42715 25283 42721
rect 25590 42712 25596 42764
rect 25648 42752 25654 42764
rect 25648 42724 27016 42752
rect 25648 42712 25654 42724
rect 18509 42687 18567 42693
rect 18509 42653 18521 42687
rect 18555 42684 18567 42687
rect 19518 42684 19524 42696
rect 18555 42656 19524 42684
rect 18555 42653 18567 42656
rect 18509 42647 18567 42653
rect 19518 42644 19524 42656
rect 19576 42644 19582 42696
rect 19613 42687 19671 42693
rect 19613 42653 19625 42687
rect 19659 42684 19671 42687
rect 19978 42684 19984 42696
rect 19659 42656 19984 42684
rect 19659 42653 19671 42656
rect 19613 42647 19671 42653
rect 19978 42644 19984 42656
rect 20036 42644 20042 42696
rect 21818 42644 21824 42696
rect 21876 42684 21882 42696
rect 22848 42684 22876 42712
rect 23566 42684 23572 42696
rect 21876 42656 22508 42684
rect 22848 42656 23572 42684
rect 21876 42644 21882 42656
rect 20533 42619 20591 42625
rect 16724 42588 17540 42616
rect 18432 42588 20484 42616
rect 16724 42576 16730 42588
rect 16390 42508 16396 42560
rect 16448 42548 16454 42560
rect 17512 42557 17540 42588
rect 16853 42551 16911 42557
rect 16853 42548 16865 42551
rect 16448 42520 16865 42548
rect 16448 42508 16454 42520
rect 16853 42517 16865 42520
rect 16899 42517 16911 42551
rect 16853 42511 16911 42517
rect 17497 42551 17555 42557
rect 17497 42517 17509 42551
rect 17543 42517 17555 42551
rect 17497 42511 17555 42517
rect 18966 42508 18972 42560
rect 19024 42548 19030 42560
rect 19429 42551 19487 42557
rect 19429 42548 19441 42551
rect 19024 42520 19441 42548
rect 19024 42508 19030 42520
rect 19429 42517 19441 42520
rect 19475 42517 19487 42551
rect 20456 42548 20484 42588
rect 20533 42585 20545 42619
rect 20579 42616 20591 42619
rect 20622 42616 20628 42628
rect 20579 42588 20628 42616
rect 20579 42585 20591 42588
rect 20533 42579 20591 42585
rect 20622 42576 20628 42588
rect 20680 42576 20686 42628
rect 21082 42576 21088 42628
rect 21140 42576 21146 42628
rect 22480 42625 22508 42656
rect 23566 42644 23572 42656
rect 23624 42644 23630 42696
rect 24949 42687 25007 42693
rect 24949 42653 24961 42687
rect 24995 42684 25007 42687
rect 25038 42684 25044 42696
rect 24995 42656 25044 42684
rect 24995 42653 25007 42656
rect 24949 42647 25007 42653
rect 25038 42644 25044 42656
rect 25096 42644 25102 42696
rect 26878 42644 26884 42696
rect 26936 42644 26942 42696
rect 26988 42684 27016 42724
rect 27430 42712 27436 42764
rect 27488 42752 27494 42764
rect 29454 42752 29460 42764
rect 27488 42724 29460 42752
rect 27488 42712 27494 42724
rect 29454 42712 29460 42724
rect 29512 42752 29518 42764
rect 30469 42755 30527 42761
rect 30469 42752 30481 42755
rect 29512 42724 30481 42752
rect 29512 42712 29518 42724
rect 30469 42721 30481 42724
rect 30515 42721 30527 42755
rect 30469 42715 30527 42721
rect 31113 42755 31171 42761
rect 31113 42721 31125 42755
rect 31159 42752 31171 42755
rect 31938 42752 31944 42764
rect 31159 42724 31944 42752
rect 31159 42721 31171 42724
rect 31113 42715 31171 42721
rect 31938 42712 31944 42724
rect 31996 42712 32002 42764
rect 32766 42712 32772 42764
rect 32824 42752 32830 42764
rect 32861 42755 32919 42761
rect 32861 42752 32873 42755
rect 32824 42724 32873 42752
rect 32824 42712 32830 42724
rect 32861 42721 32873 42724
rect 32907 42721 32919 42755
rect 32861 42715 32919 42721
rect 33594 42712 33600 42764
rect 33652 42752 33658 42764
rect 33888 42761 33916 42860
rect 35424 42857 35436 42891
rect 35470 42888 35482 42891
rect 36814 42888 36820 42900
rect 35470 42860 36820 42888
rect 35470 42857 35482 42860
rect 35424 42851 35482 42857
rect 36814 42848 36820 42860
rect 36872 42848 36878 42900
rect 33781 42755 33839 42761
rect 33781 42752 33793 42755
rect 33652 42724 33793 42752
rect 33652 42712 33658 42724
rect 33781 42721 33793 42724
rect 33827 42721 33839 42755
rect 33781 42715 33839 42721
rect 33873 42755 33931 42761
rect 33873 42721 33885 42755
rect 33919 42721 33931 42755
rect 33873 42715 33931 42721
rect 34882 42712 34888 42764
rect 34940 42752 34946 42764
rect 35161 42755 35219 42761
rect 35161 42752 35173 42755
rect 34940 42724 35173 42752
rect 34940 42712 34946 42724
rect 35161 42721 35173 42724
rect 35207 42721 35219 42755
rect 35161 42715 35219 42721
rect 26988 42656 27292 42684
rect 22465 42619 22523 42625
rect 22465 42585 22477 42619
rect 22511 42616 22523 42619
rect 27264 42616 27292 42656
rect 36538 42644 36544 42696
rect 36596 42644 36602 42696
rect 49050 42644 49056 42696
rect 49108 42644 49114 42696
rect 29733 42619 29791 42625
rect 29733 42616 29745 42619
rect 22511 42588 27200 42616
rect 27264 42588 28198 42616
rect 29012 42588 29745 42616
rect 22511 42585 22523 42588
rect 22465 42579 22523 42585
rect 27172 42560 27200 42588
rect 21542 42548 21548 42560
rect 20456 42520 21548 42548
rect 19429 42511 19487 42517
rect 21542 42508 21548 42520
rect 21600 42508 21606 42560
rect 21910 42508 21916 42560
rect 21968 42548 21974 42560
rect 22005 42551 22063 42557
rect 22005 42548 22017 42551
rect 21968 42520 22017 42548
rect 21968 42508 21974 42520
rect 22005 42517 22017 42520
rect 22051 42517 22063 42551
rect 22005 42511 22063 42517
rect 23750 42508 23756 42560
rect 23808 42548 23814 42560
rect 24581 42551 24639 42557
rect 24581 42548 24593 42551
rect 23808 42520 24593 42548
rect 23808 42508 23814 42520
rect 24581 42517 24593 42520
rect 24627 42517 24639 42551
rect 24581 42511 24639 42517
rect 25038 42508 25044 42560
rect 25096 42508 25102 42560
rect 27154 42508 27160 42560
rect 27212 42548 27218 42560
rect 27522 42548 27528 42560
rect 27212 42520 27528 42548
rect 27212 42508 27218 42520
rect 27522 42508 27528 42520
rect 27580 42548 27586 42560
rect 29012 42548 29040 42588
rect 29733 42585 29745 42588
rect 29779 42585 29791 42619
rect 29733 42579 29791 42585
rect 31389 42619 31447 42625
rect 31389 42585 31401 42619
rect 31435 42616 31447 42619
rect 31662 42616 31668 42628
rect 31435 42588 31668 42616
rect 31435 42585 31447 42588
rect 31389 42579 31447 42585
rect 27580 42520 29040 42548
rect 27580 42508 27586 42520
rect 29178 42508 29184 42560
rect 29236 42508 29242 42560
rect 29748 42548 29776 42579
rect 31662 42576 31668 42588
rect 31720 42576 31726 42628
rect 32858 42616 32864 42628
rect 32614 42588 32864 42616
rect 32858 42576 32864 42588
rect 32916 42576 32922 42628
rect 32398 42548 32404 42560
rect 29748 42520 32404 42548
rect 32398 42508 32404 42520
rect 32456 42508 32462 42560
rect 33321 42551 33379 42557
rect 33321 42517 33333 42551
rect 33367 42548 33379 42551
rect 33594 42548 33600 42560
rect 33367 42520 33600 42548
rect 33367 42517 33379 42520
rect 33321 42511 33379 42517
rect 33594 42508 33600 42520
rect 33652 42508 33658 42560
rect 33686 42508 33692 42560
rect 33744 42508 33750 42560
rect 33778 42508 33784 42560
rect 33836 42548 33842 42560
rect 36909 42551 36967 42557
rect 36909 42548 36921 42551
rect 33836 42520 36921 42548
rect 33836 42508 33842 42520
rect 36909 42517 36921 42520
rect 36955 42548 36967 42551
rect 37826 42548 37832 42560
rect 36955 42520 37832 42548
rect 36955 42517 36967 42520
rect 36909 42511 36967 42517
rect 37826 42508 37832 42520
rect 37884 42508 37890 42560
rect 47210 42508 47216 42560
rect 47268 42548 47274 42560
rect 49237 42551 49295 42557
rect 49237 42548 49249 42551
rect 47268 42520 49249 42548
rect 47268 42508 47274 42520
rect 49237 42517 49249 42520
rect 49283 42517 49295 42551
rect 49237 42511 49295 42517
rect 1104 42458 49864 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 27950 42458
rect 28002 42406 28014 42458
rect 28066 42406 28078 42458
rect 28130 42406 28142 42458
rect 28194 42406 28206 42458
rect 28258 42406 37950 42458
rect 38002 42406 38014 42458
rect 38066 42406 38078 42458
rect 38130 42406 38142 42458
rect 38194 42406 38206 42458
rect 38258 42406 47950 42458
rect 48002 42406 48014 42458
rect 48066 42406 48078 42458
rect 48130 42406 48142 42458
rect 48194 42406 48206 42458
rect 48258 42406 49864 42458
rect 1104 42384 49864 42406
rect 11882 42304 11888 42356
rect 11940 42304 11946 42356
rect 15102 42304 15108 42356
rect 15160 42344 15166 42356
rect 24394 42344 24400 42356
rect 15160 42316 24400 42344
rect 15160 42304 15166 42316
rect 24394 42304 24400 42316
rect 24452 42304 24458 42356
rect 24946 42304 24952 42356
rect 25004 42344 25010 42356
rect 26145 42347 26203 42353
rect 26145 42344 26157 42347
rect 25004 42316 26157 42344
rect 25004 42304 25010 42316
rect 26145 42313 26157 42316
rect 26191 42313 26203 42347
rect 26145 42307 26203 42313
rect 27798 42304 27804 42356
rect 27856 42344 27862 42356
rect 29089 42347 29147 42353
rect 29089 42344 29101 42347
rect 27856 42316 29101 42344
rect 27856 42304 27862 42316
rect 29089 42313 29101 42316
rect 29135 42313 29147 42347
rect 29089 42307 29147 42313
rect 29181 42347 29239 42353
rect 29181 42313 29193 42347
rect 29227 42344 29239 42347
rect 29638 42344 29644 42356
rect 29227 42316 29644 42344
rect 29227 42313 29239 42316
rect 29181 42307 29239 42313
rect 29638 42304 29644 42316
rect 29696 42304 29702 42356
rect 31478 42344 31484 42356
rect 30208 42316 31484 42344
rect 18414 42276 18420 42288
rect 18354 42262 18420 42276
rect 18340 42248 18420 42262
rect 11793 42211 11851 42217
rect 11793 42177 11805 42211
rect 11839 42208 11851 42211
rect 11839 42180 12434 42208
rect 11839 42177 11851 42180
rect 11793 42171 11851 42177
rect 12406 42072 12434 42180
rect 16298 42168 16304 42220
rect 16356 42168 16362 42220
rect 16850 42168 16856 42220
rect 16908 42168 16914 42220
rect 17126 42100 17132 42152
rect 17184 42100 17190 42152
rect 17678 42100 17684 42152
rect 17736 42140 17742 42152
rect 18340 42140 18368 42248
rect 18414 42236 18420 42248
rect 18472 42236 18478 42288
rect 19797 42279 19855 42285
rect 19797 42245 19809 42279
rect 19843 42276 19855 42279
rect 21818 42276 21824 42288
rect 19843 42248 21824 42276
rect 19843 42245 19855 42248
rect 19797 42239 19855 42245
rect 21818 42236 21824 42248
rect 21876 42236 21882 42288
rect 22554 42236 22560 42288
rect 22612 42276 22618 42288
rect 22612 42248 22770 42276
rect 22612 42236 22618 42248
rect 23566 42236 23572 42288
rect 23624 42276 23630 42288
rect 23624 42248 25162 42276
rect 23624 42236 23630 42248
rect 27154 42236 27160 42288
rect 27212 42236 27218 42288
rect 30208 42285 30236 42316
rect 31478 42304 31484 42316
rect 31536 42304 31542 42356
rect 31662 42304 31668 42356
rect 31720 42304 31726 42356
rect 32858 42344 32864 42356
rect 32692 42316 32864 42344
rect 30193 42279 30251 42285
rect 30193 42245 30205 42279
rect 30239 42245 30251 42279
rect 31846 42276 31852 42288
rect 31418 42248 31852 42276
rect 30193 42239 30251 42245
rect 31846 42236 31852 42248
rect 31904 42276 31910 42288
rect 32692 42276 32720 42316
rect 32858 42304 32864 42316
rect 32916 42304 32922 42356
rect 34238 42304 34244 42356
rect 34296 42344 34302 42356
rect 35069 42347 35127 42353
rect 35069 42344 35081 42347
rect 34296 42316 35081 42344
rect 34296 42304 34302 42316
rect 35069 42313 35081 42316
rect 35115 42344 35127 42347
rect 35115 42316 38056 42344
rect 35115 42313 35127 42316
rect 35069 42307 35127 42313
rect 31904 42248 32720 42276
rect 31904 42236 31910 42248
rect 32766 42236 32772 42288
rect 32824 42276 32830 42288
rect 33597 42279 33655 42285
rect 33597 42276 33609 42279
rect 32824 42248 33609 42276
rect 32824 42236 32830 42248
rect 33597 42245 33609 42248
rect 33643 42245 33655 42279
rect 35158 42276 35164 42288
rect 34822 42248 35164 42276
rect 33597 42239 33655 42245
rect 35158 42236 35164 42248
rect 35216 42236 35222 42288
rect 36262 42236 36268 42288
rect 36320 42276 36326 42288
rect 36449 42279 36507 42285
rect 36449 42276 36461 42279
rect 36320 42248 36461 42276
rect 36320 42236 36326 42248
rect 36449 42245 36461 42248
rect 36495 42245 36507 42279
rect 37921 42279 37979 42285
rect 37921 42276 37933 42279
rect 36449 42239 36507 42245
rect 36556 42248 37933 42276
rect 19242 42168 19248 42220
rect 19300 42208 19306 42220
rect 20346 42208 20352 42220
rect 19300 42180 20352 42208
rect 19300 42168 19306 42180
rect 20346 42168 20352 42180
rect 20404 42168 20410 42220
rect 20530 42168 20536 42220
rect 20588 42208 20594 42220
rect 22005 42211 22063 42217
rect 22005 42208 22017 42211
rect 20588 42180 22017 42208
rect 20588 42168 20594 42180
rect 22005 42177 22017 42180
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 26878 42168 26884 42220
rect 26936 42208 26942 42220
rect 29546 42208 29552 42220
rect 26936 42180 29552 42208
rect 26936 42168 26942 42180
rect 29546 42168 29552 42180
rect 29604 42168 29610 42220
rect 35250 42168 35256 42220
rect 35308 42208 35314 42220
rect 36556 42208 36584 42248
rect 37921 42245 37933 42248
rect 37967 42245 37979 42279
rect 37921 42239 37979 42245
rect 35308 42180 36584 42208
rect 37829 42211 37887 42217
rect 35308 42168 35314 42180
rect 37829 42177 37841 42211
rect 37875 42177 37887 42211
rect 37829 42171 37887 42177
rect 17736 42112 18368 42140
rect 17736 42100 17742 42112
rect 21910 42100 21916 42152
rect 21968 42140 21974 42152
rect 22281 42143 22339 42149
rect 22281 42140 22293 42143
rect 21968 42112 22293 42140
rect 21968 42100 21974 42112
rect 22281 42109 22293 42112
rect 22327 42109 22339 42143
rect 22281 42103 22339 42109
rect 24397 42143 24455 42149
rect 24397 42109 24409 42143
rect 24443 42140 24455 42143
rect 24762 42140 24768 42152
rect 24443 42112 24768 42140
rect 24443 42109 24455 42112
rect 24397 42103 24455 42109
rect 24762 42100 24768 42112
rect 24820 42140 24826 42152
rect 25130 42140 25136 42152
rect 24820 42112 25136 42140
rect 24820 42100 24826 42112
rect 25130 42100 25136 42112
rect 25188 42140 25194 42152
rect 27062 42140 27068 42152
rect 25188 42112 27068 42140
rect 25188 42100 25194 42112
rect 27062 42100 27068 42112
rect 27120 42140 27126 42152
rect 27893 42143 27951 42149
rect 27893 42140 27905 42143
rect 27120 42112 27905 42140
rect 27120 42100 27126 42112
rect 27893 42109 27905 42112
rect 27939 42109 27951 42143
rect 27893 42103 27951 42109
rect 29270 42100 29276 42152
rect 29328 42100 29334 42152
rect 29924 42143 29982 42149
rect 29924 42109 29936 42143
rect 29970 42109 29982 42143
rect 31938 42140 31944 42152
rect 29924 42103 29982 42109
rect 31220 42112 31944 42140
rect 16850 42072 16856 42084
rect 12406 42044 16856 42072
rect 16850 42032 16856 42044
rect 16908 42032 16914 42084
rect 18322 42032 18328 42084
rect 18380 42072 18386 42084
rect 18601 42075 18659 42081
rect 18601 42072 18613 42075
rect 18380 42044 18613 42072
rect 18380 42032 18386 42044
rect 18601 42041 18613 42044
rect 18647 42041 18659 42075
rect 18601 42035 18659 42041
rect 20438 42032 20444 42084
rect 20496 42072 20502 42084
rect 21082 42072 21088 42084
rect 20496 42044 21088 42072
rect 20496 42032 20502 42044
rect 21082 42032 21088 42044
rect 21140 42032 21146 42084
rect 21542 42032 21548 42084
rect 21600 42072 21606 42084
rect 21818 42072 21824 42084
rect 21600 42044 21824 42072
rect 21600 42032 21606 42044
rect 21818 42032 21824 42044
rect 21876 42032 21882 42084
rect 28721 42075 28779 42081
rect 28721 42041 28733 42075
rect 28767 42072 28779 42075
rect 29638 42072 29644 42084
rect 28767 42044 29644 42072
rect 28767 42041 28779 42044
rect 28721 42035 28779 42041
rect 29638 42032 29644 42044
rect 29696 42032 29702 42084
rect 15286 41964 15292 42016
rect 15344 42004 15350 42016
rect 16117 42007 16175 42013
rect 16117 42004 16129 42007
rect 15344 41976 16129 42004
rect 15344 41964 15350 41976
rect 16117 41973 16129 41976
rect 16163 41973 16175 42007
rect 16117 41967 16175 41973
rect 20806 41964 20812 42016
rect 20864 42004 20870 42016
rect 21361 42007 21419 42013
rect 21361 42004 21373 42007
rect 20864 41976 21373 42004
rect 20864 41964 20870 41976
rect 21361 41973 21373 41976
rect 21407 41973 21419 42007
rect 21361 41967 21419 41973
rect 23750 41964 23756 42016
rect 23808 41964 23814 42016
rect 24210 41964 24216 42016
rect 24268 42004 24274 42016
rect 24660 42007 24718 42013
rect 24660 42004 24672 42007
rect 24268 41976 24672 42004
rect 24268 41964 24274 41976
rect 24660 41973 24672 41976
rect 24706 42004 24718 42007
rect 26602 42004 26608 42016
rect 24706 41976 26608 42004
rect 24706 41973 24718 41976
rect 24660 41967 24718 41973
rect 26602 41964 26608 41976
rect 26660 41964 26666 42016
rect 29932 42004 29960 42103
rect 31220 42004 31248 42112
rect 31938 42100 31944 42112
rect 31996 42140 32002 42152
rect 32858 42140 32864 42152
rect 31996 42112 32864 42140
rect 31996 42100 32002 42112
rect 32858 42100 32864 42112
rect 32916 42140 32922 42152
rect 33321 42143 33379 42149
rect 33321 42140 33333 42143
rect 32916 42112 33333 42140
rect 32916 42100 32922 42112
rect 33321 42109 33333 42112
rect 33367 42109 33379 42143
rect 33321 42103 33379 42109
rect 36078 42100 36084 42152
rect 36136 42140 36142 42152
rect 36541 42143 36599 42149
rect 36541 42140 36553 42143
rect 36136 42112 36553 42140
rect 36136 42100 36142 42112
rect 36541 42109 36553 42112
rect 36587 42109 36599 42143
rect 36541 42103 36599 42109
rect 36630 42100 36636 42152
rect 36688 42100 36694 42152
rect 31294 42032 31300 42084
rect 31352 42072 31358 42084
rect 37844 42072 37872 42171
rect 38028 42149 38056 42316
rect 38013 42143 38071 42149
rect 38013 42109 38025 42143
rect 38059 42109 38071 42143
rect 38013 42103 38071 42109
rect 31352 42044 33456 42072
rect 31352 42032 31358 42044
rect 29932 41976 31248 42004
rect 33428 42004 33456 42044
rect 34624 42044 37872 42072
rect 34624 42004 34652 42044
rect 33428 41976 34652 42004
rect 35158 41964 35164 42016
rect 35216 42004 35222 42016
rect 36081 42007 36139 42013
rect 36081 42004 36093 42007
rect 35216 41976 36093 42004
rect 35216 41964 35222 41976
rect 36081 41973 36093 41976
rect 36127 41973 36139 42007
rect 36081 41967 36139 41973
rect 37461 42007 37519 42013
rect 37461 41973 37473 42007
rect 37507 42004 37519 42007
rect 39482 42004 39488 42016
rect 37507 41976 39488 42004
rect 37507 41973 37519 41976
rect 37461 41967 37519 41973
rect 39482 41964 39488 41976
rect 39540 41964 39546 42016
rect 1104 41914 49864 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 32950 41914
rect 33002 41862 33014 41914
rect 33066 41862 33078 41914
rect 33130 41862 33142 41914
rect 33194 41862 33206 41914
rect 33258 41862 42950 41914
rect 43002 41862 43014 41914
rect 43066 41862 43078 41914
rect 43130 41862 43142 41914
rect 43194 41862 43206 41914
rect 43258 41862 49864 41914
rect 1104 41840 49864 41862
rect 11974 41760 11980 41812
rect 12032 41760 12038 41812
rect 13722 41760 13728 41812
rect 13780 41800 13786 41812
rect 15013 41803 15071 41809
rect 15013 41800 15025 41803
rect 13780 41772 15025 41800
rect 13780 41760 13786 41772
rect 15013 41769 15025 41772
rect 15059 41769 15071 41803
rect 15013 41763 15071 41769
rect 16298 41760 16304 41812
rect 16356 41800 16362 41812
rect 21634 41800 21640 41812
rect 16356 41772 21640 41800
rect 16356 41760 16362 41772
rect 21634 41760 21640 41772
rect 21692 41760 21698 41812
rect 21910 41760 21916 41812
rect 21968 41760 21974 41812
rect 22084 41803 22142 41809
rect 22084 41769 22096 41803
rect 22130 41800 22142 41803
rect 22130 41772 23244 41800
rect 22130 41769 22142 41772
rect 22084 41763 22142 41769
rect 9490 41692 9496 41744
rect 9548 41732 9554 41744
rect 13081 41735 13139 41741
rect 13081 41732 13093 41735
rect 9548 41704 13093 41732
rect 9548 41692 9554 41704
rect 13081 41701 13093 41704
rect 13127 41701 13139 41735
rect 20717 41735 20775 41741
rect 20717 41732 20729 41735
rect 13081 41695 13139 41701
rect 19904 41704 20729 41732
rect 1302 41624 1308 41676
rect 1360 41664 1366 41676
rect 2041 41667 2099 41673
rect 2041 41664 2053 41667
rect 1360 41636 2053 41664
rect 1360 41624 1366 41636
rect 2041 41633 2053 41636
rect 2087 41633 2099 41667
rect 14274 41664 14280 41676
rect 2041 41627 2099 41633
rect 12176 41636 14280 41664
rect 1765 41599 1823 41605
rect 1765 41565 1777 41599
rect 1811 41596 1823 41599
rect 11054 41596 11060 41608
rect 1811 41568 11060 41596
rect 1811 41565 1823 41568
rect 1765 41559 1823 41565
rect 11054 41556 11060 41568
rect 11112 41556 11118 41608
rect 12176 41605 12204 41636
rect 14274 41624 14280 41636
rect 14332 41624 14338 41676
rect 15657 41667 15715 41673
rect 15657 41633 15669 41667
rect 15703 41664 15715 41667
rect 16022 41664 16028 41676
rect 15703 41636 16028 41664
rect 15703 41633 15715 41636
rect 15657 41627 15715 41633
rect 16022 41624 16028 41636
rect 16080 41624 16086 41676
rect 19904 41673 19932 41704
rect 20717 41701 20729 41704
rect 20763 41732 20775 41735
rect 21174 41732 21180 41744
rect 20763 41704 21180 41732
rect 20763 41701 20775 41704
rect 20717 41695 20775 41701
rect 21174 41692 21180 41704
rect 21232 41692 21238 41744
rect 21928 41732 21956 41760
rect 21468 41704 21956 41732
rect 23216 41732 23244 41772
rect 24486 41760 24492 41812
rect 24544 41800 24550 41812
rect 27617 41803 27675 41809
rect 27617 41800 27629 41803
rect 24544 41772 27629 41800
rect 24544 41760 24550 41772
rect 27617 41769 27629 41772
rect 27663 41769 27675 41803
rect 30098 41800 30104 41812
rect 27617 41763 27675 41769
rect 28828 41772 30104 41800
rect 23750 41732 23756 41744
rect 23216 41704 23756 41732
rect 19889 41667 19947 41673
rect 19889 41664 19901 41667
rect 16500 41636 19901 41664
rect 12161 41599 12219 41605
rect 12161 41565 12173 41599
rect 12207 41565 12219 41599
rect 12161 41559 12219 41565
rect 13265 41599 13323 41605
rect 13265 41565 13277 41599
rect 13311 41565 13323 41599
rect 13265 41559 13323 41565
rect 15381 41599 15439 41605
rect 15381 41565 15393 41599
rect 15427 41596 15439 41599
rect 16393 41599 16451 41605
rect 16393 41596 16405 41599
rect 15427 41568 16405 41596
rect 15427 41565 15439 41568
rect 15381 41559 15439 41565
rect 16393 41565 16405 41568
rect 16439 41565 16451 41599
rect 16393 41559 16451 41565
rect 13280 41528 13308 41559
rect 13354 41528 13360 41540
rect 13280 41500 13360 41528
rect 13354 41488 13360 41500
rect 13412 41488 13418 41540
rect 15473 41531 15531 41537
rect 15473 41497 15485 41531
rect 15519 41528 15531 41531
rect 16114 41528 16120 41540
rect 15519 41500 16120 41528
rect 15519 41497 15531 41500
rect 15473 41491 15531 41497
rect 16114 41488 16120 41500
rect 16172 41488 16178 41540
rect 3602 41420 3608 41472
rect 3660 41460 3666 41472
rect 16500 41460 16528 41636
rect 19889 41633 19901 41636
rect 19935 41633 19947 41667
rect 19889 41627 19947 41633
rect 20073 41667 20131 41673
rect 20073 41633 20085 41667
rect 20119 41664 20131 41667
rect 20622 41664 20628 41676
rect 20119 41636 20628 41664
rect 20119 41633 20131 41636
rect 20073 41627 20131 41633
rect 20622 41624 20628 41636
rect 20680 41624 20686 41676
rect 21266 41624 21272 41676
rect 21324 41624 21330 41676
rect 21468 41673 21496 41704
rect 23750 41692 23756 41704
rect 23808 41692 23814 41744
rect 26602 41692 26608 41744
rect 26660 41732 26666 41744
rect 27338 41732 27344 41744
rect 26660 41704 27344 41732
rect 26660 41692 26666 41704
rect 27338 41692 27344 41704
rect 27396 41692 27402 41744
rect 21453 41667 21511 41673
rect 21453 41633 21465 41667
rect 21499 41633 21511 41667
rect 21453 41627 21511 41633
rect 21821 41667 21879 41673
rect 21821 41633 21833 41667
rect 21867 41664 21879 41667
rect 22462 41664 22468 41676
rect 21867 41636 22468 41664
rect 21867 41633 21879 41636
rect 21821 41627 21879 41633
rect 22462 41624 22468 41636
rect 22520 41624 22526 41676
rect 23290 41624 23296 41676
rect 23348 41664 23354 41676
rect 23569 41667 23627 41673
rect 23569 41664 23581 41667
rect 23348 41636 23581 41664
rect 23348 41624 23354 41636
rect 23569 41633 23581 41636
rect 23615 41633 23627 41667
rect 23569 41627 23627 41633
rect 24578 41624 24584 41676
rect 24636 41664 24642 41676
rect 24857 41667 24915 41673
rect 24857 41664 24869 41667
rect 24636 41636 24869 41664
rect 24636 41624 24642 41636
rect 24857 41633 24869 41636
rect 24903 41664 24915 41667
rect 25130 41664 25136 41676
rect 24903 41636 25136 41664
rect 24903 41633 24915 41636
rect 24857 41627 24915 41633
rect 25130 41624 25136 41636
rect 25188 41624 25194 41676
rect 26418 41624 26424 41676
rect 26476 41664 26482 41676
rect 28169 41667 28227 41673
rect 28169 41664 28181 41667
rect 26476 41636 28181 41664
rect 26476 41624 26482 41636
rect 28169 41633 28181 41636
rect 28215 41633 28227 41667
rect 28169 41627 28227 41633
rect 17221 41599 17279 41605
rect 17221 41565 17233 41599
rect 17267 41596 17279 41599
rect 18506 41596 18512 41608
rect 17267 41568 18512 41596
rect 17267 41565 17279 41568
rect 17221 41559 17279 41565
rect 18506 41556 18512 41568
rect 18564 41556 18570 41608
rect 18874 41556 18880 41608
rect 18932 41556 18938 41608
rect 19797 41599 19855 41605
rect 19797 41565 19809 41599
rect 19843 41596 19855 41599
rect 21082 41596 21088 41608
rect 19843 41568 21088 41596
rect 19843 41565 19855 41568
rect 19797 41559 19855 41565
rect 21082 41556 21088 41568
rect 21140 41556 21146 41608
rect 24118 41556 24124 41608
rect 24176 41596 24182 41608
rect 24765 41599 24823 41605
rect 24176 41592 24716 41596
rect 24765 41592 24777 41599
rect 24176 41568 24777 41592
rect 24176 41556 24182 41568
rect 24688 41565 24777 41568
rect 24811 41565 24823 41599
rect 26970 41596 26976 41608
rect 24688 41564 24823 41565
rect 24765 41559 24823 41564
rect 26436 41568 26976 41596
rect 21177 41531 21235 41537
rect 21177 41528 21189 41531
rect 19444 41500 21189 41528
rect 3660 41432 16528 41460
rect 3660 41420 3666 41432
rect 17034 41420 17040 41472
rect 17092 41460 17098 41472
rect 17586 41460 17592 41472
rect 17092 41432 17592 41460
rect 17092 41420 17098 41432
rect 17586 41420 17592 41432
rect 17644 41420 17650 41472
rect 19444 41469 19472 41500
rect 21177 41497 21189 41500
rect 21223 41497 21235 41531
rect 21177 41491 21235 41497
rect 22002 41488 22008 41540
rect 22060 41528 22066 41540
rect 22554 41528 22560 41540
rect 22060 41500 22560 41528
rect 22060 41488 22066 41500
rect 22554 41488 22560 41500
rect 22612 41488 22618 41540
rect 23750 41488 23756 41540
rect 23808 41528 23814 41540
rect 25133 41531 25191 41537
rect 23808 41500 24716 41528
rect 23808 41488 23814 41500
rect 19429 41463 19487 41469
rect 19429 41429 19441 41463
rect 19475 41429 19487 41463
rect 19429 41423 19487 41429
rect 20809 41463 20867 41469
rect 20809 41429 20821 41463
rect 20855 41460 20867 41463
rect 20990 41460 20996 41472
rect 20855 41432 20996 41460
rect 20855 41429 20867 41432
rect 20809 41423 20867 41429
rect 20990 41420 20996 41432
rect 21048 41420 21054 41472
rect 22738 41420 22744 41472
rect 22796 41460 22802 41472
rect 24581 41463 24639 41469
rect 24581 41460 24593 41463
rect 22796 41432 24593 41460
rect 22796 41420 22802 41432
rect 24581 41429 24593 41432
rect 24627 41429 24639 41463
rect 24688 41460 24716 41500
rect 25133 41497 25145 41531
rect 25179 41528 25191 41531
rect 25406 41528 25412 41540
rect 25179 41500 25412 41528
rect 25179 41497 25191 41500
rect 25133 41491 25191 41497
rect 25406 41488 25412 41500
rect 25464 41488 25470 41540
rect 25590 41488 25596 41540
rect 25648 41488 25654 41540
rect 26436 41460 26464 41568
rect 26970 41556 26976 41568
rect 27028 41596 27034 41608
rect 27338 41596 27344 41608
rect 27028 41568 27344 41596
rect 27028 41556 27034 41568
rect 27338 41556 27344 41568
rect 27396 41556 27402 41608
rect 28077 41599 28135 41605
rect 28077 41596 28089 41599
rect 27724 41568 28089 41596
rect 24688 41432 26464 41460
rect 24581 41423 24639 41429
rect 26602 41420 26608 41472
rect 26660 41460 26666 41472
rect 27065 41463 27123 41469
rect 27065 41460 27077 41463
rect 26660 41432 27077 41460
rect 26660 41420 26666 41432
rect 27065 41429 27077 41432
rect 27111 41460 27123 41463
rect 27724 41460 27752 41568
rect 28077 41565 28089 41568
rect 28123 41596 28135 41599
rect 28828 41596 28856 41772
rect 30098 41760 30104 41772
rect 30156 41760 30162 41812
rect 31478 41760 31484 41812
rect 31536 41760 31542 41812
rect 32582 41760 32588 41812
rect 32640 41800 32646 41812
rect 32950 41800 32956 41812
rect 32640 41772 32956 41800
rect 32640 41760 32646 41772
rect 32950 41760 32956 41772
rect 33008 41760 33014 41812
rect 33410 41760 33416 41812
rect 33468 41800 33474 41812
rect 33689 41803 33747 41809
rect 33689 41800 33701 41803
rect 33468 41772 33701 41800
rect 33468 41760 33474 41772
rect 33689 41769 33701 41772
rect 33735 41769 33747 41803
rect 33689 41763 33747 41769
rect 35148 41803 35206 41809
rect 35148 41769 35160 41803
rect 35194 41800 35206 41803
rect 36538 41800 36544 41812
rect 35194 41772 36544 41800
rect 35194 41769 35206 41772
rect 35148 41763 35206 41769
rect 36538 41760 36544 41772
rect 36596 41760 36602 41812
rect 36633 41803 36691 41809
rect 36633 41769 36645 41803
rect 36679 41800 36691 41803
rect 36722 41800 36728 41812
rect 36679 41772 36728 41800
rect 36679 41769 36691 41772
rect 36633 41763 36691 41769
rect 36722 41760 36728 41772
rect 36780 41800 36786 41812
rect 36906 41800 36912 41812
rect 36780 41772 36912 41800
rect 36780 41760 36786 41772
rect 36906 41760 36912 41772
rect 36964 41760 36970 41812
rect 29178 41692 29184 41744
rect 29236 41732 29242 41744
rect 29236 41704 29868 41732
rect 29236 41692 29242 41704
rect 29454 41624 29460 41676
rect 29512 41664 29518 41676
rect 29733 41667 29791 41673
rect 29733 41664 29745 41667
rect 29512 41636 29745 41664
rect 29512 41624 29518 41636
rect 29733 41633 29745 41636
rect 29779 41633 29791 41667
rect 29840 41664 29868 41704
rect 30009 41667 30067 41673
rect 30009 41664 30021 41667
rect 29840 41636 30021 41664
rect 29733 41627 29791 41633
rect 30009 41633 30021 41636
rect 30055 41664 30067 41667
rect 30374 41664 30380 41676
rect 30055 41636 30380 41664
rect 30055 41633 30067 41636
rect 30009 41627 30067 41633
rect 30374 41624 30380 41636
rect 30432 41624 30438 41676
rect 30650 41624 30656 41676
rect 30708 41664 30714 41676
rect 30708 41636 31248 41664
rect 30708 41624 30714 41636
rect 28123 41568 28856 41596
rect 28123 41565 28135 41568
rect 28077 41559 28135 41565
rect 28994 41556 29000 41608
rect 29052 41556 29058 41608
rect 31220 41528 31248 41636
rect 31938 41624 31944 41676
rect 31996 41624 32002 41676
rect 32217 41667 32275 41673
rect 32217 41633 32229 41667
rect 32263 41664 32275 41667
rect 33870 41664 33876 41676
rect 32263 41636 33876 41664
rect 32263 41633 32275 41636
rect 32217 41627 32275 41633
rect 33870 41624 33876 41636
rect 33928 41664 33934 41676
rect 34330 41664 34336 41676
rect 33928 41636 34336 41664
rect 33928 41624 33934 41636
rect 34330 41624 34336 41636
rect 34388 41624 34394 41676
rect 34882 41624 34888 41676
rect 34940 41664 34946 41676
rect 35158 41664 35164 41676
rect 34940 41636 35164 41664
rect 34940 41624 34946 41636
rect 35158 41624 35164 41636
rect 35216 41624 35222 41676
rect 36556 41664 36584 41760
rect 36906 41664 36912 41676
rect 36556 41636 36912 41664
rect 36906 41624 36912 41636
rect 36964 41624 36970 41676
rect 49050 41556 49056 41608
rect 49108 41556 49114 41608
rect 31846 41528 31852 41540
rect 31220 41514 31852 41528
rect 31234 41500 31852 41514
rect 31846 41488 31852 41500
rect 31904 41488 31910 41540
rect 35250 41528 35256 41540
rect 33442 41500 35256 41528
rect 35250 41488 35256 41500
rect 35308 41488 35314 41540
rect 36446 41528 36452 41540
rect 36386 41500 36452 41528
rect 36446 41488 36452 41500
rect 36504 41488 36510 41540
rect 27111 41432 27752 41460
rect 27111 41429 27123 41432
rect 27065 41423 27123 41429
rect 27798 41420 27804 41472
rect 27856 41460 27862 41472
rect 27985 41463 28043 41469
rect 27985 41460 27997 41463
rect 27856 41432 27997 41460
rect 27856 41420 27862 41432
rect 27985 41429 27997 41432
rect 28031 41429 28043 41463
rect 27985 41423 28043 41429
rect 29546 41420 29552 41472
rect 29604 41460 29610 41472
rect 32306 41460 32312 41472
rect 29604 41432 32312 41460
rect 29604 41420 29610 41432
rect 32306 41420 32312 41432
rect 32364 41420 32370 41472
rect 36078 41420 36084 41472
rect 36136 41460 36142 41472
rect 36464 41460 36492 41488
rect 36136 41432 36492 41460
rect 36136 41420 36142 41432
rect 49234 41420 49240 41472
rect 49292 41420 49298 41472
rect 1104 41370 49864 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 27950 41370
rect 28002 41318 28014 41370
rect 28066 41318 28078 41370
rect 28130 41318 28142 41370
rect 28194 41318 28206 41370
rect 28258 41318 37950 41370
rect 38002 41318 38014 41370
rect 38066 41318 38078 41370
rect 38130 41318 38142 41370
rect 38194 41318 38206 41370
rect 38258 41318 47950 41370
rect 48002 41318 48014 41370
rect 48066 41318 48078 41370
rect 48130 41318 48142 41370
rect 48194 41318 48206 41370
rect 48258 41318 49864 41370
rect 1104 41296 49864 41318
rect 11054 41216 11060 41268
rect 11112 41256 11118 41268
rect 13265 41259 13323 41265
rect 13265 41256 13277 41259
rect 11112 41228 13277 41256
rect 11112 41216 11118 41228
rect 13265 41225 13277 41228
rect 13311 41225 13323 41259
rect 22094 41256 22100 41268
rect 13265 41219 13323 41225
rect 15948 41228 22100 41256
rect 12621 41191 12679 41197
rect 12621 41157 12633 41191
rect 12667 41188 12679 41191
rect 13173 41191 13231 41197
rect 13173 41188 13185 41191
rect 12667 41160 13185 41188
rect 12667 41157 12679 41160
rect 12621 41151 12679 41157
rect 13173 41157 13185 41160
rect 13219 41188 13231 41191
rect 15948 41188 15976 41228
rect 22094 41216 22100 41228
rect 22152 41216 22158 41268
rect 22373 41259 22431 41265
rect 22373 41225 22385 41259
rect 22419 41225 22431 41259
rect 22373 41219 22431 41225
rect 23569 41259 23627 41265
rect 23569 41225 23581 41259
rect 23615 41256 23627 41259
rect 23658 41256 23664 41268
rect 23615 41228 23664 41256
rect 23615 41225 23627 41228
rect 23569 41219 23627 41225
rect 13219 41160 15976 41188
rect 18233 41191 18291 41197
rect 13219 41157 13231 41160
rect 13173 41151 13231 41157
rect 18233 41157 18245 41191
rect 18279 41188 18291 41191
rect 18782 41188 18788 41200
rect 18279 41160 18788 41188
rect 18279 41157 18291 41160
rect 18233 41151 18291 41157
rect 18782 41148 18788 41160
rect 18840 41148 18846 41200
rect 19426 41188 19432 41200
rect 18892 41160 19432 41188
rect 1765 41123 1823 41129
rect 1765 41089 1777 41123
rect 1811 41120 1823 41123
rect 12250 41120 12256 41132
rect 1811 41092 12256 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 12250 41080 12256 41092
rect 12308 41080 12314 41132
rect 18892 41129 18920 41160
rect 19426 41148 19432 41160
rect 19484 41148 19490 41200
rect 20438 41188 20444 41200
rect 20378 41160 20444 41188
rect 20438 41148 20444 41160
rect 20496 41188 20502 41200
rect 21358 41188 21364 41200
rect 20496 41160 21364 41188
rect 20496 41148 20502 41160
rect 21358 41148 21364 41160
rect 21416 41188 21422 41200
rect 22002 41188 22008 41200
rect 21416 41160 22008 41188
rect 21416 41148 21422 41160
rect 22002 41148 22008 41160
rect 22060 41148 22066 41200
rect 22388 41188 22416 41219
rect 23658 41216 23664 41228
rect 23716 41216 23722 41268
rect 24762 41216 24768 41268
rect 24820 41216 24826 41268
rect 25222 41216 25228 41268
rect 25280 41216 25286 41268
rect 27706 41216 27712 41268
rect 27764 41216 27770 41268
rect 28077 41259 28135 41265
rect 28077 41225 28089 41259
rect 28123 41256 28135 41259
rect 28994 41256 29000 41268
rect 28123 41228 29000 41256
rect 28123 41225 28135 41228
rect 28077 41219 28135 41225
rect 28994 41216 29000 41228
rect 29052 41216 29058 41268
rect 29549 41259 29607 41265
rect 29549 41225 29561 41259
rect 29595 41256 29607 41259
rect 29730 41256 29736 41268
rect 29595 41228 29736 41256
rect 29595 41225 29607 41228
rect 29549 41219 29607 41225
rect 29730 41216 29736 41228
rect 29788 41216 29794 41268
rect 30653 41259 30711 41265
rect 30653 41256 30665 41259
rect 29840 41228 30665 41256
rect 23937 41191 23995 41197
rect 23937 41188 23949 41191
rect 22388 41160 23949 41188
rect 23937 41157 23949 41160
rect 23983 41157 23995 41191
rect 23937 41151 23995 41157
rect 28902 41148 28908 41200
rect 28960 41188 28966 41200
rect 29641 41191 29699 41197
rect 29641 41188 29653 41191
rect 28960 41160 29653 41188
rect 28960 41148 28966 41160
rect 29641 41157 29653 41160
rect 29687 41157 29699 41191
rect 29840 41188 29868 41228
rect 30653 41225 30665 41228
rect 30699 41225 30711 41259
rect 30653 41219 30711 41225
rect 30745 41259 30803 41265
rect 30745 41225 30757 41259
rect 30791 41256 30803 41259
rect 30834 41256 30840 41268
rect 30791 41228 30840 41256
rect 30791 41225 30803 41228
rect 30745 41219 30803 41225
rect 30834 41216 30840 41228
rect 30892 41216 30898 41268
rect 31573 41259 31631 41265
rect 31573 41225 31585 41259
rect 31619 41256 31631 41259
rect 32309 41259 32367 41265
rect 31619 41228 32168 41256
rect 31619 41225 31631 41228
rect 31573 41219 31631 41225
rect 29641 41151 29699 41157
rect 29748 41160 29868 41188
rect 15473 41123 15531 41129
rect 15473 41089 15485 41123
rect 15519 41089 15531 41123
rect 15473 41083 15531 41089
rect 18877 41123 18935 41129
rect 18877 41089 18889 41123
rect 18923 41089 18935 41123
rect 18877 41083 18935 41089
rect 1302 41012 1308 41064
rect 1360 41052 1366 41064
rect 2041 41055 2099 41061
rect 2041 41052 2053 41055
rect 1360 41024 2053 41052
rect 1360 41012 1366 41024
rect 2041 41021 2053 41024
rect 2087 41021 2099 41055
rect 2041 41015 2099 41021
rect 13814 40944 13820 40996
rect 13872 40984 13878 40996
rect 15102 40984 15108 40996
rect 13872 40956 15108 40984
rect 13872 40944 13878 40956
rect 15102 40944 15108 40956
rect 15160 40984 15166 40996
rect 15488 40984 15516 41083
rect 21082 41080 21088 41132
rect 21140 41120 21146 41132
rect 21269 41123 21327 41129
rect 21269 41120 21281 41123
rect 21140 41092 21281 41120
rect 21140 41080 21146 41092
rect 21269 41089 21281 41092
rect 21315 41089 21327 41123
rect 21269 41083 21327 41089
rect 22741 41123 22799 41129
rect 22741 41089 22753 41123
rect 22787 41120 22799 41123
rect 22787 41092 23520 41120
rect 22787 41089 22799 41092
rect 22741 41083 22799 41089
rect 18782 41012 18788 41064
rect 18840 41052 18846 41064
rect 19153 41055 19211 41061
rect 19153 41052 19165 41055
rect 18840 41024 19165 41052
rect 18840 41012 18846 41024
rect 19153 41021 19165 41024
rect 19199 41052 19211 41055
rect 19199 41024 22324 41052
rect 19199 41021 19211 41024
rect 19153 41015 19211 41021
rect 20990 40984 20996 40996
rect 15160 40956 15424 40984
rect 15488 40956 19012 40984
rect 15160 40944 15166 40956
rect 13538 40876 13544 40928
rect 13596 40916 13602 40928
rect 15289 40919 15347 40925
rect 15289 40916 15301 40919
rect 13596 40888 15301 40916
rect 13596 40876 13602 40888
rect 15289 40885 15301 40888
rect 15335 40885 15347 40919
rect 15396 40916 15424 40956
rect 18325 40919 18383 40925
rect 18325 40916 18337 40919
rect 15396 40888 18337 40916
rect 15289 40879 15347 40885
rect 18325 40885 18337 40888
rect 18371 40885 18383 40919
rect 18984 40916 19012 40956
rect 20548 40956 20996 40984
rect 20548 40916 20576 40956
rect 20990 40944 20996 40956
rect 21048 40944 21054 40996
rect 22296 40984 22324 41024
rect 22370 41012 22376 41064
rect 22428 41052 22434 41064
rect 22833 41055 22891 41061
rect 22833 41052 22845 41055
rect 22428 41024 22845 41052
rect 22428 41012 22434 41024
rect 22833 41021 22845 41024
rect 22879 41021 22891 41055
rect 22833 41015 22891 41021
rect 23017 41055 23075 41061
rect 23017 41021 23029 41055
rect 23063 41052 23075 41055
rect 23492 41052 23520 41092
rect 23566 41080 23572 41132
rect 23624 41120 23630 41132
rect 25133 41123 25191 41129
rect 25133 41120 25145 41123
rect 23624 41092 25145 41120
rect 23624 41080 23630 41092
rect 25133 41089 25145 41092
rect 25179 41089 25191 41123
rect 25133 41083 25191 41089
rect 25424 41092 28304 41120
rect 23934 41052 23940 41064
rect 23063 41024 23428 41052
rect 23492 41024 23940 41052
rect 23063 41021 23075 41024
rect 23017 41015 23075 41021
rect 23290 40984 23296 40996
rect 22296 40956 23296 40984
rect 23290 40944 23296 40956
rect 23348 40944 23354 40996
rect 23400 40984 23428 41024
rect 23934 41012 23940 41024
rect 23992 41012 23998 41064
rect 24026 41012 24032 41064
rect 24084 41012 24090 41064
rect 24210 41012 24216 41064
rect 24268 41012 24274 41064
rect 25424 41061 25452 41092
rect 25409 41055 25467 41061
rect 25409 41021 25421 41055
rect 25455 41021 25467 41055
rect 25409 41015 25467 41021
rect 27706 41012 27712 41064
rect 27764 41052 27770 41064
rect 28276 41061 28304 41092
rect 28350 41080 28356 41132
rect 28408 41120 28414 41132
rect 29748 41120 29776 41160
rect 28408 41092 29776 41120
rect 28408 41080 28414 41092
rect 28169 41055 28227 41061
rect 28169 41052 28181 41055
rect 27764 41024 28181 41052
rect 27764 41012 27770 41024
rect 28169 41021 28181 41024
rect 28215 41021 28227 41055
rect 28169 41015 28227 41021
rect 28261 41055 28319 41061
rect 28261 41021 28273 41055
rect 28307 41052 28319 41055
rect 28442 41052 28448 41064
rect 28307 41024 28448 41052
rect 28307 41021 28319 41024
rect 28261 41015 28319 41021
rect 28442 41012 28448 41024
rect 28500 41012 28506 41064
rect 28810 41012 28816 41064
rect 28868 41052 28874 41064
rect 29733 41055 29791 41061
rect 29733 41052 29745 41055
rect 28868 41024 29745 41052
rect 28868 41012 28874 41024
rect 29733 41021 29745 41024
rect 29779 41021 29791 41055
rect 29733 41015 29791 41021
rect 30834 41012 30840 41064
rect 30892 41012 30898 41064
rect 31018 41012 31024 41064
rect 31076 41052 31082 41064
rect 31386 41052 31392 41064
rect 31076 41024 31392 41052
rect 31076 41012 31082 41024
rect 31386 41012 31392 41024
rect 31444 41012 31450 41064
rect 24854 40984 24860 40996
rect 23400 40956 24860 40984
rect 24854 40944 24860 40956
rect 24912 40944 24918 40996
rect 25498 40944 25504 40996
rect 25556 40984 25562 40996
rect 28994 40984 29000 40996
rect 25556 40956 29000 40984
rect 25556 40944 25562 40956
rect 28994 40944 29000 40956
rect 29052 40944 29058 40996
rect 29178 40944 29184 40996
rect 29236 40944 29242 40996
rect 31588 40984 31616 41219
rect 32140 41188 32168 41228
rect 32309 41225 32321 41259
rect 32355 41256 32367 41259
rect 33410 41256 33416 41268
rect 32355 41228 33416 41256
rect 32355 41225 32367 41228
rect 32309 41219 32367 41225
rect 33410 41216 33416 41228
rect 33468 41216 33474 41268
rect 36538 41216 36544 41268
rect 36596 41216 36602 41268
rect 33965 41191 34023 41197
rect 32140 41160 32812 41188
rect 32490 41080 32496 41132
rect 32548 41120 32554 41132
rect 32784 41129 32812 41160
rect 33965 41157 33977 41191
rect 34011 41188 34023 41191
rect 34238 41188 34244 41200
rect 34011 41160 34244 41188
rect 34011 41157 34023 41160
rect 33965 41151 34023 41157
rect 34238 41148 34244 41160
rect 34296 41148 34302 41200
rect 35250 41188 35256 41200
rect 35190 41160 35256 41188
rect 35250 41148 35256 41160
rect 35308 41188 35314 41200
rect 36078 41188 36084 41200
rect 35308 41160 36084 41188
rect 35308 41148 35314 41160
rect 36078 41148 36084 41160
rect 36136 41148 36142 41200
rect 32677 41123 32735 41129
rect 32677 41120 32689 41123
rect 32548 41092 32689 41120
rect 32548 41080 32554 41092
rect 32677 41089 32689 41092
rect 32723 41089 32735 41123
rect 32677 41083 32735 41089
rect 32769 41123 32827 41129
rect 32769 41089 32781 41123
rect 32815 41120 32827 41123
rect 33318 41120 33324 41132
rect 32815 41092 33324 41120
rect 32815 41089 32827 41092
rect 32769 41083 32827 41089
rect 33318 41080 33324 41092
rect 33376 41080 33382 41132
rect 35434 41080 35440 41132
rect 35492 41120 35498 41132
rect 35713 41123 35771 41129
rect 35713 41120 35725 41123
rect 35492 41092 35725 41120
rect 35492 41080 35498 41092
rect 35713 41089 35725 41092
rect 35759 41089 35771 41123
rect 35713 41083 35771 41089
rect 36449 41123 36507 41129
rect 36449 41089 36461 41123
rect 36495 41120 36507 41123
rect 37182 41120 37188 41132
rect 36495 41092 37188 41120
rect 36495 41089 36507 41092
rect 36449 41083 36507 41089
rect 37182 41080 37188 41092
rect 37240 41080 37246 41132
rect 37274 41080 37280 41132
rect 37332 41120 37338 41132
rect 37461 41123 37519 41129
rect 37461 41120 37473 41123
rect 37332 41092 37473 41120
rect 37332 41080 37338 41092
rect 37461 41089 37473 41092
rect 37507 41089 37519 41123
rect 37461 41083 37519 41089
rect 38838 41080 38844 41132
rect 38896 41080 38902 41132
rect 49326 41080 49332 41132
rect 49384 41080 49390 41132
rect 32950 41012 32956 41064
rect 33008 41012 33014 41064
rect 33689 41055 33747 41061
rect 33689 41021 33701 41055
rect 33735 41052 33747 41055
rect 34514 41052 34520 41064
rect 33735 41024 34520 41052
rect 33735 41021 33747 41024
rect 33689 41015 33747 41021
rect 34514 41012 34520 41024
rect 34572 41012 34578 41064
rect 35986 41012 35992 41064
rect 36044 41052 36050 41064
rect 36633 41055 36691 41061
rect 36633 41052 36645 41055
rect 36044 41024 36645 41052
rect 36044 41012 36050 41024
rect 36633 41021 36645 41024
rect 36679 41021 36691 41055
rect 36633 41015 36691 41021
rect 36722 41012 36728 41064
rect 36780 41052 36786 41064
rect 37734 41052 37740 41064
rect 36780 41024 37740 41052
rect 36780 41012 36786 41024
rect 37734 41012 37740 41024
rect 37792 41012 37798 41064
rect 29748 40956 31616 40984
rect 29748 40928 29776 40956
rect 35066 40944 35072 40996
rect 35124 40984 35130 40996
rect 35124 40956 36216 40984
rect 35124 40944 35130 40956
rect 18984 40888 20576 40916
rect 18325 40879 18383 40885
rect 20622 40876 20628 40928
rect 20680 40876 20686 40928
rect 20898 40876 20904 40928
rect 20956 40916 20962 40928
rect 22370 40916 22376 40928
rect 20956 40888 22376 40916
rect 20956 40876 20962 40888
rect 22370 40876 22376 40888
rect 22428 40876 22434 40928
rect 28350 40876 28356 40928
rect 28408 40916 28414 40928
rect 28718 40916 28724 40928
rect 28408 40888 28724 40916
rect 28408 40876 28414 40888
rect 28718 40876 28724 40888
rect 28776 40876 28782 40928
rect 29730 40876 29736 40928
rect 29788 40876 29794 40928
rect 30285 40919 30343 40925
rect 30285 40885 30297 40919
rect 30331 40916 30343 40919
rect 31386 40916 31392 40928
rect 30331 40888 31392 40916
rect 30331 40885 30343 40888
rect 30285 40879 30343 40885
rect 31386 40876 31392 40888
rect 31444 40876 31450 40928
rect 32490 40876 32496 40928
rect 32548 40916 32554 40928
rect 33505 40919 33563 40925
rect 33505 40916 33517 40919
rect 32548 40888 33517 40916
rect 32548 40876 32554 40888
rect 33505 40885 33517 40888
rect 33551 40885 33563 40919
rect 33505 40879 33563 40885
rect 34606 40876 34612 40928
rect 34664 40916 34670 40928
rect 36081 40919 36139 40925
rect 36081 40916 36093 40919
rect 34664 40888 36093 40916
rect 34664 40876 34670 40888
rect 36081 40885 36093 40888
rect 36127 40885 36139 40919
rect 36188 40916 36216 40956
rect 38746 40916 38752 40928
rect 36188 40888 38752 40916
rect 36081 40879 36139 40885
rect 38746 40876 38752 40888
rect 38804 40876 38810 40928
rect 39206 40876 39212 40928
rect 39264 40876 39270 40928
rect 49142 40876 49148 40928
rect 49200 40876 49206 40928
rect 1104 40826 49864 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 32950 40826
rect 33002 40774 33014 40826
rect 33066 40774 33078 40826
rect 33130 40774 33142 40826
rect 33194 40774 33206 40826
rect 33258 40774 42950 40826
rect 43002 40774 43014 40826
rect 43066 40774 43078 40826
rect 43130 40774 43142 40826
rect 43194 40774 43206 40826
rect 43258 40774 49864 40826
rect 1104 40752 49864 40774
rect 12250 40672 12256 40724
rect 12308 40672 12314 40724
rect 17126 40672 17132 40724
rect 17184 40712 17190 40724
rect 17862 40712 17868 40724
rect 17184 40684 17868 40712
rect 17184 40672 17190 40684
rect 17862 40672 17868 40684
rect 17920 40672 17926 40724
rect 19429 40715 19487 40721
rect 19429 40681 19441 40715
rect 19475 40712 19487 40715
rect 19886 40712 19892 40724
rect 19475 40684 19892 40712
rect 19475 40681 19487 40684
rect 19429 40675 19487 40681
rect 19886 40672 19892 40684
rect 19944 40672 19950 40724
rect 20898 40712 20904 40724
rect 19996 40684 20904 40712
rect 9582 40604 9588 40656
rect 9640 40644 9646 40656
rect 13081 40647 13139 40653
rect 13081 40644 13093 40647
rect 9640 40616 13093 40644
rect 9640 40604 9646 40616
rect 13081 40613 13093 40616
rect 13127 40613 13139 40647
rect 19996 40644 20024 40684
rect 20898 40672 20904 40684
rect 20956 40672 20962 40724
rect 20990 40672 20996 40724
rect 21048 40712 21054 40724
rect 23566 40712 23572 40724
rect 21048 40684 23572 40712
rect 21048 40672 21054 40684
rect 23566 40672 23572 40684
rect 23624 40672 23630 40724
rect 24946 40672 24952 40724
rect 25004 40712 25010 40724
rect 26789 40715 26847 40721
rect 26789 40712 26801 40715
rect 25004 40684 26801 40712
rect 25004 40672 25010 40684
rect 26789 40681 26801 40684
rect 26835 40681 26847 40715
rect 26789 40675 26847 40681
rect 28077 40715 28135 40721
rect 28077 40681 28089 40715
rect 28123 40712 28135 40715
rect 29086 40712 29092 40724
rect 28123 40684 29092 40712
rect 28123 40681 28135 40684
rect 28077 40675 28135 40681
rect 29086 40672 29092 40684
rect 29144 40672 29150 40724
rect 35066 40712 35072 40724
rect 29196 40684 35072 40712
rect 13081 40607 13139 40613
rect 19904 40616 20024 40644
rect 16942 40576 16948 40588
rect 13280 40548 16948 40576
rect 13280 40517 13308 40548
rect 16942 40536 16948 40548
rect 17000 40536 17006 40588
rect 17126 40536 17132 40588
rect 17184 40576 17190 40588
rect 19904 40585 19932 40616
rect 22094 40604 22100 40656
rect 22152 40644 22158 40656
rect 25498 40644 25504 40656
rect 22152 40616 25504 40644
rect 22152 40604 22158 40616
rect 25498 40604 25504 40616
rect 25556 40604 25562 40656
rect 29196 40644 29224 40684
rect 35066 40672 35072 40684
rect 35124 40672 35130 40724
rect 37090 40712 37096 40724
rect 35268 40684 37096 40712
rect 28552 40616 29224 40644
rect 19889 40579 19947 40585
rect 17184 40548 19380 40576
rect 17184 40536 17190 40548
rect 13265 40511 13323 40517
rect 13265 40477 13277 40511
rect 13311 40477 13323 40511
rect 13265 40471 13323 40477
rect 15654 40468 15660 40520
rect 15712 40468 15718 40520
rect 15930 40468 15936 40520
rect 15988 40508 15994 40520
rect 16117 40511 16175 40517
rect 16117 40508 16129 40511
rect 15988 40480 16129 40508
rect 15988 40468 15994 40480
rect 16117 40477 16129 40480
rect 16163 40477 16175 40511
rect 16117 40471 16175 40477
rect 18417 40511 18475 40517
rect 18417 40477 18429 40511
rect 18463 40508 18475 40511
rect 19242 40508 19248 40520
rect 18463 40480 19248 40508
rect 18463 40477 18475 40480
rect 18417 40471 18475 40477
rect 19242 40468 19248 40480
rect 19300 40468 19306 40520
rect 12161 40443 12219 40449
rect 12161 40409 12173 40443
rect 12207 40440 12219 40443
rect 12207 40412 12434 40440
rect 12207 40409 12219 40412
rect 12161 40403 12219 40409
rect 12406 40372 12434 40412
rect 16022 40400 16028 40452
rect 16080 40440 16086 40452
rect 16393 40443 16451 40449
rect 16393 40440 16405 40443
rect 16080 40412 16405 40440
rect 16080 40400 16086 40412
rect 16393 40409 16405 40412
rect 16439 40440 16451 40443
rect 16666 40440 16672 40452
rect 16439 40412 16672 40440
rect 16439 40409 16451 40412
rect 16393 40403 16451 40409
rect 16666 40400 16672 40412
rect 16724 40400 16730 40452
rect 16850 40400 16856 40452
rect 16908 40400 16914 40452
rect 18601 40443 18659 40449
rect 18601 40409 18613 40443
rect 18647 40440 18659 40443
rect 18690 40440 18696 40452
rect 18647 40412 18696 40440
rect 18647 40409 18659 40412
rect 18601 40403 18659 40409
rect 18690 40400 18696 40412
rect 18748 40400 18754 40452
rect 18414 40372 18420 40384
rect 12406 40344 18420 40372
rect 18414 40332 18420 40344
rect 18472 40332 18478 40384
rect 19352 40372 19380 40548
rect 19889 40545 19901 40579
rect 19935 40545 19947 40579
rect 19889 40539 19947 40545
rect 19981 40579 20039 40585
rect 19981 40545 19993 40579
rect 20027 40576 20039 40579
rect 20070 40576 20076 40588
rect 20027 40548 20076 40576
rect 20027 40545 20039 40548
rect 19981 40539 20039 40545
rect 20070 40536 20076 40548
rect 20128 40536 20134 40588
rect 20530 40536 20536 40588
rect 20588 40576 20594 40588
rect 20625 40579 20683 40585
rect 20625 40576 20637 40579
rect 20588 40548 20637 40576
rect 20588 40536 20594 40548
rect 20625 40545 20637 40548
rect 20671 40545 20683 40579
rect 20625 40539 20683 40545
rect 22554 40536 22560 40588
rect 22612 40576 22618 40588
rect 22649 40579 22707 40585
rect 22649 40576 22661 40579
rect 22612 40548 22661 40576
rect 22612 40536 22618 40548
rect 22649 40545 22661 40548
rect 22695 40545 22707 40579
rect 22649 40539 22707 40545
rect 23842 40536 23848 40588
rect 23900 40536 23906 40588
rect 27338 40536 27344 40588
rect 27396 40536 27402 40588
rect 23753 40511 23811 40517
rect 23753 40477 23765 40511
rect 23799 40508 23811 40511
rect 24302 40508 24308 40520
rect 23799 40480 24308 40508
rect 23799 40477 23811 40480
rect 23753 40471 23811 40477
rect 24302 40468 24308 40480
rect 24360 40468 24366 40520
rect 25409 40511 25467 40517
rect 25409 40477 25421 40511
rect 25455 40508 25467 40511
rect 28445 40511 28503 40517
rect 28445 40508 28457 40511
rect 25455 40480 28457 40508
rect 25455 40477 25467 40480
rect 25409 40471 25467 40477
rect 28445 40477 28457 40480
rect 28491 40477 28503 40511
rect 28445 40471 28503 40477
rect 19797 40443 19855 40449
rect 19797 40409 19809 40443
rect 19843 40440 19855 40443
rect 20806 40440 20812 40452
rect 19843 40412 20812 40440
rect 19843 40409 19855 40412
rect 19797 40403 19855 40409
rect 20806 40400 20812 40412
rect 20864 40400 20870 40452
rect 20898 40400 20904 40452
rect 20956 40400 20962 40452
rect 21358 40400 21364 40452
rect 21416 40400 21422 40452
rect 26234 40400 26240 40452
rect 26292 40440 26298 40452
rect 27249 40443 27307 40449
rect 27249 40440 27261 40443
rect 26292 40412 27261 40440
rect 26292 40400 26298 40412
rect 27249 40409 27261 40412
rect 27295 40440 27307 40443
rect 28552 40440 28580 40616
rect 29822 40604 29828 40656
rect 29880 40644 29886 40656
rect 30929 40647 30987 40653
rect 29880 40616 30696 40644
rect 29880 40604 29886 40616
rect 28721 40579 28779 40585
rect 28721 40545 28733 40579
rect 28767 40576 28779 40579
rect 29362 40576 29368 40588
rect 28767 40548 29368 40576
rect 28767 40545 28779 40548
rect 28721 40539 28779 40545
rect 29362 40536 29368 40548
rect 29420 40536 29426 40588
rect 29638 40536 29644 40588
rect 29696 40576 29702 40588
rect 29696 40548 30236 40576
rect 29696 40536 29702 40548
rect 28626 40468 28632 40520
rect 28684 40508 28690 40520
rect 30101 40511 30159 40517
rect 30101 40508 30113 40511
rect 28684 40480 30113 40508
rect 28684 40468 28690 40480
rect 30101 40477 30113 40480
rect 30147 40477 30159 40511
rect 30208 40508 30236 40548
rect 30282 40536 30288 40588
rect 30340 40536 30346 40588
rect 30668 40576 30696 40616
rect 30929 40613 30941 40647
rect 30975 40644 30987 40647
rect 30975 40616 31754 40644
rect 30975 40613 30987 40616
rect 30929 40607 30987 40613
rect 31389 40579 31447 40585
rect 31389 40576 31401 40579
rect 30668 40548 31401 40576
rect 31389 40545 31401 40548
rect 31435 40545 31447 40579
rect 31389 40539 31447 40545
rect 31478 40536 31484 40588
rect 31536 40536 31542 40588
rect 31726 40576 31754 40616
rect 34330 40604 34336 40656
rect 34388 40644 34394 40656
rect 35268 40644 35296 40684
rect 37090 40672 37096 40684
rect 37148 40672 37154 40724
rect 37182 40672 37188 40724
rect 37240 40712 37246 40724
rect 38197 40715 38255 40721
rect 38197 40712 38209 40715
rect 37240 40684 38209 40712
rect 37240 40672 37246 40684
rect 38197 40681 38209 40684
rect 38243 40681 38255 40715
rect 47394 40712 47400 40724
rect 38197 40675 38255 40681
rect 41386 40684 47400 40712
rect 41386 40644 41414 40684
rect 47394 40672 47400 40684
rect 47452 40672 47458 40724
rect 34388 40616 35296 40644
rect 36832 40616 41414 40644
rect 34388 40604 34394 40616
rect 31726 40548 32812 40576
rect 32784 40520 32812 40548
rect 32858 40536 32864 40588
rect 32916 40576 32922 40588
rect 33137 40579 33195 40585
rect 33137 40576 33149 40579
rect 32916 40548 33149 40576
rect 32916 40536 32922 40548
rect 33137 40545 33149 40548
rect 33183 40545 33195 40579
rect 33137 40539 33195 40545
rect 33318 40536 33324 40588
rect 33376 40576 33382 40588
rect 36832 40576 36860 40616
rect 33376 40548 36860 40576
rect 33376 40536 33382 40548
rect 37090 40536 37096 40588
rect 37148 40576 37154 40588
rect 37185 40579 37243 40585
rect 37185 40576 37197 40579
rect 37148 40548 37197 40576
rect 37148 40536 37154 40548
rect 37185 40545 37197 40548
rect 37231 40545 37243 40579
rect 37185 40539 37243 40545
rect 37642 40536 37648 40588
rect 37700 40536 37706 40588
rect 37826 40536 37832 40588
rect 37884 40576 37890 40588
rect 38749 40579 38807 40585
rect 38749 40576 38761 40579
rect 37884 40548 38761 40576
rect 37884 40536 37890 40548
rect 38749 40545 38761 40548
rect 38795 40545 38807 40579
rect 38749 40539 38807 40545
rect 30558 40508 30564 40520
rect 30208 40480 30564 40508
rect 30101 40471 30159 40477
rect 30558 40468 30564 40480
rect 30616 40468 30622 40520
rect 30926 40468 30932 40520
rect 30984 40508 30990 40520
rect 31297 40511 31355 40517
rect 31297 40508 31309 40511
rect 30984 40480 31309 40508
rect 30984 40468 30990 40480
rect 31297 40477 31309 40480
rect 31343 40477 31355 40511
rect 31297 40471 31355 40477
rect 32398 40468 32404 40520
rect 32456 40468 32462 40520
rect 32766 40468 32772 40520
rect 32824 40468 32830 40520
rect 34514 40468 34520 40520
rect 34572 40508 34578 40520
rect 35158 40508 35164 40520
rect 34572 40480 35164 40508
rect 34572 40468 34578 40480
rect 35158 40468 35164 40480
rect 35216 40468 35222 40520
rect 38565 40511 38623 40517
rect 38565 40477 38577 40511
rect 38611 40508 38623 40511
rect 49142 40508 49148 40520
rect 38611 40480 49148 40508
rect 38611 40477 38623 40480
rect 38565 40471 38623 40477
rect 49142 40468 49148 40480
rect 49200 40468 49206 40520
rect 33686 40440 33692 40452
rect 27295 40412 28580 40440
rect 29748 40412 33692 40440
rect 27295 40409 27307 40412
rect 27249 40403 27307 40409
rect 20990 40372 20996 40384
rect 19352 40344 20996 40372
rect 20990 40332 20996 40344
rect 21048 40332 21054 40384
rect 22462 40332 22468 40384
rect 22520 40372 22526 40384
rect 23293 40375 23351 40381
rect 23293 40372 23305 40375
rect 22520 40344 23305 40372
rect 22520 40332 22526 40344
rect 23293 40341 23305 40344
rect 23339 40341 23351 40375
rect 23293 40335 23351 40341
rect 23661 40375 23719 40381
rect 23661 40341 23673 40375
rect 23707 40372 23719 40375
rect 25866 40372 25872 40384
rect 23707 40344 25872 40372
rect 23707 40341 23719 40344
rect 23661 40335 23719 40341
rect 25866 40332 25872 40344
rect 25924 40332 25930 40384
rect 26418 40332 26424 40384
rect 26476 40372 26482 40384
rect 27157 40375 27215 40381
rect 27157 40372 27169 40375
rect 26476 40344 27169 40372
rect 26476 40332 26482 40344
rect 27157 40341 27169 40344
rect 27203 40341 27215 40375
rect 27157 40335 27215 40341
rect 28537 40375 28595 40381
rect 28537 40341 28549 40375
rect 28583 40372 28595 40375
rect 28718 40372 28724 40384
rect 28583 40344 28724 40372
rect 28583 40341 28595 40344
rect 28537 40335 28595 40341
rect 28718 40332 28724 40344
rect 28776 40332 28782 40384
rect 29748 40381 29776 40412
rect 33686 40400 33692 40412
rect 33744 40400 33750 40452
rect 35437 40443 35495 40449
rect 35437 40409 35449 40443
rect 35483 40409 35495 40443
rect 35437 40403 35495 40409
rect 29733 40375 29791 40381
rect 29733 40341 29745 40375
rect 29779 40341 29791 40375
rect 29733 40335 29791 40341
rect 30098 40332 30104 40384
rect 30156 40372 30162 40384
rect 30193 40375 30251 40381
rect 30193 40372 30205 40375
rect 30156 40344 30205 40372
rect 30156 40332 30162 40344
rect 30193 40341 30205 40344
rect 30239 40341 30251 40375
rect 30193 40335 30251 40341
rect 31754 40332 31760 40384
rect 31812 40372 31818 40384
rect 33962 40372 33968 40384
rect 31812 40344 33968 40372
rect 31812 40332 31818 40344
rect 33962 40332 33968 40344
rect 34020 40332 34026 40384
rect 35452 40372 35480 40403
rect 36078 40400 36084 40452
rect 36136 40400 36142 40452
rect 39206 40440 39212 40452
rect 37568 40412 39212 40440
rect 37568 40372 37596 40412
rect 39206 40400 39212 40412
rect 39264 40400 39270 40452
rect 47210 40440 47216 40452
rect 41386 40412 47216 40440
rect 35452 40344 37596 40372
rect 37642 40332 37648 40384
rect 37700 40372 37706 40384
rect 38657 40375 38715 40381
rect 38657 40372 38669 40375
rect 37700 40344 38669 40372
rect 37700 40332 37706 40344
rect 38657 40341 38669 40344
rect 38703 40372 38715 40375
rect 41386 40372 41414 40412
rect 47210 40400 47216 40412
rect 47268 40400 47274 40452
rect 38703 40344 41414 40372
rect 38703 40341 38715 40344
rect 38657 40335 38715 40341
rect 1104 40282 49864 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 27950 40282
rect 28002 40230 28014 40282
rect 28066 40230 28078 40282
rect 28130 40230 28142 40282
rect 28194 40230 28206 40282
rect 28258 40230 37950 40282
rect 38002 40230 38014 40282
rect 38066 40230 38078 40282
rect 38130 40230 38142 40282
rect 38194 40230 38206 40282
rect 38258 40230 47950 40282
rect 48002 40230 48014 40282
rect 48066 40230 48078 40282
rect 48130 40230 48142 40282
rect 48194 40230 48206 40282
rect 48258 40230 49864 40282
rect 1104 40208 49864 40230
rect 12802 40128 12808 40180
rect 12860 40168 12866 40180
rect 14277 40171 14335 40177
rect 14277 40168 14289 40171
rect 12860 40140 14289 40168
rect 12860 40128 12866 40140
rect 14277 40137 14289 40140
rect 14323 40137 14335 40171
rect 14277 40131 14335 40137
rect 17310 40128 17316 40180
rect 17368 40168 17374 40180
rect 18141 40171 18199 40177
rect 18141 40168 18153 40171
rect 17368 40140 18153 40168
rect 17368 40128 17374 40140
rect 18141 40137 18153 40140
rect 18187 40137 18199 40171
rect 18141 40131 18199 40137
rect 18509 40171 18567 40177
rect 18509 40137 18521 40171
rect 18555 40168 18567 40171
rect 18874 40168 18880 40180
rect 18555 40140 18880 40168
rect 18555 40137 18567 40140
rect 18509 40131 18567 40137
rect 18874 40128 18880 40140
rect 18932 40128 18938 40180
rect 20622 40168 20628 40180
rect 19904 40140 20628 40168
rect 8386 40100 8392 40112
rect 1780 40072 8392 40100
rect 1780 40041 1808 40072
rect 8386 40060 8392 40072
rect 8444 40060 8450 40112
rect 9306 40060 9312 40112
rect 9364 40100 9370 40112
rect 9582 40100 9588 40112
rect 9364 40072 9588 40100
rect 9364 40060 9370 40072
rect 9582 40060 9588 40072
rect 9640 40060 9646 40112
rect 16850 40060 16856 40112
rect 16908 40100 16914 40112
rect 17678 40100 17684 40112
rect 16908 40072 17684 40100
rect 16908 40060 16914 40072
rect 17678 40060 17684 40072
rect 17736 40060 17742 40112
rect 19518 40060 19524 40112
rect 19576 40100 19582 40112
rect 19904 40109 19932 40140
rect 20622 40128 20628 40140
rect 20680 40128 20686 40180
rect 20806 40128 20812 40180
rect 20864 40168 20870 40180
rect 21361 40171 21419 40177
rect 20864 40140 21312 40168
rect 20864 40128 20870 40140
rect 19889 40103 19947 40109
rect 19889 40100 19901 40103
rect 19576 40072 19901 40100
rect 19576 40060 19582 40072
rect 19889 40069 19901 40072
rect 19935 40069 19947 40103
rect 21284 40100 21312 40140
rect 21361 40137 21373 40171
rect 21407 40168 21419 40171
rect 21818 40168 21824 40180
rect 21407 40140 21824 40168
rect 21407 40137 21419 40140
rect 21361 40131 21419 40137
rect 21818 40128 21824 40140
rect 21876 40128 21882 40180
rect 22278 40128 22284 40180
rect 22336 40128 22342 40180
rect 23750 40128 23756 40180
rect 23808 40168 23814 40180
rect 26329 40171 26387 40177
rect 26329 40168 26341 40171
rect 23808 40140 26341 40168
rect 23808 40128 23814 40140
rect 26329 40137 26341 40140
rect 26375 40137 26387 40171
rect 26329 40131 26387 40137
rect 26694 40128 26700 40180
rect 26752 40168 26758 40180
rect 27525 40171 27583 40177
rect 27525 40168 27537 40171
rect 26752 40140 27537 40168
rect 26752 40128 26758 40140
rect 27525 40137 27537 40140
rect 27571 40168 27583 40171
rect 27798 40168 27804 40180
rect 27571 40140 27804 40168
rect 27571 40137 27583 40140
rect 27525 40131 27583 40137
rect 27798 40128 27804 40140
rect 27856 40128 27862 40180
rect 29730 40128 29736 40180
rect 29788 40168 29794 40180
rect 30285 40171 30343 40177
rect 30285 40168 30297 40171
rect 29788 40140 30297 40168
rect 29788 40128 29794 40140
rect 30285 40137 30297 40140
rect 30331 40168 30343 40171
rect 31478 40168 31484 40180
rect 30331 40140 31484 40168
rect 30331 40137 30343 40140
rect 30285 40131 30343 40137
rect 31478 40128 31484 40140
rect 31536 40128 31542 40180
rect 34422 40168 34428 40180
rect 31864 40140 34428 40168
rect 22462 40100 22468 40112
rect 21284 40072 22468 40100
rect 19889 40063 19947 40069
rect 22462 40060 22468 40072
rect 22520 40060 22526 40112
rect 22649 40103 22707 40109
rect 22649 40069 22661 40103
rect 22695 40100 22707 40103
rect 22830 40100 22836 40112
rect 22695 40072 22836 40100
rect 22695 40069 22707 40072
rect 22649 40063 22707 40069
rect 22830 40060 22836 40072
rect 22888 40060 22894 40112
rect 23845 40103 23903 40109
rect 23845 40069 23857 40103
rect 23891 40100 23903 40103
rect 24946 40100 24952 40112
rect 23891 40072 24952 40100
rect 23891 40069 23903 40072
rect 23845 40063 23903 40069
rect 24946 40060 24952 40072
rect 25004 40060 25010 40112
rect 25498 40060 25504 40112
rect 25556 40060 25562 40112
rect 27430 40060 27436 40112
rect 27488 40100 27494 40112
rect 30650 40100 30656 40112
rect 27488 40072 27844 40100
rect 30038 40072 30656 40100
rect 27488 40060 27494 40072
rect 1765 40035 1823 40041
rect 1765 40001 1777 40035
rect 1811 40001 1823 40035
rect 1765 39995 1823 40001
rect 14642 39992 14648 40044
rect 14700 39992 14706 40044
rect 14737 40035 14795 40041
rect 14737 40001 14749 40035
rect 14783 40032 14795 40035
rect 15470 40032 15476 40044
rect 14783 40004 15476 40032
rect 14783 40001 14795 40004
rect 14737 39995 14795 40001
rect 15470 39992 15476 40004
rect 15528 39992 15534 40044
rect 15565 40035 15623 40041
rect 15565 40001 15577 40035
rect 15611 40032 15623 40035
rect 16117 40035 16175 40041
rect 16117 40032 16129 40035
rect 15611 40004 16129 40032
rect 15611 40001 15623 40004
rect 15565 39995 15623 40001
rect 16117 40001 16129 40004
rect 16163 40032 16175 40035
rect 16298 40032 16304 40044
rect 16163 40004 16304 40032
rect 16163 40001 16175 40004
rect 16117 39995 16175 40001
rect 16298 39992 16304 40004
rect 16356 39992 16362 40044
rect 19426 40032 19432 40044
rect 18616 40004 19432 40032
rect 2038 39924 2044 39976
rect 2096 39924 2102 39976
rect 14918 39924 14924 39976
rect 14976 39924 14982 39976
rect 18616 39973 18644 40004
rect 19426 39992 19432 40004
rect 19484 39992 19490 40044
rect 20990 39992 20996 40044
rect 21048 40032 21054 40044
rect 21358 40032 21364 40044
rect 21048 40004 21364 40032
rect 21048 39992 21054 40004
rect 21358 39992 21364 40004
rect 21416 39992 21422 40044
rect 21726 39992 21732 40044
rect 21784 40032 21790 40044
rect 23937 40035 23995 40041
rect 21784 40004 22508 40032
rect 21784 39992 21790 40004
rect 18601 39967 18659 39973
rect 18601 39964 18613 39967
rect 17604 39936 18613 39964
rect 3326 39856 3332 39908
rect 3384 39896 3390 39908
rect 17604 39905 17632 39936
rect 18601 39933 18613 39936
rect 18647 39933 18659 39967
rect 18601 39927 18659 39933
rect 18782 39924 18788 39976
rect 18840 39924 18846 39976
rect 19610 39924 19616 39976
rect 19668 39924 19674 39976
rect 22186 39964 22192 39976
rect 19720 39936 22192 39964
rect 17589 39899 17647 39905
rect 17589 39896 17601 39899
rect 3384 39868 17601 39896
rect 3384 39856 3390 39868
rect 17589 39865 17601 39868
rect 17635 39865 17647 39899
rect 17589 39859 17647 39865
rect 17678 39856 17684 39908
rect 17736 39896 17742 39908
rect 19720 39896 19748 39936
rect 22186 39924 22192 39936
rect 22244 39924 22250 39976
rect 17736 39868 19748 39896
rect 22480 39896 22508 40004
rect 23937 40001 23949 40035
rect 23983 40032 23995 40035
rect 23983 40004 24348 40032
rect 23983 40001 23995 40004
rect 23937 39995 23995 40001
rect 22554 39924 22560 39976
rect 22612 39964 22618 39976
rect 22741 39967 22799 39973
rect 22741 39964 22753 39967
rect 22612 39936 22753 39964
rect 22612 39924 22618 39936
rect 22741 39933 22753 39936
rect 22787 39933 22799 39967
rect 22741 39927 22799 39933
rect 22833 39967 22891 39973
rect 22833 39933 22845 39967
rect 22879 39933 22891 39967
rect 22833 39927 22891 39933
rect 24029 39967 24087 39973
rect 24029 39933 24041 39967
rect 24075 39933 24087 39967
rect 24320 39964 24348 40004
rect 24578 39992 24584 40044
rect 24636 39992 24642 40044
rect 24857 39967 24915 39973
rect 24320 39936 24716 39964
rect 24029 39927 24087 39933
rect 22848 39896 22876 39927
rect 22480 39868 22876 39896
rect 17736 39856 17742 39868
rect 23750 39856 23756 39908
rect 23808 39896 23814 39908
rect 24044 39896 24072 39927
rect 23808 39868 24072 39896
rect 23808 39856 23814 39868
rect 7558 39788 7564 39840
rect 7616 39828 7622 39840
rect 12710 39828 12716 39840
rect 7616 39800 12716 39828
rect 7616 39788 7622 39800
rect 12710 39788 12716 39800
rect 12768 39788 12774 39840
rect 14366 39788 14372 39840
rect 14424 39828 14430 39840
rect 16209 39831 16267 39837
rect 16209 39828 16221 39831
rect 14424 39800 16221 39828
rect 14424 39788 14430 39800
rect 16209 39797 16221 39800
rect 16255 39797 16267 39831
rect 16209 39791 16267 39797
rect 22738 39788 22744 39840
rect 22796 39828 22802 39840
rect 23477 39831 23535 39837
rect 23477 39828 23489 39831
rect 22796 39800 23489 39828
rect 22796 39788 22802 39800
rect 23477 39797 23489 39800
rect 23523 39797 23535 39831
rect 23477 39791 23535 39797
rect 23934 39788 23940 39840
rect 23992 39828 23998 39840
rect 24486 39828 24492 39840
rect 23992 39800 24492 39828
rect 23992 39788 23998 39800
rect 24486 39788 24492 39800
rect 24544 39788 24550 39840
rect 24688 39828 24716 39936
rect 24857 39933 24869 39967
rect 24903 39964 24915 39967
rect 26878 39964 26884 39976
rect 24903 39936 26884 39964
rect 24903 39933 24915 39936
rect 24857 39927 24915 39933
rect 26878 39924 26884 39936
rect 26936 39924 26942 39976
rect 27338 39924 27344 39976
rect 27396 39964 27402 39976
rect 27617 39967 27675 39973
rect 27617 39964 27629 39967
rect 27396 39936 27629 39964
rect 27396 39924 27402 39936
rect 27617 39933 27629 39936
rect 27663 39933 27675 39967
rect 27617 39927 27675 39933
rect 27709 39967 27767 39973
rect 27709 39933 27721 39967
rect 27755 39933 27767 39967
rect 27816 39964 27844 40072
rect 30650 40060 30656 40072
rect 30708 40060 30714 40112
rect 31389 40103 31447 40109
rect 31389 40069 31401 40103
rect 31435 40100 31447 40103
rect 31754 40100 31760 40112
rect 31435 40072 31760 40100
rect 31435 40069 31447 40072
rect 31389 40063 31447 40069
rect 31754 40060 31760 40072
rect 31812 40060 31818 40112
rect 31110 39992 31116 40044
rect 31168 40032 31174 40044
rect 31481 40035 31539 40041
rect 31481 40032 31493 40035
rect 31168 40004 31493 40032
rect 31168 39992 31174 40004
rect 31481 40001 31493 40004
rect 31527 40001 31539 40035
rect 31481 39995 31539 40001
rect 28537 39967 28595 39973
rect 28537 39964 28549 39967
rect 27816 39936 28549 39964
rect 27709 39927 27767 39933
rect 28537 39933 28549 39936
rect 28583 39933 28595 39967
rect 28537 39927 28595 39933
rect 28813 39967 28871 39973
rect 28813 39933 28825 39967
rect 28859 39964 28871 39967
rect 30190 39964 30196 39976
rect 28859 39936 30196 39964
rect 28859 39933 28871 39936
rect 28813 39927 28871 39933
rect 26510 39896 26516 39908
rect 25884 39868 26516 39896
rect 25884 39828 25912 39868
rect 26510 39856 26516 39868
rect 26568 39856 26574 39908
rect 27724 39896 27752 39927
rect 30190 39924 30196 39936
rect 30248 39924 30254 39976
rect 31570 39924 31576 39976
rect 31628 39924 31634 39976
rect 26620 39868 27752 39896
rect 31021 39899 31079 39905
rect 24688 39800 25912 39828
rect 25958 39788 25964 39840
rect 26016 39828 26022 39840
rect 26620 39828 26648 39868
rect 31021 39865 31033 39899
rect 31067 39896 31079 39899
rect 31864 39896 31892 40140
rect 34422 40128 34428 40140
rect 34480 40128 34486 40180
rect 35434 40128 35440 40180
rect 35492 40168 35498 40180
rect 36170 40168 36176 40180
rect 35492 40140 36176 40168
rect 35492 40128 35498 40140
rect 36170 40128 36176 40140
rect 36228 40168 36234 40180
rect 36265 40171 36323 40177
rect 36265 40168 36277 40171
rect 36228 40140 36277 40168
rect 36228 40128 36234 40140
rect 36265 40137 36277 40140
rect 36311 40137 36323 40171
rect 36265 40131 36323 40137
rect 38657 40171 38715 40177
rect 38657 40137 38669 40171
rect 38703 40168 38715 40171
rect 38746 40168 38752 40180
rect 38703 40140 38752 40168
rect 38703 40137 38715 40140
rect 38657 40131 38715 40137
rect 38746 40128 38752 40140
rect 38804 40128 38810 40180
rect 32858 40100 32864 40112
rect 32324 40072 32864 40100
rect 32324 40044 32352 40072
rect 32858 40060 32864 40072
rect 32916 40060 32922 40112
rect 33870 40100 33876 40112
rect 33810 40072 33876 40100
rect 33870 40060 33876 40072
rect 33928 40100 33934 40112
rect 35250 40100 35256 40112
rect 33928 40072 35256 40100
rect 33928 40060 33934 40072
rect 35250 40060 35256 40072
rect 35308 40060 35314 40112
rect 39025 40103 39083 40109
rect 39025 40069 39037 40103
rect 39071 40069 39083 40103
rect 39025 40063 39083 40069
rect 32306 39992 32312 40044
rect 32364 39992 32370 40044
rect 34514 39992 34520 40044
rect 34572 39992 34578 40044
rect 32585 39967 32643 39973
rect 32585 39933 32597 39967
rect 32631 39964 32643 39967
rect 33594 39964 33600 39976
rect 32631 39936 33600 39964
rect 32631 39933 32643 39936
rect 32585 39927 32643 39933
rect 33594 39924 33600 39936
rect 33652 39964 33658 39976
rect 33870 39964 33876 39976
rect 33652 39936 33876 39964
rect 33652 39924 33658 39936
rect 33870 39924 33876 39936
rect 33928 39924 33934 39976
rect 34422 39924 34428 39976
rect 34480 39964 34486 39976
rect 34793 39967 34851 39973
rect 34793 39964 34805 39967
rect 34480 39936 34805 39964
rect 34480 39924 34486 39936
rect 34793 39933 34805 39936
rect 34839 39964 34851 39967
rect 35342 39964 35348 39976
rect 34839 39936 35348 39964
rect 34839 39933 34851 39936
rect 34793 39927 34851 39933
rect 35342 39924 35348 39936
rect 35400 39924 35406 39976
rect 39040 39964 39068 40063
rect 39114 39992 39120 40044
rect 39172 39992 39178 40044
rect 49050 39992 49056 40044
rect 49108 39992 49114 40044
rect 38120 39936 39068 39964
rect 38120 39905 38148 39936
rect 38105 39899 38163 39905
rect 38105 39896 38117 39899
rect 31067 39868 31892 39896
rect 33980 39868 34652 39896
rect 31067 39865 31079 39868
rect 31021 39859 31079 39865
rect 26016 39800 26648 39828
rect 26016 39788 26022 39800
rect 27154 39788 27160 39840
rect 27212 39788 27218 39840
rect 27798 39788 27804 39840
rect 27856 39828 27862 39840
rect 28902 39828 28908 39840
rect 27856 39800 28908 39828
rect 27856 39788 27862 39800
rect 28902 39788 28908 39800
rect 28960 39828 28966 39840
rect 33980 39828 34008 39868
rect 28960 39800 34008 39828
rect 28960 39788 28966 39800
rect 34054 39788 34060 39840
rect 34112 39788 34118 39840
rect 34624 39828 34652 39868
rect 37476 39868 38117 39896
rect 37476 39828 37504 39868
rect 38105 39865 38117 39868
rect 38151 39865 38163 39899
rect 38105 39859 38163 39865
rect 34624 39800 37504 39828
rect 37550 39788 37556 39840
rect 37608 39828 37614 39840
rect 38470 39828 38476 39840
rect 37608 39800 38476 39828
rect 37608 39788 37614 39800
rect 38470 39788 38476 39800
rect 38528 39788 38534 39840
rect 39040 39828 39068 39936
rect 39301 39967 39359 39973
rect 39301 39933 39313 39967
rect 39347 39964 39359 39967
rect 39390 39964 39396 39976
rect 39347 39936 39396 39964
rect 39347 39933 39359 39936
rect 39301 39927 39359 39933
rect 39390 39924 39396 39936
rect 39448 39924 39454 39976
rect 49237 39831 49295 39837
rect 49237 39828 49249 39831
rect 39040 39800 49249 39828
rect 49237 39797 49249 39800
rect 49283 39797 49295 39831
rect 49237 39791 49295 39797
rect 1104 39738 49864 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 32950 39738
rect 33002 39686 33014 39738
rect 33066 39686 33078 39738
rect 33130 39686 33142 39738
rect 33194 39686 33206 39738
rect 33258 39686 42950 39738
rect 43002 39686 43014 39738
rect 43066 39686 43078 39738
rect 43130 39686 43142 39738
rect 43194 39686 43206 39738
rect 43258 39686 49864 39738
rect 1104 39664 49864 39686
rect 1670 39584 1676 39636
rect 1728 39624 1734 39636
rect 7558 39624 7564 39636
rect 1728 39596 7564 39624
rect 1728 39584 1734 39596
rect 7558 39584 7564 39596
rect 7616 39584 7622 39636
rect 13357 39627 13415 39633
rect 13357 39624 13369 39627
rect 7668 39596 13369 39624
rect 7668 39488 7696 39596
rect 13357 39593 13369 39596
rect 13403 39593 13415 39627
rect 13357 39587 13415 39593
rect 14642 39584 14648 39636
rect 14700 39624 14706 39636
rect 14921 39627 14979 39633
rect 14921 39624 14933 39627
rect 14700 39596 14933 39624
rect 14700 39584 14706 39596
rect 14921 39593 14933 39596
rect 14967 39593 14979 39627
rect 14921 39587 14979 39593
rect 16666 39584 16672 39636
rect 16724 39624 16730 39636
rect 17405 39627 17463 39633
rect 17405 39624 17417 39627
rect 16724 39596 17417 39624
rect 16724 39584 16730 39596
rect 17405 39593 17417 39596
rect 17451 39593 17463 39627
rect 17405 39587 17463 39593
rect 17770 39584 17776 39636
rect 17828 39624 17834 39636
rect 18141 39627 18199 39633
rect 18141 39624 18153 39627
rect 17828 39596 18153 39624
rect 17828 39584 17834 39596
rect 18141 39593 18153 39596
rect 18187 39593 18199 39627
rect 18141 39587 18199 39593
rect 18248 39596 21680 39624
rect 1780 39460 7696 39488
rect 10689 39491 10747 39497
rect 1780 39429 1808 39460
rect 10689 39457 10701 39491
rect 10735 39488 10747 39491
rect 14458 39488 14464 39500
rect 10735 39460 14464 39488
rect 10735 39457 10747 39460
rect 10689 39451 10747 39457
rect 14458 39448 14464 39460
rect 14516 39488 14522 39500
rect 15657 39491 15715 39497
rect 15657 39488 15669 39491
rect 14516 39460 15669 39488
rect 14516 39448 14522 39460
rect 15657 39457 15669 39460
rect 15703 39488 15715 39491
rect 15930 39488 15936 39500
rect 15703 39460 15936 39488
rect 15703 39457 15715 39460
rect 15657 39451 15715 39457
rect 15930 39448 15936 39460
rect 15988 39448 15994 39500
rect 16298 39448 16304 39500
rect 16356 39488 16362 39500
rect 18248 39488 18276 39596
rect 21542 39556 21548 39568
rect 20364 39528 21548 39556
rect 20364 39497 20392 39528
rect 21542 39516 21548 39528
rect 21600 39516 21606 39568
rect 21652 39556 21680 39596
rect 21726 39584 21732 39636
rect 21784 39624 21790 39636
rect 22462 39624 22468 39636
rect 21784 39596 22468 39624
rect 21784 39584 21790 39596
rect 22462 39584 22468 39596
rect 22520 39584 22526 39636
rect 24394 39624 24400 39636
rect 22940 39596 24400 39624
rect 22940 39556 22968 39596
rect 24394 39584 24400 39596
rect 24452 39584 24458 39636
rect 24581 39627 24639 39633
rect 24581 39593 24593 39627
rect 24627 39624 24639 39627
rect 25038 39624 25044 39636
rect 24627 39596 25044 39624
rect 24627 39593 24639 39596
rect 24581 39587 24639 39593
rect 25038 39584 25044 39596
rect 25096 39584 25102 39636
rect 25866 39584 25872 39636
rect 25924 39584 25930 39636
rect 26881 39627 26939 39633
rect 26881 39593 26893 39627
rect 26927 39624 26939 39627
rect 28626 39624 28632 39636
rect 26927 39596 28632 39624
rect 26927 39593 26939 39596
rect 26881 39587 26939 39593
rect 28626 39584 28632 39596
rect 28684 39584 28690 39636
rect 29086 39584 29092 39636
rect 29144 39624 29150 39636
rect 30006 39624 30012 39636
rect 29144 39596 30012 39624
rect 29144 39584 29150 39596
rect 30006 39584 30012 39596
rect 30064 39584 30070 39636
rect 31560 39627 31618 39633
rect 31560 39593 31572 39627
rect 31606 39624 31618 39627
rect 31754 39624 31760 39636
rect 31606 39596 31760 39624
rect 31606 39593 31618 39596
rect 31560 39587 31618 39593
rect 31754 39584 31760 39596
rect 31812 39584 31818 39636
rect 31938 39584 31944 39636
rect 31996 39624 32002 39636
rect 33045 39627 33103 39633
rect 33045 39624 33057 39627
rect 31996 39596 33057 39624
rect 31996 39584 32002 39596
rect 33045 39593 33057 39596
rect 33091 39593 33103 39627
rect 33045 39587 33103 39593
rect 34054 39584 34060 39636
rect 34112 39624 34118 39636
rect 34112 39596 36308 39624
rect 34112 39584 34118 39596
rect 21652 39528 22968 39556
rect 23014 39516 23020 39568
rect 23072 39516 23078 39568
rect 29733 39559 29791 39565
rect 29733 39525 29745 39559
rect 29779 39525 29791 39559
rect 29733 39519 29791 39525
rect 16356 39460 18276 39488
rect 18693 39491 18751 39497
rect 16356 39448 16362 39460
rect 18693 39457 18705 39491
rect 18739 39457 18751 39491
rect 18693 39451 18751 39457
rect 20349 39491 20407 39497
rect 20349 39457 20361 39491
rect 20395 39457 20407 39491
rect 20349 39451 20407 39457
rect 1765 39423 1823 39429
rect 1765 39389 1777 39423
rect 1811 39389 1823 39423
rect 1765 39383 1823 39389
rect 12710 39380 12716 39432
rect 12768 39420 12774 39432
rect 13630 39420 13636 39432
rect 12768 39392 13636 39420
rect 12768 39380 12774 39392
rect 13630 39380 13636 39392
rect 13688 39380 13694 39432
rect 17862 39380 17868 39432
rect 17920 39420 17926 39432
rect 18708 39420 18736 39451
rect 20898 39448 20904 39500
rect 20956 39488 20962 39500
rect 21450 39488 21456 39500
rect 20956 39460 21456 39488
rect 20956 39448 20962 39460
rect 21450 39448 21456 39460
rect 21508 39448 21514 39500
rect 22646 39448 22652 39500
rect 22704 39488 22710 39500
rect 23569 39491 23627 39497
rect 23569 39488 23581 39491
rect 22704 39460 23581 39488
rect 22704 39448 22710 39460
rect 23569 39457 23581 39460
rect 23615 39457 23627 39491
rect 23569 39451 23627 39457
rect 25130 39448 25136 39500
rect 25188 39448 25194 39500
rect 26513 39491 26571 39497
rect 26513 39457 26525 39491
rect 26559 39488 26571 39491
rect 26878 39488 26884 39500
rect 26559 39460 26884 39488
rect 26559 39457 26571 39460
rect 26513 39451 26571 39457
rect 26878 39448 26884 39460
rect 26936 39448 26942 39500
rect 27062 39448 27068 39500
rect 27120 39488 27126 39500
rect 27341 39491 27399 39497
rect 27341 39488 27353 39491
rect 27120 39460 27353 39488
rect 27120 39448 27126 39460
rect 27341 39457 27353 39460
rect 27387 39457 27399 39491
rect 27341 39451 27399 39457
rect 28626 39448 28632 39500
rect 28684 39488 28690 39500
rect 28684 39460 28856 39488
rect 28684 39448 28690 39460
rect 17920 39392 18736 39420
rect 20073 39423 20131 39429
rect 17920 39380 17926 39392
rect 20073 39389 20085 39423
rect 20119 39420 20131 39423
rect 22833 39423 22891 39429
rect 22833 39420 22845 39423
rect 20119 39392 22845 39420
rect 20119 39389 20131 39392
rect 20073 39383 20131 39389
rect 22833 39389 22845 39392
rect 22879 39389 22891 39423
rect 22833 39383 22891 39389
rect 24949 39423 25007 39429
rect 24949 39389 24961 39423
rect 24995 39420 25007 39423
rect 25406 39420 25412 39432
rect 24995 39392 25412 39420
rect 24995 39389 25007 39392
rect 24949 39383 25007 39389
rect 25406 39380 25412 39392
rect 25464 39380 25470 39432
rect 25777 39423 25835 39429
rect 25777 39389 25789 39423
rect 25823 39420 25835 39423
rect 26237 39423 26295 39429
rect 26237 39420 26249 39423
rect 25823 39392 26249 39420
rect 25823 39389 25835 39392
rect 25777 39383 25835 39389
rect 26237 39389 26249 39392
rect 26283 39389 26295 39423
rect 28828 39420 28856 39460
rect 28948 39448 28954 39500
rect 29006 39488 29012 39500
rect 29748 39488 29776 39519
rect 32766 39516 32772 39568
rect 32824 39556 32830 39568
rect 34072 39556 34100 39584
rect 34330 39556 34336 39568
rect 32824 39528 34100 39556
rect 34164 39528 34336 39556
rect 32824 39516 32830 39528
rect 29006 39460 29776 39488
rect 30285 39491 30343 39497
rect 29006 39448 29012 39460
rect 30285 39457 30297 39491
rect 30331 39457 30343 39491
rect 30285 39451 30343 39457
rect 31297 39491 31355 39497
rect 31297 39457 31309 39491
rect 31343 39488 31355 39491
rect 32306 39488 32312 39500
rect 31343 39460 32312 39488
rect 31343 39457 31355 39460
rect 31297 39451 31355 39457
rect 29822 39420 29828 39432
rect 28828 39392 29828 39420
rect 26237 39383 26295 39389
rect 29822 39380 29828 39392
rect 29880 39380 29886 39432
rect 1302 39312 1308 39364
rect 1360 39352 1366 39364
rect 2501 39355 2559 39361
rect 2501 39352 2513 39355
rect 1360 39324 2513 39352
rect 1360 39312 1366 39324
rect 2501 39321 2513 39324
rect 2547 39321 2559 39355
rect 2501 39315 2559 39321
rect 10965 39355 11023 39361
rect 10965 39321 10977 39355
rect 11011 39321 11023 39355
rect 13265 39355 13323 39361
rect 12190 39324 12756 39352
rect 10965 39315 11023 39321
rect 10980 39284 11008 39315
rect 12618 39284 12624 39296
rect 10980 39256 12624 39284
rect 12618 39244 12624 39256
rect 12676 39244 12682 39296
rect 12728 39284 12756 39324
rect 13265 39321 13277 39355
rect 13311 39352 13323 39355
rect 15838 39352 15844 39364
rect 13311 39324 15844 39352
rect 13311 39321 13323 39324
rect 13265 39315 13323 39321
rect 15838 39312 15844 39324
rect 15896 39312 15902 39364
rect 15933 39355 15991 39361
rect 15933 39321 15945 39355
rect 15979 39352 15991 39355
rect 16206 39352 16212 39364
rect 15979 39324 16212 39352
rect 15979 39321 15991 39324
rect 15933 39315 15991 39321
rect 16206 39312 16212 39324
rect 16264 39312 16270 39364
rect 18509 39355 18567 39361
rect 16316 39324 16422 39352
rect 16316 39284 16344 39324
rect 18509 39321 18521 39355
rect 18555 39352 18567 39355
rect 18690 39352 18696 39364
rect 18555 39324 18696 39352
rect 18555 39321 18567 39324
rect 18509 39315 18567 39321
rect 18690 39312 18696 39324
rect 18748 39312 18754 39364
rect 21269 39355 21327 39361
rect 21269 39352 21281 39355
rect 19720 39324 21281 39352
rect 16574 39284 16580 39296
rect 12728 39256 16580 39284
rect 16574 39244 16580 39256
rect 16632 39284 16638 39296
rect 16850 39284 16856 39296
rect 16632 39256 16856 39284
rect 16632 39244 16638 39256
rect 16850 39244 16856 39256
rect 16908 39244 16914 39296
rect 18598 39244 18604 39296
rect 18656 39244 18662 39296
rect 19720 39293 19748 39324
rect 21269 39321 21281 39324
rect 21315 39321 21327 39355
rect 21269 39315 21327 39321
rect 21361 39355 21419 39361
rect 21361 39321 21373 39355
rect 21407 39352 21419 39355
rect 22738 39352 22744 39364
rect 21407 39324 22744 39352
rect 21407 39321 21419 39324
rect 21361 39315 21419 39321
rect 22738 39312 22744 39324
rect 22796 39312 22802 39364
rect 23290 39312 23296 39364
rect 23348 39352 23354 39364
rect 23477 39355 23535 39361
rect 23477 39352 23489 39355
rect 23348 39324 23489 39352
rect 23348 39312 23354 39324
rect 23477 39321 23489 39324
rect 23523 39321 23535 39355
rect 23477 39315 23535 39321
rect 26970 39312 26976 39364
rect 27028 39352 27034 39364
rect 27614 39352 27620 39364
rect 27028 39324 27620 39352
rect 27028 39312 27034 39324
rect 27614 39312 27620 39324
rect 27672 39312 27678 39364
rect 28626 39312 28632 39364
rect 28684 39312 28690 39364
rect 28902 39312 28908 39364
rect 28960 39352 28966 39364
rect 30101 39355 30159 39361
rect 30101 39352 30113 39355
rect 28960 39324 30113 39352
rect 28960 39312 28966 39324
rect 30101 39321 30113 39324
rect 30147 39321 30159 39355
rect 30300 39352 30328 39451
rect 32306 39448 32312 39460
rect 32364 39448 32370 39500
rect 33686 39448 33692 39500
rect 33744 39488 33750 39500
rect 34054 39488 34060 39500
rect 33744 39460 34060 39488
rect 33744 39448 33750 39460
rect 34054 39448 34060 39460
rect 34112 39448 34118 39500
rect 34164 39497 34192 39528
rect 34330 39516 34336 39528
rect 34388 39516 34394 39568
rect 36280 39556 36308 39596
rect 37366 39584 37372 39636
rect 37424 39624 37430 39636
rect 39298 39624 39304 39636
rect 37424 39596 39304 39624
rect 37424 39584 37430 39596
rect 39298 39584 39304 39596
rect 39356 39584 39362 39636
rect 38841 39559 38899 39565
rect 36280 39528 38700 39556
rect 34149 39491 34207 39497
rect 34149 39457 34161 39491
rect 34195 39457 34207 39491
rect 34882 39488 34888 39500
rect 34149 39451 34207 39457
rect 34256 39460 34888 39488
rect 33134 39380 33140 39432
rect 33192 39420 33198 39432
rect 34256 39420 34284 39460
rect 34882 39448 34888 39460
rect 34940 39448 34946 39500
rect 35342 39448 35348 39500
rect 35400 39488 35406 39500
rect 38565 39491 38623 39497
rect 38565 39488 38577 39491
rect 35400 39460 38577 39488
rect 35400 39448 35406 39460
rect 38565 39457 38577 39460
rect 38611 39457 38623 39491
rect 38672 39488 38700 39528
rect 38841 39525 38853 39559
rect 38887 39556 38899 39559
rect 41322 39556 41328 39568
rect 38887 39528 41328 39556
rect 38887 39525 38899 39528
rect 38841 39519 38899 39525
rect 41322 39516 41328 39528
rect 41380 39516 41386 39568
rect 38930 39488 38936 39500
rect 38672 39460 38936 39488
rect 38565 39451 38623 39457
rect 38930 39448 38936 39460
rect 38988 39448 38994 39500
rect 39206 39448 39212 39500
rect 39264 39488 39270 39500
rect 39393 39491 39451 39497
rect 39393 39488 39405 39491
rect 39264 39460 39405 39488
rect 39264 39448 39270 39460
rect 39393 39457 39405 39460
rect 39439 39457 39451 39491
rect 39393 39451 39451 39457
rect 33192 39392 34284 39420
rect 33192 39380 33198 39392
rect 34514 39380 34520 39432
rect 34572 39420 34578 39432
rect 34977 39423 35035 39429
rect 34977 39420 34989 39423
rect 34572 39392 34989 39420
rect 34572 39380 34578 39392
rect 34977 39389 34989 39392
rect 35023 39389 35035 39423
rect 38381 39423 38439 39429
rect 38381 39420 38393 39423
rect 34977 39383 35035 39389
rect 37476 39392 38393 39420
rect 33410 39352 33416 39364
rect 30300 39324 31984 39352
rect 32798 39324 33416 39352
rect 30101 39315 30159 39321
rect 19705 39287 19763 39293
rect 19705 39253 19717 39287
rect 19751 39253 19763 39287
rect 19705 39247 19763 39253
rect 20162 39244 20168 39296
rect 20220 39244 20226 39296
rect 20898 39244 20904 39296
rect 20956 39244 20962 39296
rect 22462 39244 22468 39296
rect 22520 39284 22526 39296
rect 22557 39287 22615 39293
rect 22557 39284 22569 39287
rect 22520 39256 22569 39284
rect 22520 39244 22526 39256
rect 22557 39253 22569 39256
rect 22603 39284 22615 39287
rect 22646 39284 22652 39296
rect 22603 39256 22652 39284
rect 22603 39253 22615 39256
rect 22557 39247 22615 39253
rect 22646 39244 22652 39256
rect 22704 39284 22710 39296
rect 23385 39287 23443 39293
rect 23385 39284 23397 39287
rect 22704 39256 23397 39284
rect 22704 39244 22710 39256
rect 23385 39253 23397 39256
rect 23431 39253 23443 39287
rect 23385 39247 23443 39253
rect 25041 39287 25099 39293
rect 25041 39253 25053 39287
rect 25087 39284 25099 39287
rect 26050 39284 26056 39296
rect 25087 39256 26056 39284
rect 25087 39253 25099 39256
rect 25041 39247 25099 39253
rect 26050 39244 26056 39256
rect 26108 39244 26114 39296
rect 26326 39244 26332 39296
rect 26384 39244 26390 39296
rect 27246 39244 27252 39296
rect 27304 39284 27310 39296
rect 29914 39284 29920 39296
rect 27304 39256 29920 39284
rect 27304 39244 27310 39256
rect 29914 39244 29920 39256
rect 29972 39244 29978 39296
rect 30193 39287 30251 39293
rect 30193 39253 30205 39287
rect 30239 39284 30251 39287
rect 31754 39284 31760 39296
rect 30239 39256 31760 39284
rect 30239 39253 30251 39256
rect 30193 39247 30251 39253
rect 31754 39244 31760 39256
rect 31812 39244 31818 39296
rect 31956 39284 31984 39324
rect 33410 39312 33416 39324
rect 33468 39312 33474 39364
rect 34057 39355 34115 39361
rect 34057 39321 34069 39355
rect 34103 39352 34115 39355
rect 34146 39352 34152 39364
rect 34103 39324 34152 39352
rect 34103 39321 34115 39324
rect 34057 39315 34115 39321
rect 34146 39312 34152 39324
rect 34204 39312 34210 39364
rect 34992 39352 35020 39383
rect 37476 39364 37504 39392
rect 38381 39389 38393 39392
rect 38427 39420 38439 39423
rect 49234 39420 49240 39432
rect 38427 39392 49240 39420
rect 38427 39389 38439 39392
rect 38381 39383 38439 39389
rect 49234 39380 49240 39392
rect 49292 39380 49298 39432
rect 35158 39352 35164 39364
rect 34992 39324 35164 39352
rect 35158 39312 35164 39324
rect 35216 39312 35222 39364
rect 35250 39312 35256 39364
rect 35308 39312 35314 39364
rect 36262 39312 36268 39364
rect 36320 39312 36326 39364
rect 37001 39355 37059 39361
rect 37001 39321 37013 39355
rect 37047 39321 37059 39355
rect 37001 39315 37059 39321
rect 32306 39284 32312 39296
rect 31956 39256 32312 39284
rect 32306 39244 32312 39256
rect 32364 39244 32370 39296
rect 33594 39244 33600 39296
rect 33652 39244 33658 39296
rect 33962 39244 33968 39296
rect 34020 39244 34026 39296
rect 36078 39244 36084 39296
rect 36136 39284 36142 39296
rect 36906 39284 36912 39296
rect 36136 39256 36912 39284
rect 36136 39244 36142 39256
rect 36906 39244 36912 39256
rect 36964 39284 36970 39296
rect 37016 39284 37044 39315
rect 37458 39312 37464 39364
rect 37516 39312 37522 39364
rect 39114 39352 39120 39364
rect 38028 39324 39120 39352
rect 38028 39293 38056 39324
rect 39114 39312 39120 39324
rect 39172 39312 39178 39364
rect 39298 39312 39304 39364
rect 39356 39312 39362 39364
rect 49142 39312 49148 39364
rect 49200 39312 49206 39364
rect 36964 39256 37044 39284
rect 38013 39287 38071 39293
rect 36964 39244 36970 39256
rect 38013 39253 38025 39287
rect 38059 39253 38071 39287
rect 38013 39247 38071 39253
rect 38470 39244 38476 39296
rect 38528 39244 38534 39296
rect 39206 39244 39212 39296
rect 39264 39244 39270 39296
rect 49234 39244 49240 39296
rect 49292 39244 49298 39296
rect 1104 39194 49864 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 27950 39194
rect 28002 39142 28014 39194
rect 28066 39142 28078 39194
rect 28130 39142 28142 39194
rect 28194 39142 28206 39194
rect 28258 39142 37950 39194
rect 38002 39142 38014 39194
rect 38066 39142 38078 39194
rect 38130 39142 38142 39194
rect 38194 39142 38206 39194
rect 38258 39142 47950 39194
rect 48002 39142 48014 39194
rect 48066 39142 48078 39194
rect 48130 39142 48142 39194
rect 48194 39142 48206 39194
rect 48258 39142 49864 39194
rect 1104 39120 49864 39142
rect 15010 39040 15016 39092
rect 15068 39080 15074 39092
rect 15473 39083 15531 39089
rect 15473 39080 15485 39083
rect 15068 39052 15485 39080
rect 15068 39040 15074 39052
rect 15473 39049 15485 39052
rect 15519 39049 15531 39083
rect 15473 39043 15531 39049
rect 15654 39040 15660 39092
rect 15712 39080 15718 39092
rect 15841 39083 15899 39089
rect 15841 39080 15853 39083
rect 15712 39052 15853 39080
rect 15712 39040 15718 39052
rect 15841 39049 15853 39052
rect 15887 39049 15899 39083
rect 15841 39043 15899 39049
rect 16942 39040 16948 39092
rect 17000 39040 17006 39092
rect 17310 39040 17316 39092
rect 17368 39040 17374 39092
rect 17770 39040 17776 39092
rect 17828 39080 17834 39092
rect 17957 39083 18015 39089
rect 17957 39080 17969 39083
rect 17828 39052 17969 39080
rect 17828 39040 17834 39052
rect 17957 39049 17969 39052
rect 18003 39049 18015 39083
rect 17957 39043 18015 39049
rect 18414 39040 18420 39092
rect 18472 39040 18478 39092
rect 19720 39052 21312 39080
rect 14642 38972 14648 39024
rect 14700 39012 14706 39024
rect 17126 39012 17132 39024
rect 14700 38984 17132 39012
rect 14700 38972 14706 38984
rect 17126 38972 17132 38984
rect 17184 38972 17190 39024
rect 17405 39015 17463 39021
rect 17405 38981 17417 39015
rect 17451 39012 17463 39015
rect 19334 39012 19340 39024
rect 17451 38984 19340 39012
rect 17451 38981 17463 38984
rect 17405 38975 17463 38981
rect 19334 38972 19340 38984
rect 19392 38972 19398 39024
rect 15013 38947 15071 38953
rect 15013 38913 15025 38947
rect 15059 38944 15071 38947
rect 17678 38944 17684 38956
rect 15059 38916 17684 38944
rect 15059 38913 15071 38916
rect 15013 38907 15071 38913
rect 17678 38904 17684 38916
rect 17736 38904 17742 38956
rect 18322 38904 18328 38956
rect 18380 38904 18386 38956
rect 19518 38944 19524 38956
rect 18432 38916 19524 38944
rect 15933 38879 15991 38885
rect 15933 38845 15945 38879
rect 15979 38876 15991 38879
rect 16022 38876 16028 38888
rect 15979 38848 16028 38876
rect 15979 38845 15991 38848
rect 15933 38839 15991 38845
rect 16022 38836 16028 38848
rect 16080 38836 16086 38888
rect 16114 38836 16120 38888
rect 16172 38836 16178 38888
rect 17589 38879 17647 38885
rect 17589 38845 17601 38879
rect 17635 38876 17647 38879
rect 18432 38876 18460 38916
rect 19518 38904 19524 38916
rect 19576 38904 19582 38956
rect 19610 38904 19616 38956
rect 19668 38944 19674 38956
rect 19720 38953 19748 39052
rect 20990 38972 20996 39024
rect 21048 38972 21054 39024
rect 19705 38947 19763 38953
rect 19705 38944 19717 38947
rect 19668 38916 19717 38944
rect 19668 38904 19674 38916
rect 19705 38913 19717 38916
rect 19751 38913 19763 38947
rect 21284 38944 21312 39052
rect 21450 39040 21456 39092
rect 21508 39040 21514 39092
rect 21542 39040 21548 39092
rect 21600 39080 21606 39092
rect 23750 39080 23756 39092
rect 21600 39052 23756 39080
rect 21600 39040 21606 39052
rect 23750 39040 23756 39052
rect 23808 39040 23814 39092
rect 24026 39040 24032 39092
rect 24084 39080 24090 39092
rect 24213 39083 24271 39089
rect 24213 39080 24225 39083
rect 24084 39052 24225 39080
rect 24084 39040 24090 39052
rect 24213 39049 24225 39052
rect 24259 39049 24271 39083
rect 24213 39043 24271 39049
rect 24670 39040 24676 39092
rect 24728 39040 24734 39092
rect 26326 39040 26332 39092
rect 26384 39080 26390 39092
rect 27525 39083 27583 39089
rect 27525 39080 27537 39083
rect 26384 39052 27537 39080
rect 26384 39040 26390 39052
rect 27525 39049 27537 39052
rect 27571 39049 27583 39083
rect 27525 39043 27583 39049
rect 27614 39040 27620 39092
rect 27672 39080 27678 39092
rect 27672 39052 30144 39080
rect 27672 39040 27678 39052
rect 21358 38972 21364 39024
rect 21416 39012 21422 39024
rect 22738 39012 22744 39024
rect 21416 38984 22744 39012
rect 21416 38972 21422 38984
rect 22738 38972 22744 38984
rect 22796 38972 22802 39024
rect 25774 39012 25780 39024
rect 23952 38984 25780 39012
rect 21450 38944 21456 38956
rect 21284 38916 21456 38944
rect 19705 38907 19763 38913
rect 21450 38904 21456 38916
rect 21508 38944 21514 38956
rect 22005 38947 22063 38953
rect 22005 38944 22017 38947
rect 21508 38916 22017 38944
rect 21508 38904 21514 38916
rect 22005 38913 22017 38916
rect 22051 38913 22063 38947
rect 22005 38907 22063 38913
rect 17635 38848 18460 38876
rect 18509 38879 18567 38885
rect 17635 38845 17647 38848
rect 17589 38839 17647 38845
rect 18509 38845 18521 38879
rect 18555 38845 18567 38879
rect 18509 38839 18567 38845
rect 19981 38879 20039 38885
rect 19981 38845 19993 38879
rect 20027 38876 20039 38879
rect 21542 38876 21548 38888
rect 20027 38848 21548 38876
rect 20027 38845 20039 38848
rect 19981 38839 20039 38845
rect 16206 38768 16212 38820
rect 16264 38808 16270 38820
rect 18524 38808 18552 38839
rect 21542 38836 21548 38848
rect 21600 38836 21606 38888
rect 22281 38879 22339 38885
rect 22281 38876 22293 38879
rect 22066 38848 22293 38876
rect 16264 38780 18552 38808
rect 16264 38768 16270 38780
rect 21818 38768 21824 38820
rect 21876 38808 21882 38820
rect 22066 38808 22094 38848
rect 22281 38845 22293 38848
rect 22327 38876 22339 38879
rect 23952 38876 23980 38984
rect 25774 38972 25780 38984
rect 25832 38972 25838 39024
rect 27798 39012 27804 39024
rect 25884 38984 27804 39012
rect 24578 38904 24584 38956
rect 24636 38904 24642 38956
rect 25884 38944 25912 38984
rect 27798 38972 27804 38984
rect 27856 38972 27862 39024
rect 30116 39012 30144 39052
rect 30190 39040 30196 39092
rect 30248 39040 30254 39092
rect 31021 39083 31079 39089
rect 31021 39049 31033 39083
rect 31067 39080 31079 39083
rect 31294 39080 31300 39092
rect 31067 39052 31300 39080
rect 31067 39049 31079 39052
rect 31021 39043 31079 39049
rect 31294 39040 31300 39052
rect 31352 39040 31358 39092
rect 31754 39040 31760 39092
rect 31812 39080 31818 39092
rect 31812 39052 31984 39080
rect 31812 39040 31818 39052
rect 30926 39012 30932 39024
rect 30116 38984 30932 39012
rect 30926 38972 30932 38984
rect 30984 38972 30990 39024
rect 31570 38972 31576 39024
rect 31628 39012 31634 39024
rect 31846 39012 31852 39024
rect 31628 38984 31852 39012
rect 31628 38972 31634 38984
rect 31846 38972 31852 38984
rect 31904 38972 31910 39024
rect 31956 39012 31984 39052
rect 33594 39040 33600 39092
rect 33652 39080 33658 39092
rect 34425 39083 34483 39089
rect 34425 39080 34437 39083
rect 33652 39052 34437 39080
rect 33652 39040 33658 39052
rect 34425 39049 34437 39052
rect 34471 39049 34483 39083
rect 34425 39043 34483 39049
rect 35250 39040 35256 39092
rect 35308 39080 35314 39092
rect 36909 39083 36967 39089
rect 36909 39080 36921 39083
rect 35308 39052 36921 39080
rect 35308 39040 35314 39052
rect 36909 39049 36921 39052
rect 36955 39080 36967 39083
rect 37826 39080 37832 39092
rect 36955 39052 37832 39080
rect 36955 39049 36967 39052
rect 36909 39043 36967 39049
rect 37826 39040 37832 39052
rect 37884 39040 37890 39092
rect 38654 39040 38660 39092
rect 38712 39080 38718 39092
rect 39117 39083 39175 39089
rect 39117 39080 39129 39083
rect 38712 39052 39129 39080
rect 38712 39040 38718 39052
rect 39117 39049 39129 39052
rect 39163 39049 39175 39083
rect 39117 39043 39175 39049
rect 34606 39012 34612 39024
rect 31956 38984 34612 39012
rect 34606 38972 34612 38984
rect 34664 38972 34670 39024
rect 36170 38972 36176 39024
rect 36228 38972 36234 39024
rect 37642 38972 37648 39024
rect 37700 39012 37706 39024
rect 37700 38984 41414 39012
rect 37700 38972 37706 38984
rect 24675 38916 25912 38944
rect 24675 38876 24703 38916
rect 27246 38904 27252 38956
rect 27304 38944 27310 38956
rect 27304 38916 27752 38944
rect 27304 38904 27310 38916
rect 22327 38848 23980 38876
rect 24044 38848 24703 38876
rect 22327 38845 22339 38848
rect 22281 38839 22339 38845
rect 21876 38780 22094 38808
rect 21876 38768 21882 38780
rect 14829 38743 14887 38749
rect 14829 38709 14841 38743
rect 14875 38740 14887 38743
rect 15102 38740 15108 38752
rect 14875 38712 15108 38740
rect 14875 38709 14887 38712
rect 14829 38703 14887 38709
rect 15102 38700 15108 38712
rect 15160 38700 15166 38752
rect 15838 38700 15844 38752
rect 15896 38740 15902 38752
rect 21082 38740 21088 38752
rect 15896 38712 21088 38740
rect 15896 38700 15902 38712
rect 21082 38700 21088 38712
rect 21140 38740 21146 38752
rect 24044 38740 24072 38848
rect 24762 38836 24768 38888
rect 24820 38836 24826 38888
rect 27338 38836 27344 38888
rect 27396 38876 27402 38888
rect 27724 38885 27752 38916
rect 29822 38904 29828 38956
rect 29880 38944 29886 38956
rect 30650 38944 30656 38956
rect 29880 38916 30656 38944
rect 29880 38904 29886 38916
rect 30650 38904 30656 38916
rect 30708 38904 30714 38956
rect 31389 38947 31447 38953
rect 31389 38913 31401 38947
rect 31435 38944 31447 38947
rect 32214 38944 32220 38956
rect 31435 38916 32220 38944
rect 31435 38913 31447 38916
rect 31389 38907 31447 38913
rect 32214 38904 32220 38916
rect 32272 38904 32278 38956
rect 33137 38947 33195 38953
rect 33137 38913 33149 38947
rect 33183 38944 33195 38947
rect 33594 38944 33600 38956
rect 33183 38916 33600 38944
rect 33183 38913 33195 38916
rect 33137 38907 33195 38913
rect 33594 38904 33600 38916
rect 33652 38904 33658 38956
rect 33962 38904 33968 38956
rect 34020 38944 34026 38956
rect 34333 38947 34391 38953
rect 34333 38944 34345 38947
rect 34020 38916 34345 38944
rect 34020 38904 34026 38916
rect 34333 38913 34345 38916
rect 34379 38913 34391 38947
rect 34333 38907 34391 38913
rect 35158 38904 35164 38956
rect 35216 38904 35222 38956
rect 38102 38904 38108 38956
rect 38160 38944 38166 38956
rect 39025 38947 39083 38953
rect 39025 38944 39037 38947
rect 38160 38916 39037 38944
rect 38160 38904 38166 38916
rect 39025 38913 39037 38916
rect 39071 38944 39083 38947
rect 39298 38944 39304 38956
rect 39071 38916 39304 38944
rect 39071 38913 39083 38916
rect 39025 38907 39083 38913
rect 39298 38904 39304 38916
rect 39356 38904 39362 38956
rect 41386 38944 41414 38984
rect 49234 38944 49240 38956
rect 41386 38916 49240 38944
rect 49234 38904 49240 38916
rect 49292 38904 49298 38956
rect 27617 38879 27675 38885
rect 27617 38876 27629 38879
rect 27396 38848 27629 38876
rect 27396 38836 27402 38848
rect 27617 38845 27629 38848
rect 27663 38845 27675 38879
rect 27617 38839 27675 38845
rect 27709 38879 27767 38885
rect 27709 38845 27721 38879
rect 27755 38845 27767 38879
rect 27709 38839 27767 38845
rect 28442 38836 28448 38888
rect 28500 38836 28506 38888
rect 28721 38879 28779 38885
rect 28721 38845 28733 38879
rect 28767 38876 28779 38879
rect 29178 38876 29184 38888
rect 28767 38848 29184 38876
rect 28767 38845 28779 38848
rect 28721 38839 28779 38845
rect 29178 38836 29184 38848
rect 29236 38836 29242 38888
rect 29270 38836 29276 38888
rect 29328 38876 29334 38888
rect 31481 38879 31539 38885
rect 31481 38876 31493 38879
rect 29328 38848 31493 38876
rect 29328 38836 29334 38848
rect 31481 38845 31493 38848
rect 31527 38845 31539 38879
rect 31481 38839 31539 38845
rect 31665 38879 31723 38885
rect 31665 38845 31677 38879
rect 31711 38876 31723 38879
rect 32674 38876 32680 38888
rect 31711 38848 32680 38876
rect 31711 38845 31723 38848
rect 31665 38839 31723 38845
rect 32674 38836 32680 38848
rect 32732 38836 32738 38888
rect 33229 38879 33287 38885
rect 33229 38845 33241 38879
rect 33275 38845 33287 38879
rect 33229 38839 33287 38845
rect 33413 38879 33471 38885
rect 33413 38845 33425 38879
rect 33459 38876 33471 38879
rect 33686 38876 33692 38888
rect 33459 38848 33692 38876
rect 33459 38845 33471 38848
rect 33413 38839 33471 38845
rect 24486 38768 24492 38820
rect 24544 38808 24550 38820
rect 25593 38811 25651 38817
rect 25593 38808 25605 38811
rect 24544 38780 25605 38808
rect 24544 38768 24550 38780
rect 25593 38777 25605 38780
rect 25639 38777 25651 38811
rect 33134 38808 33140 38820
rect 25593 38771 25651 38777
rect 29748 38780 33140 38808
rect 21140 38712 24072 38740
rect 21140 38700 21146 38712
rect 24578 38700 24584 38752
rect 24636 38740 24642 38752
rect 24762 38740 24768 38752
rect 24636 38712 24768 38740
rect 24636 38700 24642 38712
rect 24762 38700 24768 38712
rect 24820 38700 24826 38752
rect 26234 38700 26240 38752
rect 26292 38740 26298 38752
rect 27157 38743 27215 38749
rect 27157 38740 27169 38743
rect 26292 38712 27169 38740
rect 26292 38700 26298 38712
rect 27157 38709 27169 38712
rect 27203 38709 27215 38743
rect 27157 38703 27215 38709
rect 27338 38700 27344 38752
rect 27396 38740 27402 38752
rect 29748 38740 29776 38780
rect 33134 38768 33140 38780
rect 33192 38768 33198 38820
rect 33244 38808 33272 38839
rect 33686 38836 33692 38848
rect 33744 38836 33750 38888
rect 33870 38836 33876 38888
rect 33928 38876 33934 38888
rect 34517 38879 34575 38885
rect 34517 38876 34529 38879
rect 33928 38848 34529 38876
rect 33928 38836 33934 38848
rect 34517 38845 34529 38848
rect 34563 38845 34575 38879
rect 34517 38839 34575 38845
rect 35434 38836 35440 38888
rect 35492 38836 35498 38888
rect 36906 38836 36912 38888
rect 36964 38876 36970 38888
rect 39209 38879 39267 38885
rect 39209 38876 39221 38879
rect 36964 38848 39221 38876
rect 36964 38836 36970 38848
rect 39209 38845 39221 38848
rect 39255 38845 39267 38879
rect 39209 38839 39267 38845
rect 35066 38808 35072 38820
rect 33244 38780 35072 38808
rect 35066 38768 35072 38780
rect 35124 38768 35130 38820
rect 38838 38808 38844 38820
rect 36832 38780 38844 38808
rect 27396 38712 29776 38740
rect 27396 38700 27402 38712
rect 29914 38700 29920 38752
rect 29972 38740 29978 38752
rect 32769 38743 32827 38749
rect 32769 38740 32781 38743
rect 29972 38712 32781 38740
rect 29972 38700 29978 38712
rect 32769 38709 32781 38712
rect 32815 38709 32827 38743
rect 32769 38703 32827 38709
rect 33965 38743 34023 38749
rect 33965 38709 33977 38743
rect 34011 38740 34023 38743
rect 36832 38740 36860 38780
rect 38838 38768 38844 38780
rect 38896 38768 38902 38820
rect 34011 38712 36860 38740
rect 34011 38709 34023 38712
rect 33965 38703 34023 38709
rect 38654 38700 38660 38752
rect 38712 38700 38718 38752
rect 1104 38650 49864 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 32950 38650
rect 33002 38598 33014 38650
rect 33066 38598 33078 38650
rect 33130 38598 33142 38650
rect 33194 38598 33206 38650
rect 33258 38598 42950 38650
rect 43002 38598 43014 38650
rect 43066 38598 43078 38650
rect 43130 38598 43142 38650
rect 43194 38598 43206 38650
rect 43258 38598 49864 38650
rect 1104 38576 49864 38598
rect 8386 38496 8392 38548
rect 8444 38496 8450 38548
rect 12434 38496 12440 38548
rect 12492 38496 12498 38548
rect 12710 38496 12716 38548
rect 12768 38536 12774 38548
rect 14366 38536 14372 38548
rect 12768 38508 14372 38536
rect 12768 38496 12774 38508
rect 14366 38496 14372 38508
rect 14424 38496 14430 38548
rect 16853 38539 16911 38545
rect 16853 38536 16865 38539
rect 14476 38508 16865 38536
rect 1762 38428 1768 38480
rect 1820 38468 1826 38480
rect 14476 38468 14504 38508
rect 16853 38505 16865 38508
rect 16899 38505 16911 38539
rect 16853 38499 16911 38505
rect 17862 38496 17868 38548
rect 17920 38536 17926 38548
rect 18966 38536 18972 38548
rect 17920 38508 18972 38536
rect 17920 38496 17926 38508
rect 18966 38496 18972 38508
rect 19024 38496 19030 38548
rect 19521 38539 19579 38545
rect 19521 38505 19533 38539
rect 19567 38536 19579 38539
rect 20162 38536 20168 38548
rect 19567 38508 20168 38536
rect 19567 38505 19579 38508
rect 19521 38499 19579 38505
rect 20162 38496 20168 38508
rect 20220 38496 20226 38548
rect 21266 38496 21272 38548
rect 21324 38536 21330 38548
rect 22097 38539 22155 38545
rect 22097 38536 22109 38539
rect 21324 38508 22109 38536
rect 21324 38496 21330 38508
rect 22097 38505 22109 38508
rect 22143 38505 22155 38539
rect 22097 38499 22155 38505
rect 24946 38496 24952 38548
rect 25004 38536 25010 38548
rect 25133 38539 25191 38545
rect 25133 38536 25145 38539
rect 25004 38508 25145 38536
rect 25004 38496 25010 38508
rect 25133 38505 25145 38508
rect 25179 38505 25191 38539
rect 25133 38499 25191 38505
rect 25682 38496 25688 38548
rect 25740 38536 25746 38548
rect 26329 38539 26387 38545
rect 26329 38536 26341 38539
rect 25740 38508 26341 38536
rect 25740 38496 25746 38508
rect 26329 38505 26341 38508
rect 26375 38536 26387 38539
rect 26375 38508 27752 38536
rect 26375 38505 26387 38508
rect 26329 38499 26387 38505
rect 1820 38440 9674 38468
rect 1820 38428 1826 38440
rect 1302 38360 1308 38412
rect 1360 38400 1366 38412
rect 2041 38403 2099 38409
rect 2041 38400 2053 38403
rect 1360 38372 2053 38400
rect 1360 38360 1366 38372
rect 2041 38369 2053 38372
rect 2087 38369 2099 38403
rect 9646 38400 9674 38440
rect 12820 38440 14504 38468
rect 12820 38400 12848 38440
rect 16206 38428 16212 38480
rect 16264 38428 16270 38480
rect 17034 38428 17040 38480
rect 17092 38468 17098 38480
rect 20070 38468 20076 38480
rect 17092 38440 20076 38468
rect 17092 38428 17098 38440
rect 20070 38428 20076 38440
rect 20128 38428 20134 38480
rect 21818 38468 21824 38480
rect 20180 38440 21824 38468
rect 9646 38372 12848 38400
rect 12989 38403 13047 38409
rect 2041 38363 2099 38369
rect 12989 38369 13001 38403
rect 13035 38369 13047 38403
rect 12989 38363 13047 38369
rect 1765 38335 1823 38341
rect 1765 38301 1777 38335
rect 1811 38332 1823 38335
rect 12710 38332 12716 38344
rect 1811 38304 12716 38332
rect 1811 38301 1823 38304
rect 1765 38295 1823 38301
rect 12710 38292 12716 38304
rect 12768 38292 12774 38344
rect 12802 38292 12808 38344
rect 12860 38332 12866 38344
rect 12897 38335 12955 38341
rect 12897 38332 12909 38335
rect 12860 38304 12909 38332
rect 12860 38292 12866 38304
rect 12897 38301 12909 38304
rect 12943 38301 12955 38335
rect 13004 38332 13032 38363
rect 14458 38360 14464 38412
rect 14516 38360 14522 38412
rect 18874 38400 18880 38412
rect 16776 38372 18880 38400
rect 16776 38341 16804 38372
rect 18874 38360 18880 38372
rect 18932 38360 18938 38412
rect 20180 38409 20208 38440
rect 21818 38428 21824 38440
rect 21876 38428 21882 38480
rect 23293 38471 23351 38477
rect 23293 38437 23305 38471
rect 23339 38437 23351 38471
rect 23293 38431 23351 38437
rect 20165 38403 20223 38409
rect 20165 38369 20177 38403
rect 20211 38369 20223 38403
rect 20165 38363 20223 38369
rect 22738 38360 22744 38412
rect 22796 38360 22802 38412
rect 16761 38335 16819 38341
rect 13004 38304 13216 38332
rect 12897 38295 12955 38301
rect 8297 38267 8355 38273
rect 8297 38233 8309 38267
rect 8343 38264 8355 38267
rect 13188 38264 13216 38304
rect 16761 38301 16773 38335
rect 16807 38301 16819 38335
rect 16761 38295 16819 38301
rect 16850 38292 16856 38344
rect 16908 38332 16914 38344
rect 18693 38335 18751 38341
rect 18693 38332 18705 38335
rect 16908 38304 18705 38332
rect 16908 38292 16914 38304
rect 18693 38301 18705 38304
rect 18739 38301 18751 38335
rect 18693 38295 18751 38301
rect 19426 38292 19432 38344
rect 19484 38332 19490 38344
rect 19889 38335 19947 38341
rect 19889 38332 19901 38335
rect 19484 38304 19901 38332
rect 19484 38292 19490 38304
rect 19889 38301 19901 38304
rect 19935 38301 19947 38335
rect 19889 38295 19947 38301
rect 19978 38292 19984 38344
rect 20036 38292 20042 38344
rect 21726 38292 21732 38344
rect 21784 38332 21790 38344
rect 23308 38332 23336 38431
rect 25590 38428 25596 38480
rect 25648 38468 25654 38480
rect 27724 38468 27752 38508
rect 28534 38496 28540 38548
rect 28592 38536 28598 38548
rect 28592 38508 31754 38536
rect 28592 38496 28598 38508
rect 29638 38468 29644 38480
rect 25648 38440 27660 38468
rect 27724 38440 29644 38468
rect 25648 38428 25654 38440
rect 23937 38403 23995 38409
rect 23937 38369 23949 38403
rect 23983 38400 23995 38403
rect 24670 38400 24676 38412
rect 23983 38372 24676 38400
rect 23983 38369 23995 38372
rect 23937 38363 23995 38369
rect 24670 38360 24676 38372
rect 24728 38360 24734 38412
rect 25774 38360 25780 38412
rect 25832 38360 25838 38412
rect 26878 38360 26884 38412
rect 26936 38400 26942 38412
rect 26936 38372 27384 38400
rect 26936 38360 26942 38372
rect 21784 38304 23336 38332
rect 23753 38335 23811 38341
rect 21784 38292 21790 38304
rect 23753 38301 23765 38335
rect 23799 38332 23811 38335
rect 27154 38332 27160 38344
rect 23799 38304 27160 38332
rect 23799 38301 23811 38304
rect 23753 38295 23811 38301
rect 27154 38292 27160 38304
rect 27212 38292 27218 38344
rect 27356 38332 27384 38372
rect 27430 38360 27436 38412
rect 27488 38400 27494 38412
rect 27632 38409 27660 38440
rect 29638 38428 29644 38440
rect 29696 38428 29702 38480
rect 31726 38468 31754 38508
rect 32122 38496 32128 38548
rect 32180 38536 32186 38548
rect 37461 38539 37519 38545
rect 32180 38508 37412 38536
rect 32180 38496 32186 38508
rect 36265 38471 36323 38477
rect 36265 38468 36277 38471
rect 31726 38440 36277 38468
rect 36265 38437 36277 38440
rect 36311 38437 36323 38471
rect 37384 38468 37412 38508
rect 37461 38505 37473 38539
rect 37507 38536 37519 38539
rect 39206 38536 39212 38548
rect 37507 38508 39212 38536
rect 37507 38505 37519 38508
rect 37461 38499 37519 38505
rect 39206 38496 39212 38508
rect 39264 38496 39270 38548
rect 38289 38471 38347 38477
rect 37384 38440 38148 38468
rect 36265 38431 36323 38437
rect 27525 38403 27583 38409
rect 27525 38400 27537 38403
rect 27488 38372 27537 38400
rect 27488 38360 27494 38372
rect 27525 38369 27537 38372
rect 27571 38369 27583 38403
rect 27525 38363 27583 38369
rect 27617 38403 27675 38409
rect 27617 38369 27629 38403
rect 27663 38369 27675 38403
rect 27617 38363 27675 38369
rect 31938 38360 31944 38412
rect 31996 38400 32002 38412
rect 33505 38403 33563 38409
rect 33505 38400 33517 38403
rect 31996 38372 33517 38400
rect 31996 38360 32002 38372
rect 33505 38369 33517 38372
rect 33551 38369 33563 38403
rect 33505 38363 33563 38369
rect 33689 38403 33747 38409
rect 33689 38369 33701 38403
rect 33735 38400 33747 38403
rect 35434 38400 35440 38412
rect 33735 38372 35440 38400
rect 33735 38369 33747 38372
rect 33689 38363 33747 38369
rect 35434 38360 35440 38372
rect 35492 38360 35498 38412
rect 36814 38360 36820 38412
rect 36872 38360 36878 38412
rect 37734 38360 37740 38412
rect 37792 38400 37798 38412
rect 38013 38403 38071 38409
rect 38013 38400 38025 38403
rect 37792 38372 38025 38400
rect 37792 38360 37798 38372
rect 38013 38369 38025 38372
rect 38059 38369 38071 38403
rect 38120 38400 38148 38440
rect 38289 38437 38301 38471
rect 38335 38468 38347 38471
rect 39666 38468 39672 38480
rect 38335 38440 39672 38468
rect 38335 38437 38347 38440
rect 38289 38431 38347 38437
rect 39666 38428 39672 38440
rect 39724 38428 39730 38480
rect 38749 38403 38807 38409
rect 38749 38400 38761 38403
rect 38120 38372 38761 38400
rect 38013 38363 38071 38369
rect 38749 38369 38761 38372
rect 38795 38369 38807 38403
rect 38749 38363 38807 38369
rect 38930 38360 38936 38412
rect 38988 38360 38994 38412
rect 27356 38304 28396 38332
rect 14737 38267 14795 38273
rect 14737 38264 14749 38267
rect 8343 38236 13032 38264
rect 13188 38236 14749 38264
rect 8343 38233 8355 38236
rect 8297 38227 8355 38233
rect 12805 38199 12863 38205
rect 12805 38165 12817 38199
rect 12851 38196 12863 38199
rect 12894 38196 12900 38208
rect 12851 38168 12900 38196
rect 12851 38165 12863 38168
rect 12805 38159 12863 38165
rect 12894 38156 12900 38168
rect 12952 38156 12958 38208
rect 13004 38196 13032 38236
rect 14737 38233 14749 38236
rect 14783 38264 14795 38267
rect 14826 38264 14832 38276
rect 14783 38236 14832 38264
rect 14783 38233 14795 38236
rect 14737 38227 14795 38233
rect 14826 38224 14832 38236
rect 14884 38224 14890 38276
rect 16666 38264 16672 38276
rect 15962 38236 16672 38264
rect 16666 38224 16672 38236
rect 16724 38224 16730 38276
rect 17313 38267 17371 38273
rect 17313 38233 17325 38267
rect 17359 38264 17371 38267
rect 17957 38267 18015 38273
rect 17359 38236 17908 38264
rect 17359 38233 17371 38236
rect 17313 38227 17371 38233
rect 15102 38196 15108 38208
rect 13004 38168 15108 38196
rect 15102 38156 15108 38168
rect 15160 38156 15166 38208
rect 17402 38156 17408 38208
rect 17460 38156 17466 38208
rect 17880 38196 17908 38236
rect 17957 38233 17969 38267
rect 18003 38264 18015 38267
rect 18598 38264 18604 38276
rect 18003 38236 18604 38264
rect 18003 38233 18015 38236
rect 17957 38227 18015 38233
rect 18598 38224 18604 38236
rect 18656 38264 18662 38276
rect 20717 38267 20775 38273
rect 20717 38264 20729 38267
rect 18656 38236 20729 38264
rect 18656 38224 18662 38236
rect 20717 38233 20729 38236
rect 20763 38233 20775 38267
rect 20717 38227 20775 38233
rect 21450 38224 21456 38276
rect 21508 38224 21514 38276
rect 22465 38267 22523 38273
rect 22465 38233 22477 38267
rect 22511 38264 22523 38267
rect 22511 38236 23244 38264
rect 22511 38233 22523 38236
rect 22465 38227 22523 38233
rect 20898 38196 20904 38208
rect 17880 38168 20904 38196
rect 20898 38156 20904 38168
rect 20956 38156 20962 38208
rect 22554 38156 22560 38208
rect 22612 38156 22618 38208
rect 23216 38196 23244 38236
rect 23290 38224 23296 38276
rect 23348 38264 23354 38276
rect 23348 38236 25820 38264
rect 23348 38224 23354 38236
rect 23566 38196 23572 38208
rect 23216 38168 23572 38196
rect 23566 38156 23572 38168
rect 23624 38156 23630 38208
rect 23658 38156 23664 38208
rect 23716 38156 23722 38208
rect 25314 38156 25320 38208
rect 25372 38196 25378 38208
rect 25501 38199 25559 38205
rect 25501 38196 25513 38199
rect 25372 38168 25513 38196
rect 25372 38156 25378 38168
rect 25501 38165 25513 38168
rect 25547 38165 25559 38199
rect 25501 38159 25559 38165
rect 25593 38199 25651 38205
rect 25593 38165 25605 38199
rect 25639 38196 25651 38199
rect 25682 38196 25688 38208
rect 25639 38168 25688 38196
rect 25639 38165 25651 38168
rect 25593 38159 25651 38165
rect 25682 38156 25688 38168
rect 25740 38156 25746 38208
rect 25792 38196 25820 38236
rect 26418 38224 26424 38276
rect 26476 38264 26482 38276
rect 26476 38236 27476 38264
rect 26476 38224 26482 38236
rect 27448 38208 27476 38236
rect 27614 38224 27620 38276
rect 27672 38264 27678 38276
rect 28261 38267 28319 38273
rect 28261 38264 28273 38267
rect 27672 38236 28273 38264
rect 27672 38224 27678 38236
rect 28261 38233 28273 38236
rect 28307 38233 28319 38267
rect 28368 38264 28396 38304
rect 28442 38292 28448 38344
rect 28500 38332 28506 38344
rect 29089 38335 29147 38341
rect 29089 38332 29101 38335
rect 28500 38304 29101 38332
rect 28500 38292 28506 38304
rect 29089 38301 29101 38304
rect 29135 38332 29147 38335
rect 29733 38335 29791 38341
rect 29733 38332 29745 38335
rect 29135 38304 29745 38332
rect 29135 38301 29147 38304
rect 29089 38295 29147 38301
rect 29733 38301 29745 38304
rect 29779 38301 29791 38335
rect 29733 38295 29791 38301
rect 32214 38292 32220 38344
rect 32272 38292 32278 38344
rect 36630 38332 36636 38344
rect 32968 38304 36636 38332
rect 30009 38267 30067 38273
rect 30009 38264 30021 38267
rect 28368 38236 30021 38264
rect 28261 38227 28319 38233
rect 30009 38233 30021 38236
rect 30055 38233 30067 38267
rect 31294 38264 31300 38276
rect 31234 38236 31300 38264
rect 30009 38227 30067 38233
rect 27065 38199 27123 38205
rect 27065 38196 27077 38199
rect 25792 38168 27077 38196
rect 27065 38165 27077 38168
rect 27111 38165 27123 38199
rect 27065 38159 27123 38165
rect 27430 38156 27436 38208
rect 27488 38156 27494 38208
rect 30024 38196 30052 38227
rect 31294 38224 31300 38236
rect 31352 38224 31358 38276
rect 31570 38264 31576 38276
rect 31404 38236 31576 38264
rect 31404 38196 31432 38236
rect 31570 38224 31576 38236
rect 31628 38224 31634 38276
rect 30024 38168 31432 38196
rect 31478 38156 31484 38208
rect 31536 38196 31542 38208
rect 32968 38196 32996 38304
rect 36630 38292 36636 38304
rect 36688 38292 36694 38344
rect 37921 38335 37979 38341
rect 37921 38301 37933 38335
rect 37967 38332 37979 38335
rect 38654 38332 38660 38344
rect 37967 38304 38660 38332
rect 37967 38301 37979 38304
rect 37921 38295 37979 38301
rect 38654 38292 38660 38304
rect 38712 38292 38718 38344
rect 33060 38236 34836 38264
rect 33060 38205 33088 38236
rect 31536 38168 32996 38196
rect 33045 38199 33103 38205
rect 31536 38156 31542 38168
rect 33045 38165 33057 38199
rect 33091 38165 33103 38199
rect 33045 38159 33103 38165
rect 33410 38156 33416 38208
rect 33468 38156 33474 38208
rect 33870 38156 33876 38208
rect 33928 38196 33934 38208
rect 34238 38196 34244 38208
rect 33928 38168 34244 38196
rect 33928 38156 33934 38168
rect 34238 38156 34244 38168
rect 34296 38156 34302 38208
rect 34808 38196 34836 38236
rect 34882 38224 34888 38276
rect 34940 38224 34946 38276
rect 35158 38224 35164 38276
rect 35216 38264 35222 38276
rect 35621 38267 35679 38273
rect 35621 38264 35633 38267
rect 35216 38236 35633 38264
rect 35216 38224 35222 38236
rect 35621 38233 35633 38236
rect 35667 38233 35679 38267
rect 35621 38227 35679 38233
rect 36170 38224 36176 38276
rect 36228 38264 36234 38276
rect 37829 38267 37887 38273
rect 37829 38264 37841 38267
rect 36228 38236 37841 38264
rect 36228 38224 36234 38236
rect 37829 38233 37841 38236
rect 37875 38233 37887 38267
rect 38838 38264 38844 38276
rect 37829 38227 37887 38233
rect 38672 38236 38844 38264
rect 36446 38196 36452 38208
rect 34808 38168 36452 38196
rect 36446 38156 36452 38168
rect 36504 38156 36510 38208
rect 36630 38156 36636 38208
rect 36688 38156 36694 38208
rect 36722 38156 36728 38208
rect 36780 38156 36786 38208
rect 38672 38205 38700 38236
rect 38838 38224 38844 38236
rect 38896 38224 38902 38276
rect 49142 38224 49148 38276
rect 49200 38224 49206 38276
rect 38657 38199 38715 38205
rect 38657 38165 38669 38199
rect 38703 38165 38715 38199
rect 38657 38159 38715 38165
rect 49234 38156 49240 38208
rect 49292 38156 49298 38208
rect 1104 38106 49864 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 27950 38106
rect 28002 38054 28014 38106
rect 28066 38054 28078 38106
rect 28130 38054 28142 38106
rect 28194 38054 28206 38106
rect 28258 38054 37950 38106
rect 38002 38054 38014 38106
rect 38066 38054 38078 38106
rect 38130 38054 38142 38106
rect 38194 38054 38206 38106
rect 38258 38054 47950 38106
rect 48002 38054 48014 38106
rect 48066 38054 48078 38106
rect 48130 38054 48142 38106
rect 48194 38054 48206 38106
rect 48258 38054 49864 38106
rect 1104 38032 49864 38054
rect 15194 37992 15200 38004
rect 12406 37964 15200 37992
rect 8481 37927 8539 37933
rect 8481 37893 8493 37927
rect 8527 37924 8539 37927
rect 12406 37924 12434 37964
rect 15194 37952 15200 37964
rect 15252 37952 15258 38004
rect 17957 37995 18015 38001
rect 17957 37961 17969 37995
rect 18003 37992 18015 37995
rect 18506 37992 18512 38004
rect 18003 37964 18512 37992
rect 18003 37961 18015 37964
rect 17957 37955 18015 37961
rect 18506 37952 18512 37964
rect 18564 37952 18570 38004
rect 20714 37952 20720 38004
rect 20772 37952 20778 38004
rect 21085 37995 21143 38001
rect 21085 37961 21097 37995
rect 21131 37992 21143 37995
rect 21634 37992 21640 38004
rect 21131 37964 21640 37992
rect 21131 37961 21143 37964
rect 21085 37955 21143 37961
rect 16666 37924 16672 37936
rect 8527 37896 12434 37924
rect 16054 37896 16672 37924
rect 8527 37893 8539 37896
rect 8481 37887 8539 37893
rect 16666 37884 16672 37896
rect 16724 37884 16730 37936
rect 19337 37927 19395 37933
rect 19337 37924 19349 37927
rect 17512 37896 19349 37924
rect 1762 37816 1768 37868
rect 1820 37816 1826 37868
rect 12894 37816 12900 37868
rect 12952 37856 12958 37868
rect 12989 37859 13047 37865
rect 12989 37856 13001 37859
rect 12952 37828 13001 37856
rect 12952 37816 12958 37828
rect 12989 37825 13001 37828
rect 13035 37825 13047 37859
rect 12989 37819 13047 37825
rect 14458 37816 14464 37868
rect 14516 37856 14522 37868
rect 17512 37865 17540 37896
rect 19337 37893 19349 37896
rect 19383 37893 19395 37927
rect 19337 37887 19395 37893
rect 20257 37927 20315 37933
rect 20257 37893 20269 37927
rect 20303 37924 20315 37927
rect 21100 37924 21128 37955
rect 21634 37952 21640 37964
rect 21692 37952 21698 38004
rect 22554 37952 22560 38004
rect 22612 37992 22618 38004
rect 25685 37995 25743 38001
rect 25685 37992 25697 37995
rect 22612 37964 25697 37992
rect 22612 37952 22618 37964
rect 25685 37961 25697 37964
rect 25731 37961 25743 37995
rect 28442 37992 28448 38004
rect 25685 37955 25743 37961
rect 27172 37964 28448 37992
rect 20303 37896 21128 37924
rect 21177 37927 21235 37933
rect 20303 37893 20315 37896
rect 20257 37887 20315 37893
rect 21177 37893 21189 37927
rect 21223 37924 21235 37927
rect 21542 37924 21548 37936
rect 21223 37896 21548 37924
rect 21223 37893 21235 37896
rect 21177 37887 21235 37893
rect 21542 37884 21548 37896
rect 21600 37884 21606 37936
rect 24949 37927 25007 37933
rect 24949 37893 24961 37927
rect 24995 37924 25007 37927
rect 26234 37924 26240 37936
rect 24995 37896 26240 37924
rect 24995 37893 25007 37896
rect 24949 37887 25007 37893
rect 26234 37884 26240 37896
rect 26292 37884 26298 37936
rect 27172 37868 27200 37964
rect 28442 37952 28448 37964
rect 28500 37952 28506 38004
rect 28810 37952 28816 38004
rect 28868 37992 28874 38004
rect 28905 37995 28963 38001
rect 28905 37992 28917 37995
rect 28868 37964 28917 37992
rect 28868 37952 28874 37964
rect 28905 37961 28917 37964
rect 28951 37961 28963 37995
rect 28905 37955 28963 37961
rect 30926 37952 30932 38004
rect 30984 37992 30990 38004
rect 31481 37995 31539 38001
rect 31481 37992 31493 37995
rect 30984 37964 31493 37992
rect 30984 37952 30990 37964
rect 31481 37961 31493 37964
rect 31527 37961 31539 37995
rect 35158 37992 35164 38004
rect 31481 37955 31539 37961
rect 32416 37964 35164 37992
rect 28166 37884 28172 37936
rect 28224 37884 28230 37936
rect 29914 37924 29920 37936
rect 29748 37896 29920 37924
rect 14553 37859 14611 37865
rect 14553 37856 14565 37859
rect 14516 37828 14565 37856
rect 14516 37816 14522 37828
rect 14553 37825 14565 37828
rect 14599 37825 14611 37859
rect 14553 37819 14611 37825
rect 17497 37859 17555 37865
rect 17497 37825 17509 37859
rect 17543 37825 17555 37859
rect 17497 37819 17555 37825
rect 18325 37859 18383 37865
rect 18325 37825 18337 37859
rect 18371 37856 18383 37859
rect 20990 37856 20996 37868
rect 18371 37828 20996 37856
rect 18371 37825 18383 37828
rect 18325 37819 18383 37825
rect 20990 37816 20996 37828
rect 21048 37816 21054 37868
rect 21450 37816 21456 37868
rect 21508 37856 21514 37868
rect 22002 37856 22008 37868
rect 21508 37828 22008 37856
rect 21508 37816 21514 37828
rect 22002 37816 22008 37828
rect 22060 37816 22066 37868
rect 23382 37816 23388 37868
rect 23440 37816 23446 37868
rect 23750 37816 23756 37868
rect 23808 37856 23814 37868
rect 24762 37856 24768 37868
rect 23808 37828 24768 37856
rect 23808 37816 23814 37828
rect 24762 37816 24768 37828
rect 24820 37816 24826 37868
rect 24854 37816 24860 37868
rect 24912 37816 24918 37868
rect 25866 37816 25872 37868
rect 25924 37856 25930 37868
rect 26053 37859 26111 37865
rect 26053 37856 26065 37859
rect 25924 37828 26065 37856
rect 25924 37816 25930 37828
rect 26053 37825 26065 37828
rect 26099 37825 26111 37859
rect 26053 37819 26111 37825
rect 27154 37816 27160 37868
rect 27212 37816 27218 37868
rect 29748 37865 29776 37896
rect 29914 37884 29920 37896
rect 29972 37884 29978 37936
rect 31294 37924 31300 37936
rect 31234 37896 31300 37924
rect 31294 37884 31300 37896
rect 31352 37884 31358 37936
rect 29733 37859 29791 37865
rect 29733 37825 29745 37859
rect 29779 37825 29791 37859
rect 29733 37819 29791 37825
rect 32030 37816 32036 37868
rect 32088 37816 32094 37868
rect 32416 37856 32444 37964
rect 35158 37952 35164 37964
rect 35216 37952 35222 38004
rect 36722 37952 36728 38004
rect 36780 37992 36786 38004
rect 38657 37995 38715 38001
rect 38657 37992 38669 37995
rect 36780 37964 38669 37992
rect 36780 37952 36786 37964
rect 38657 37961 38669 37964
rect 38703 37961 38715 37995
rect 38657 37955 38715 37961
rect 39114 37952 39120 38004
rect 39172 37952 39178 38004
rect 34422 37924 34428 37936
rect 33994 37896 34428 37924
rect 34422 37884 34428 37896
rect 34480 37884 34486 37936
rect 36446 37884 36452 37936
rect 36504 37924 36510 37936
rect 37829 37927 37887 37933
rect 37829 37924 37841 37927
rect 36504 37896 37841 37924
rect 36504 37884 36510 37896
rect 37829 37893 37841 37896
rect 37875 37893 37887 37927
rect 49234 37924 49240 37936
rect 37829 37887 37887 37893
rect 38120 37896 49240 37924
rect 32493 37859 32551 37865
rect 32493 37856 32505 37859
rect 32416 37828 32505 37856
rect 32493 37825 32505 37828
rect 32539 37825 32551 37859
rect 35621 37859 35679 37865
rect 35621 37856 35633 37859
rect 32493 37819 32551 37825
rect 34164 37828 35633 37856
rect 1302 37748 1308 37800
rect 1360 37788 1366 37800
rect 2041 37791 2099 37797
rect 2041 37788 2053 37791
rect 1360 37760 2053 37788
rect 1360 37748 1366 37760
rect 2041 37757 2053 37760
rect 2087 37757 2099 37791
rect 2041 37751 2099 37757
rect 14829 37791 14887 37797
rect 14829 37757 14841 37791
rect 14875 37788 14887 37791
rect 16114 37788 16120 37800
rect 14875 37760 16120 37788
rect 14875 37757 14887 37760
rect 14829 37751 14887 37757
rect 16114 37748 16120 37760
rect 16172 37748 16178 37800
rect 18417 37791 18475 37797
rect 18417 37757 18429 37791
rect 18463 37757 18475 37791
rect 18417 37751 18475 37757
rect 18601 37791 18659 37797
rect 18601 37757 18613 37791
rect 18647 37788 18659 37791
rect 19334 37788 19340 37800
rect 18647 37760 19340 37788
rect 18647 37757 18659 37760
rect 18601 37751 18659 37757
rect 18432 37720 18460 37751
rect 19334 37748 19340 37760
rect 19392 37748 19398 37800
rect 19426 37748 19432 37800
rect 19484 37748 19490 37800
rect 19518 37748 19524 37800
rect 19576 37748 19582 37800
rect 20438 37748 20444 37800
rect 20496 37788 20502 37800
rect 21269 37791 21327 37797
rect 21269 37788 21281 37791
rect 20496 37760 21281 37788
rect 20496 37748 20502 37760
rect 21269 37757 21281 37760
rect 21315 37757 21327 37791
rect 21269 37751 21327 37757
rect 22281 37791 22339 37797
rect 22281 37757 22293 37791
rect 22327 37788 22339 37791
rect 24029 37791 24087 37797
rect 24029 37788 24041 37791
rect 22327 37760 23336 37788
rect 22327 37757 22339 37760
rect 22281 37751 22339 37757
rect 20070 37720 20076 37732
rect 18432 37692 20076 37720
rect 20070 37680 20076 37692
rect 20128 37680 20134 37732
rect 8570 37612 8576 37664
rect 8628 37612 8634 37664
rect 13814 37612 13820 37664
rect 13872 37652 13878 37664
rect 14918 37652 14924 37664
rect 13872 37624 14924 37652
rect 13872 37612 13878 37624
rect 14918 37612 14924 37624
rect 14976 37652 14982 37664
rect 16301 37655 16359 37661
rect 16301 37652 16313 37655
rect 14976 37624 16313 37652
rect 14976 37612 14982 37624
rect 16301 37621 16313 37624
rect 16347 37621 16359 37655
rect 16301 37615 16359 37621
rect 16482 37612 16488 37664
rect 16540 37652 16546 37664
rect 18969 37655 19027 37661
rect 18969 37652 18981 37655
rect 16540 37624 18981 37652
rect 16540 37612 16546 37624
rect 18969 37621 18981 37624
rect 19015 37621 19027 37655
rect 23308 37652 23336 37760
rect 23400 37760 24041 37788
rect 23400 37732 23428 37760
rect 24029 37757 24041 37760
rect 24075 37757 24087 37791
rect 24029 37751 24087 37757
rect 25038 37748 25044 37800
rect 25096 37748 25102 37800
rect 25222 37748 25228 37800
rect 25280 37788 25286 37800
rect 26145 37791 26203 37797
rect 26145 37788 26157 37791
rect 25280 37760 26157 37788
rect 25280 37748 25286 37760
rect 23382 37680 23388 37732
rect 23440 37680 23446 37732
rect 23474 37680 23480 37732
rect 23532 37720 23538 37732
rect 24489 37723 24547 37729
rect 24489 37720 24501 37723
rect 23532 37692 24501 37720
rect 23532 37680 23538 37692
rect 24489 37689 24501 37692
rect 24535 37689 24547 37723
rect 24489 37683 24547 37689
rect 23842 37652 23848 37664
rect 23308 37624 23848 37652
rect 18969 37615 19027 37621
rect 23842 37612 23848 37624
rect 23900 37612 23906 37664
rect 25792 37652 25820 37760
rect 26145 37757 26157 37760
rect 26191 37757 26203 37791
rect 26145 37751 26203 37757
rect 26237 37791 26295 37797
rect 26237 37757 26249 37791
rect 26283 37757 26295 37791
rect 26237 37751 26295 37757
rect 25866 37680 25872 37732
rect 25924 37720 25930 37732
rect 26252 37720 26280 37751
rect 27062 37748 27068 37800
rect 27120 37788 27126 37800
rect 27433 37791 27491 37797
rect 27433 37788 27445 37791
rect 27120 37760 27445 37788
rect 27120 37748 27126 37760
rect 27433 37757 27445 37760
rect 27479 37757 27491 37791
rect 27433 37751 27491 37757
rect 28166 37748 28172 37800
rect 28224 37788 28230 37800
rect 28626 37788 28632 37800
rect 28224 37760 28632 37788
rect 28224 37748 28230 37760
rect 28626 37748 28632 37760
rect 28684 37748 28690 37800
rect 30009 37791 30067 37797
rect 30009 37757 30021 37791
rect 30055 37788 30067 37791
rect 31846 37788 31852 37800
rect 30055 37760 31852 37788
rect 30055 37757 30067 37760
rect 30009 37751 30067 37757
rect 31846 37748 31852 37760
rect 31904 37748 31910 37800
rect 32048 37720 32076 37816
rect 32769 37791 32827 37797
rect 32769 37757 32781 37791
rect 32815 37788 32827 37791
rect 33778 37788 33784 37800
rect 32815 37760 33784 37788
rect 32815 37757 32827 37760
rect 32769 37751 32827 37757
rect 33778 37748 33784 37760
rect 33836 37748 33842 37800
rect 25924 37692 26280 37720
rect 31036 37692 32076 37720
rect 25924 37680 25930 37692
rect 31036 37652 31064 37692
rect 25792 37624 31064 37652
rect 31110 37612 31116 37664
rect 31168 37652 31174 37664
rect 34164 37652 34192 37828
rect 35621 37825 35633 37828
rect 35667 37825 35679 37859
rect 35621 37819 35679 37825
rect 35434 37788 35440 37800
rect 35360 37760 35440 37788
rect 35253 37723 35311 37729
rect 35253 37689 35265 37723
rect 35299 37720 35311 37723
rect 35360 37720 35388 37760
rect 35434 37748 35440 37760
rect 35492 37748 35498 37800
rect 35299 37692 35388 37720
rect 35636 37720 35664 37819
rect 36998 37816 37004 37868
rect 37056 37856 37062 37868
rect 37921 37859 37979 37865
rect 37921 37856 37933 37859
rect 37056 37828 37933 37856
rect 37056 37816 37062 37828
rect 37921 37825 37933 37828
rect 37967 37825 37979 37859
rect 37921 37819 37979 37825
rect 35710 37748 35716 37800
rect 35768 37748 35774 37800
rect 35802 37748 35808 37800
rect 35860 37748 35866 37800
rect 37826 37748 37832 37800
rect 37884 37788 37890 37800
rect 38013 37791 38071 37797
rect 38013 37788 38025 37791
rect 37884 37760 38025 37788
rect 37884 37748 37890 37760
rect 38013 37757 38025 37760
rect 38059 37757 38071 37791
rect 38013 37751 38071 37757
rect 38120 37720 38148 37896
rect 49234 37884 49240 37896
rect 49292 37884 49298 37936
rect 39025 37859 39083 37865
rect 39025 37825 39037 37859
rect 39071 37856 39083 37859
rect 39071 37828 45554 37856
rect 39071 37825 39083 37828
rect 39025 37819 39083 37825
rect 38562 37748 38568 37800
rect 38620 37788 38626 37800
rect 39209 37791 39267 37797
rect 39209 37788 39221 37791
rect 38620 37760 39221 37788
rect 38620 37748 38626 37760
rect 39209 37757 39221 37760
rect 39255 37757 39267 37791
rect 39209 37751 39267 37757
rect 35636 37692 38148 37720
rect 45526 37720 45554 37828
rect 49326 37816 49332 37868
rect 49384 37816 49390 37868
rect 49145 37723 49203 37729
rect 49145 37720 49157 37723
rect 45526 37692 49157 37720
rect 35299 37689 35311 37692
rect 35253 37683 35311 37689
rect 49145 37689 49157 37692
rect 49191 37689 49203 37723
rect 49145 37683 49203 37689
rect 31168 37624 34192 37652
rect 31168 37612 31174 37624
rect 34238 37612 34244 37664
rect 34296 37612 34302 37664
rect 34698 37612 34704 37664
rect 34756 37652 34762 37664
rect 35710 37652 35716 37664
rect 34756 37624 35716 37652
rect 34756 37612 34762 37624
rect 35710 37612 35716 37624
rect 35768 37612 35774 37664
rect 37461 37655 37519 37661
rect 37461 37621 37473 37655
rect 37507 37652 37519 37655
rect 39850 37652 39856 37664
rect 37507 37624 39856 37652
rect 37507 37621 37519 37624
rect 37461 37615 37519 37621
rect 39850 37612 39856 37624
rect 39908 37612 39914 37664
rect 1104 37562 49864 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 32950 37562
rect 33002 37510 33014 37562
rect 33066 37510 33078 37562
rect 33130 37510 33142 37562
rect 33194 37510 33206 37562
rect 33258 37510 42950 37562
rect 43002 37510 43014 37562
rect 43066 37510 43078 37562
rect 43130 37510 43142 37562
rect 43194 37510 43206 37562
rect 43258 37510 49864 37562
rect 1104 37488 49864 37510
rect 14366 37408 14372 37460
rect 14424 37448 14430 37460
rect 14424 37420 18552 37448
rect 14424 37408 14430 37420
rect 12986 37272 12992 37324
rect 13044 37312 13050 37324
rect 13633 37315 13691 37321
rect 13633 37312 13645 37315
rect 13044 37284 13645 37312
rect 13044 37272 13050 37284
rect 13633 37281 13645 37284
rect 13679 37281 13691 37315
rect 13633 37275 13691 37281
rect 12526 37204 12532 37256
rect 12584 37244 12590 37256
rect 13357 37247 13415 37253
rect 13357 37244 13369 37247
rect 12584 37216 13369 37244
rect 12584 37204 12590 37216
rect 13357 37213 13369 37216
rect 13403 37213 13415 37247
rect 13648 37244 13676 37275
rect 14642 37272 14648 37324
rect 14700 37312 14706 37324
rect 14921 37315 14979 37321
rect 14921 37312 14933 37315
rect 14700 37284 14933 37312
rect 14700 37272 14706 37284
rect 14921 37281 14933 37284
rect 14967 37281 14979 37315
rect 14921 37275 14979 37281
rect 15102 37272 15108 37324
rect 15160 37272 15166 37324
rect 16117 37315 16175 37321
rect 16117 37281 16129 37315
rect 16163 37312 16175 37315
rect 16206 37312 16212 37324
rect 16163 37284 16212 37312
rect 16163 37281 16175 37284
rect 16117 37275 16175 37281
rect 16206 37272 16212 37284
rect 16264 37312 16270 37324
rect 18414 37312 18420 37324
rect 16264 37284 18420 37312
rect 16264 37272 16270 37284
rect 18414 37272 18420 37284
rect 18472 37272 18478 37324
rect 18524 37312 18552 37420
rect 20990 37408 20996 37460
rect 21048 37448 21054 37460
rect 21729 37451 21787 37457
rect 21729 37448 21741 37451
rect 21048 37420 21741 37448
rect 21048 37408 21054 37420
rect 21729 37417 21741 37420
rect 21775 37417 21787 37451
rect 28258 37448 28264 37460
rect 21729 37411 21787 37417
rect 22066 37420 28264 37448
rect 18874 37340 18880 37392
rect 18932 37380 18938 37392
rect 22066 37380 22094 37420
rect 28258 37408 28264 37420
rect 28316 37448 28322 37460
rect 31110 37448 31116 37460
rect 28316 37420 31116 37448
rect 28316 37408 28322 37420
rect 31110 37408 31116 37420
rect 31168 37408 31174 37460
rect 31294 37408 31300 37460
rect 31352 37448 31358 37460
rect 31352 37420 32260 37448
rect 31352 37408 31358 37420
rect 18932 37352 22094 37380
rect 18932 37340 18938 37352
rect 18601 37315 18659 37321
rect 18601 37312 18613 37315
rect 18524 37284 18613 37312
rect 18601 37281 18613 37284
rect 18647 37312 18659 37315
rect 19242 37312 19248 37324
rect 18647 37284 19248 37312
rect 18647 37281 18659 37284
rect 18601 37275 18659 37281
rect 19242 37272 19248 37284
rect 19300 37272 19306 37324
rect 20349 37315 20407 37321
rect 20349 37281 20361 37315
rect 20395 37312 20407 37315
rect 22370 37312 22376 37324
rect 20395 37284 22376 37312
rect 20395 37281 20407 37284
rect 20349 37275 20407 37281
rect 22370 37272 22376 37284
rect 22428 37272 22434 37324
rect 23569 37315 23627 37321
rect 23569 37281 23581 37315
rect 23615 37312 23627 37315
rect 23934 37312 23940 37324
rect 23615 37284 23940 37312
rect 23615 37281 23627 37284
rect 23569 37275 23627 37281
rect 23934 37272 23940 37284
rect 23992 37272 23998 37324
rect 24026 37272 24032 37324
rect 24084 37312 24090 37324
rect 26789 37315 26847 37321
rect 26789 37312 26801 37315
rect 24084 37284 26801 37312
rect 24084 37272 24090 37284
rect 26789 37281 26801 37284
rect 26835 37281 26847 37315
rect 26789 37275 26847 37281
rect 27062 37272 27068 37324
rect 27120 37312 27126 37324
rect 28350 37312 28356 37324
rect 27120 37284 28356 37312
rect 27120 37272 27126 37284
rect 28350 37272 28356 37284
rect 28408 37312 28414 37324
rect 28408 37284 28948 37312
rect 28408 37272 28414 37284
rect 13906 37244 13912 37256
rect 13648 37216 13912 37244
rect 13357 37207 13415 37213
rect 13906 37204 13912 37216
rect 13964 37204 13970 37256
rect 14458 37204 14464 37256
rect 14516 37244 14522 37256
rect 15838 37244 15844 37256
rect 14516 37216 15844 37244
rect 14516 37204 14522 37216
rect 15838 37204 15844 37216
rect 15896 37204 15902 37256
rect 17586 37204 17592 37256
rect 17644 37204 17650 37256
rect 20073 37247 20131 37253
rect 20073 37213 20085 37247
rect 20119 37244 20131 37247
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 20119 37216 21097 37244
rect 20119 37213 20131 37216
rect 20073 37207 20131 37213
rect 21085 37213 21097 37216
rect 21131 37213 21143 37247
rect 21085 37207 21143 37213
rect 23290 37204 23296 37256
rect 23348 37244 23354 37256
rect 23385 37247 23443 37253
rect 23385 37244 23397 37247
rect 23348 37216 23397 37244
rect 23348 37204 23354 37216
rect 23385 37213 23397 37216
rect 23431 37213 23443 37247
rect 23385 37207 23443 37213
rect 27433 37247 27491 37253
rect 27433 37213 27445 37247
rect 27479 37244 27491 37247
rect 27614 37244 27620 37256
rect 27479 37216 27620 37244
rect 27479 37213 27491 37216
rect 27433 37207 27491 37213
rect 27614 37204 27620 37216
rect 27672 37204 27678 37256
rect 5350 37136 5356 37188
rect 5408 37176 5414 37188
rect 13449 37179 13507 37185
rect 13449 37176 13461 37179
rect 5408 37148 13461 37176
rect 5408 37136 5414 37148
rect 13449 37145 13461 37148
rect 13495 37145 13507 37179
rect 15746 37176 15752 37188
rect 13449 37139 13507 37145
rect 14384 37148 15752 37176
rect 12989 37111 13047 37117
rect 12989 37077 13001 37111
rect 13035 37108 13047 37111
rect 14384 37108 14412 37148
rect 15746 37136 15752 37148
rect 15804 37136 15810 37188
rect 16666 37136 16672 37188
rect 16724 37136 16730 37188
rect 17604 37176 17632 37204
rect 18417 37179 18475 37185
rect 18417 37176 18429 37179
rect 17604 37148 18429 37176
rect 18417 37145 18429 37148
rect 18463 37145 18475 37179
rect 18417 37139 18475 37145
rect 19886 37136 19892 37188
rect 19944 37176 19950 37188
rect 19944 37148 22094 37176
rect 19944 37136 19950 37148
rect 13035 37080 14412 37108
rect 14461 37111 14519 37117
rect 13035 37077 13047 37080
rect 12989 37071 13047 37077
rect 14461 37077 14473 37111
rect 14507 37108 14519 37111
rect 14734 37108 14740 37120
rect 14507 37080 14740 37108
rect 14507 37077 14519 37080
rect 14461 37071 14519 37077
rect 14734 37068 14740 37080
rect 14792 37068 14798 37120
rect 14829 37111 14887 37117
rect 14829 37077 14841 37111
rect 14875 37108 14887 37111
rect 15010 37108 15016 37120
rect 14875 37080 15016 37108
rect 14875 37077 14887 37080
rect 14829 37071 14887 37077
rect 15010 37068 15016 37080
rect 15068 37068 15074 37120
rect 16206 37068 16212 37120
rect 16264 37108 16270 37120
rect 17589 37111 17647 37117
rect 17589 37108 17601 37111
rect 16264 37080 17601 37108
rect 16264 37068 16270 37080
rect 17589 37077 17601 37080
rect 17635 37077 17647 37111
rect 17589 37071 17647 37077
rect 17678 37068 17684 37120
rect 17736 37108 17742 37120
rect 18049 37111 18107 37117
rect 18049 37108 18061 37111
rect 17736 37080 18061 37108
rect 17736 37068 17742 37080
rect 18049 37077 18061 37080
rect 18095 37077 18107 37111
rect 18049 37071 18107 37077
rect 18509 37111 18567 37117
rect 18509 37077 18521 37111
rect 18555 37108 18567 37111
rect 18782 37108 18788 37120
rect 18555 37080 18788 37108
rect 18555 37077 18567 37080
rect 18509 37071 18567 37077
rect 18782 37068 18788 37080
rect 18840 37068 18846 37120
rect 19705 37111 19763 37117
rect 19705 37077 19717 37111
rect 19751 37108 19763 37111
rect 19794 37108 19800 37120
rect 19751 37080 19800 37108
rect 19751 37077 19763 37080
rect 19705 37071 19763 37077
rect 19794 37068 19800 37080
rect 19852 37068 19858 37120
rect 20165 37111 20223 37117
rect 20165 37077 20177 37111
rect 20211 37108 20223 37111
rect 21726 37108 21732 37120
rect 20211 37080 21732 37108
rect 20211 37077 20223 37080
rect 20165 37071 20223 37077
rect 21726 37068 21732 37080
rect 21784 37068 21790 37120
rect 22066 37108 22094 37148
rect 26050 37136 26056 37188
rect 26108 37176 26114 37188
rect 26108 37148 26556 37176
rect 26108 37136 26114 37148
rect 26528 37120 26556 37148
rect 27522 37136 27528 37188
rect 27580 37176 27586 37188
rect 28169 37179 28227 37185
rect 28169 37176 28181 37179
rect 27580 37148 28181 37176
rect 27580 37136 27586 37148
rect 28169 37145 28181 37148
rect 28215 37145 28227 37179
rect 28920 37176 28948 37284
rect 30006 37272 30012 37324
rect 30064 37312 30070 37324
rect 30926 37312 30932 37324
rect 30064 37284 30932 37312
rect 30064 37272 30070 37284
rect 30926 37272 30932 37284
rect 30984 37272 30990 37324
rect 32232 37312 32260 37420
rect 33410 37408 33416 37460
rect 33468 37448 33474 37460
rect 34241 37451 34299 37457
rect 34241 37448 34253 37451
rect 33468 37420 34253 37448
rect 33468 37408 33474 37420
rect 34241 37417 34253 37420
rect 34287 37417 34299 37451
rect 34241 37411 34299 37417
rect 32232 37284 32444 37312
rect 29914 37204 29920 37256
rect 29972 37244 29978 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 29972 37216 30665 37244
rect 29972 37204 29978 37216
rect 30653 37213 30665 37216
rect 30699 37213 30711 37247
rect 32232 37244 32260 37284
rect 32062 37216 32260 37244
rect 30653 37207 30711 37213
rect 30466 37176 30472 37188
rect 28920 37148 30472 37176
rect 28169 37139 28227 37145
rect 30466 37136 30472 37148
rect 30524 37136 30530 37188
rect 22925 37111 22983 37117
rect 22925 37108 22937 37111
rect 22066 37080 22937 37108
rect 22925 37077 22937 37080
rect 22971 37077 22983 37111
rect 22925 37071 22983 37077
rect 23290 37068 23296 37120
rect 23348 37068 23354 37120
rect 26234 37068 26240 37120
rect 26292 37068 26298 37120
rect 26510 37068 26516 37120
rect 26568 37108 26574 37120
rect 26605 37111 26663 37117
rect 26605 37108 26617 37111
rect 26568 37080 26617 37108
rect 26568 37068 26574 37080
rect 26605 37077 26617 37080
rect 26651 37077 26663 37111
rect 26605 37071 26663 37077
rect 26697 37111 26755 37117
rect 26697 37077 26709 37111
rect 26743 37108 26755 37111
rect 30374 37108 30380 37120
rect 26743 37080 30380 37108
rect 26743 37077 26755 37080
rect 26697 37071 26755 37077
rect 30374 37068 30380 37080
rect 30432 37068 30438 37120
rect 30668 37108 30696 37207
rect 32306 37204 32312 37256
rect 32364 37204 32370 37256
rect 32416 37244 32444 37284
rect 33318 37272 33324 37324
rect 33376 37312 33382 37324
rect 33413 37315 33471 37321
rect 33413 37312 33425 37315
rect 33376 37284 33425 37312
rect 33376 37272 33382 37284
rect 33413 37281 33425 37284
rect 33459 37281 33471 37315
rect 33413 37275 33471 37281
rect 35621 37315 35679 37321
rect 35621 37281 35633 37315
rect 35667 37312 35679 37315
rect 36814 37312 36820 37324
rect 35667 37284 36820 37312
rect 35667 37281 35679 37284
rect 35621 37275 35679 37281
rect 36814 37272 36820 37284
rect 36872 37272 36878 37324
rect 36906 37272 36912 37324
rect 36964 37312 36970 37324
rect 38105 37315 38163 37321
rect 38105 37312 38117 37315
rect 36964 37284 38117 37312
rect 36964 37272 36970 37284
rect 38105 37281 38117 37284
rect 38151 37281 38163 37315
rect 38105 37275 38163 37281
rect 33134 37244 33140 37256
rect 32416 37216 33140 37244
rect 33134 37204 33140 37216
rect 33192 37204 33198 37256
rect 34146 37204 34152 37256
rect 34204 37244 34210 37256
rect 35345 37247 35403 37253
rect 35345 37244 35357 37247
rect 34204 37216 35357 37244
rect 34204 37204 34210 37216
rect 35345 37213 35357 37216
rect 35391 37213 35403 37247
rect 35345 37207 35403 37213
rect 37642 37204 37648 37256
rect 37700 37244 37706 37256
rect 37921 37247 37979 37253
rect 37921 37244 37933 37247
rect 37700 37216 37933 37244
rect 37700 37204 37706 37216
rect 37921 37213 37933 37216
rect 37967 37213 37979 37247
rect 37921 37207 37979 37213
rect 32324 37176 32352 37204
rect 32766 37176 32772 37188
rect 32324 37148 32772 37176
rect 32306 37108 32312 37120
rect 30668 37080 32312 37108
rect 32306 37068 32312 37080
rect 32364 37068 32370 37120
rect 32416 37117 32444 37148
rect 32766 37136 32772 37148
rect 32824 37136 32830 37188
rect 33229 37179 33287 37185
rect 33229 37145 33241 37179
rect 33275 37176 33287 37179
rect 33410 37176 33416 37188
rect 33275 37148 33416 37176
rect 33275 37145 33287 37148
rect 33229 37139 33287 37145
rect 33410 37136 33416 37148
rect 33468 37136 33474 37188
rect 36354 37136 36360 37188
rect 36412 37136 36418 37188
rect 38654 37176 38660 37188
rect 37108 37148 38660 37176
rect 32401 37111 32459 37117
rect 32401 37077 32413 37111
rect 32447 37077 32459 37111
rect 32401 37071 32459 37077
rect 32490 37068 32496 37120
rect 32548 37108 32554 37120
rect 32861 37111 32919 37117
rect 32861 37108 32873 37111
rect 32548 37080 32873 37108
rect 32548 37068 32554 37080
rect 32861 37077 32873 37080
rect 32907 37077 32919 37111
rect 32861 37071 32919 37077
rect 33321 37111 33379 37117
rect 33321 37077 33333 37111
rect 33367 37108 33379 37111
rect 35802 37108 35808 37120
rect 33367 37080 35808 37108
rect 33367 37077 33379 37080
rect 33321 37071 33379 37077
rect 35802 37068 35808 37080
rect 35860 37068 35866 37120
rect 37108 37117 37136 37148
rect 38654 37136 38660 37148
rect 38712 37176 38718 37188
rect 39390 37176 39396 37188
rect 38712 37148 39396 37176
rect 38712 37136 38718 37148
rect 39390 37136 39396 37148
rect 39448 37136 39454 37188
rect 37093 37111 37151 37117
rect 37093 37077 37105 37111
rect 37139 37077 37151 37111
rect 37093 37071 37151 37077
rect 37550 37068 37556 37120
rect 37608 37068 37614 37120
rect 37642 37068 37648 37120
rect 37700 37108 37706 37120
rect 38013 37111 38071 37117
rect 38013 37108 38025 37111
rect 37700 37080 38025 37108
rect 37700 37068 37706 37080
rect 38013 37077 38025 37080
rect 38059 37077 38071 37111
rect 38013 37071 38071 37077
rect 1104 37018 49864 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 27950 37018
rect 28002 36966 28014 37018
rect 28066 36966 28078 37018
rect 28130 36966 28142 37018
rect 28194 36966 28206 37018
rect 28258 36966 37950 37018
rect 38002 36966 38014 37018
rect 38066 36966 38078 37018
rect 38130 36966 38142 37018
rect 38194 36966 38206 37018
rect 38258 36966 47950 37018
rect 48002 36966 48014 37018
rect 48066 36966 48078 37018
rect 48130 36966 48142 37018
rect 48194 36966 48206 37018
rect 48258 36966 49864 37018
rect 1104 36944 49864 36966
rect 12710 36864 12716 36916
rect 12768 36904 12774 36916
rect 12805 36907 12863 36913
rect 12805 36904 12817 36907
rect 12768 36876 12817 36904
rect 12768 36864 12774 36876
rect 12805 36873 12817 36876
rect 12851 36904 12863 36907
rect 13446 36904 13452 36916
rect 12851 36876 13452 36904
rect 12851 36873 12863 36876
rect 12805 36867 12863 36873
rect 13446 36864 13452 36876
rect 13504 36864 13510 36916
rect 14458 36904 14464 36916
rect 13648 36876 14464 36904
rect 13648 36836 13676 36876
rect 14458 36864 14464 36876
rect 14516 36864 14522 36916
rect 18506 36864 18512 36916
rect 18564 36904 18570 36916
rect 18601 36907 18659 36913
rect 18601 36904 18613 36907
rect 18564 36876 18613 36904
rect 18564 36864 18570 36876
rect 18601 36873 18613 36876
rect 18647 36873 18659 36907
rect 18601 36867 18659 36873
rect 19058 36864 19064 36916
rect 19116 36904 19122 36916
rect 19521 36907 19579 36913
rect 19116 36876 19472 36904
rect 19116 36864 19122 36876
rect 13556 36808 13676 36836
rect 1762 36728 1768 36780
rect 1820 36728 1826 36780
rect 4890 36728 4896 36780
rect 4948 36768 4954 36780
rect 5350 36768 5356 36780
rect 4948 36740 5356 36768
rect 4948 36728 4954 36740
rect 5350 36728 5356 36740
rect 5408 36728 5414 36780
rect 12713 36771 12771 36777
rect 12713 36737 12725 36771
rect 12759 36768 12771 36771
rect 13446 36768 13452 36780
rect 12759 36740 13452 36768
rect 12759 36737 12771 36740
rect 12713 36731 12771 36737
rect 13446 36728 13452 36740
rect 13504 36728 13510 36780
rect 13556 36777 13584 36808
rect 13814 36796 13820 36848
rect 13872 36796 13878 36848
rect 16666 36836 16672 36848
rect 16224 36808 16672 36836
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36737 13599 36771
rect 13541 36731 13599 36737
rect 14918 36728 14924 36780
rect 14976 36768 14982 36780
rect 16224 36768 16252 36808
rect 16666 36796 16672 36808
rect 16724 36836 16730 36848
rect 19444 36836 19472 36876
rect 19521 36873 19533 36907
rect 19567 36904 19579 36907
rect 19610 36904 19616 36916
rect 19567 36876 19616 36904
rect 19567 36873 19579 36876
rect 19521 36867 19579 36873
rect 19610 36864 19616 36876
rect 19668 36864 19674 36916
rect 21085 36907 21143 36913
rect 21085 36873 21097 36907
rect 21131 36904 21143 36907
rect 22186 36904 22192 36916
rect 21131 36876 22192 36904
rect 21131 36873 21143 36876
rect 21085 36867 21143 36873
rect 22186 36864 22192 36876
rect 22244 36864 22250 36916
rect 22465 36907 22523 36913
rect 22465 36873 22477 36907
rect 22511 36904 22523 36907
rect 26234 36904 26240 36916
rect 22511 36876 26240 36904
rect 22511 36873 22523 36876
rect 22465 36867 22523 36873
rect 26234 36864 26240 36876
rect 26292 36864 26298 36916
rect 26344 36876 29224 36904
rect 20806 36836 20812 36848
rect 16724 36808 17618 36836
rect 18524 36808 19380 36836
rect 19444 36808 20812 36836
rect 16724 36796 16730 36808
rect 18524 36780 18552 36808
rect 14976 36740 16252 36768
rect 16301 36771 16359 36777
rect 14976 36728 14982 36740
rect 16301 36737 16313 36771
rect 16347 36768 16359 36771
rect 16758 36768 16764 36780
rect 16347 36740 16764 36768
rect 16347 36737 16359 36740
rect 16301 36731 16359 36737
rect 16758 36728 16764 36740
rect 16816 36728 16822 36780
rect 18506 36728 18512 36780
rect 18564 36728 18570 36780
rect 19352 36768 19380 36808
rect 20806 36796 20812 36808
rect 20864 36796 20870 36848
rect 22002 36796 22008 36848
rect 22060 36836 22066 36848
rect 22060 36808 23612 36836
rect 22060 36796 22066 36808
rect 19429 36771 19487 36777
rect 19429 36768 19441 36771
rect 19352 36740 19441 36768
rect 19429 36737 19441 36740
rect 19475 36737 19487 36771
rect 19429 36731 19487 36737
rect 21818 36728 21824 36780
rect 21876 36768 21882 36780
rect 23584 36777 23612 36808
rect 24394 36796 24400 36848
rect 24452 36796 24458 36848
rect 26344 36836 26372 36876
rect 27706 36836 27712 36848
rect 25148 36808 26372 36836
rect 26436 36808 27712 36836
rect 22373 36771 22431 36777
rect 22373 36768 22385 36771
rect 21876 36740 22385 36768
rect 21876 36728 21882 36740
rect 22373 36737 22385 36740
rect 22419 36737 22431 36771
rect 22373 36731 22431 36737
rect 23569 36771 23627 36777
rect 23569 36737 23581 36771
rect 23615 36737 23627 36771
rect 25148 36768 25176 36808
rect 23569 36731 23627 36737
rect 25056 36740 25176 36768
rect 1302 36660 1308 36712
rect 1360 36700 1366 36712
rect 2041 36703 2099 36709
rect 2041 36700 2053 36703
rect 1360 36672 2053 36700
rect 1360 36660 1366 36672
rect 2041 36669 2053 36672
rect 2087 36669 2099 36703
rect 2041 36663 2099 36669
rect 12986 36660 12992 36712
rect 13044 36660 13050 36712
rect 13354 36660 13360 36712
rect 13412 36700 13418 36712
rect 13412 36672 14872 36700
rect 13412 36660 13418 36672
rect 14844 36632 14872 36672
rect 15838 36660 15844 36712
rect 15896 36700 15902 36712
rect 16850 36700 16856 36712
rect 15896 36672 16856 36700
rect 15896 36660 15902 36672
rect 16850 36660 16856 36672
rect 16908 36660 16914 36712
rect 17126 36660 17132 36712
rect 17184 36660 17190 36712
rect 19242 36660 19248 36712
rect 19300 36700 19306 36712
rect 19705 36703 19763 36709
rect 19705 36700 19717 36703
rect 19300 36672 19717 36700
rect 19300 36660 19306 36672
rect 19705 36669 19717 36672
rect 19751 36700 19763 36703
rect 19794 36700 19800 36712
rect 19751 36672 19800 36700
rect 19751 36669 19763 36672
rect 19705 36663 19763 36669
rect 19794 36660 19800 36672
rect 19852 36660 19858 36712
rect 21174 36660 21180 36712
rect 21232 36660 21238 36712
rect 21358 36660 21364 36712
rect 21416 36660 21422 36712
rect 22646 36660 22652 36712
rect 22704 36660 22710 36712
rect 22738 36660 22744 36712
rect 22796 36700 22802 36712
rect 23842 36700 23848 36712
rect 22796 36672 23848 36700
rect 22796 36660 22802 36672
rect 23842 36660 23848 36672
rect 23900 36660 23906 36712
rect 24578 36660 24584 36712
rect 24636 36700 24642 36712
rect 25056 36700 25084 36740
rect 25222 36728 25228 36780
rect 25280 36768 25286 36780
rect 26145 36771 26203 36777
rect 26145 36768 26157 36771
rect 25280 36740 26157 36768
rect 25280 36728 25286 36740
rect 26145 36737 26157 36740
rect 26191 36737 26203 36771
rect 26145 36731 26203 36737
rect 26237 36771 26295 36777
rect 26237 36737 26249 36771
rect 26283 36768 26295 36771
rect 26436 36768 26464 36808
rect 27706 36796 27712 36808
rect 27764 36796 27770 36848
rect 28166 36796 28172 36848
rect 28224 36796 28230 36848
rect 29196 36845 29224 36876
rect 30742 36864 30748 36916
rect 30800 36904 30806 36916
rect 32674 36904 32680 36916
rect 30800 36876 32680 36904
rect 30800 36864 30806 36876
rect 32674 36864 32680 36876
rect 32732 36864 32738 36916
rect 33502 36864 33508 36916
rect 33560 36904 33566 36916
rect 34149 36907 34207 36913
rect 33560 36876 34100 36904
rect 33560 36864 33566 36876
rect 29181 36839 29239 36845
rect 29181 36805 29193 36839
rect 29227 36805 29239 36839
rect 29914 36836 29920 36848
rect 29181 36799 29239 36805
rect 29656 36808 29920 36836
rect 26283 36740 26464 36768
rect 26283 36737 26295 36740
rect 26237 36731 26295 36737
rect 24636 36672 25084 36700
rect 24636 36660 24642 36672
rect 25130 36660 25136 36712
rect 25188 36700 25194 36712
rect 25317 36703 25375 36709
rect 25317 36700 25329 36703
rect 25188 36672 25329 36700
rect 25188 36660 25194 36672
rect 25317 36669 25329 36672
rect 25363 36700 25375 36703
rect 25958 36700 25964 36712
rect 25363 36672 25964 36700
rect 25363 36669 25375 36672
rect 25317 36663 25375 36669
rect 25958 36660 25964 36672
rect 26016 36660 26022 36712
rect 26050 36660 26056 36712
rect 26108 36700 26114 36712
rect 26252 36700 26280 36731
rect 27154 36728 27160 36780
rect 27212 36728 27218 36780
rect 29656 36777 29684 36808
rect 29914 36796 29920 36808
rect 29972 36796 29978 36848
rect 31294 36836 31300 36848
rect 31142 36808 31300 36836
rect 31294 36796 31300 36808
rect 31352 36796 31358 36848
rect 34072 36836 34100 36876
rect 34149 36873 34161 36907
rect 34195 36904 34207 36907
rect 35342 36904 35348 36916
rect 34195 36876 35348 36904
rect 34195 36873 34207 36876
rect 34149 36867 34207 36873
rect 35342 36864 35348 36876
rect 35400 36864 35406 36916
rect 36725 36907 36783 36913
rect 36725 36873 36737 36907
rect 36771 36904 36783 36907
rect 36814 36904 36820 36916
rect 36771 36876 36820 36904
rect 36771 36873 36783 36876
rect 36725 36867 36783 36873
rect 36814 36864 36820 36876
rect 36872 36864 36878 36916
rect 38746 36864 38752 36916
rect 38804 36864 38810 36916
rect 35253 36839 35311 36845
rect 35253 36836 35265 36839
rect 34072 36808 35265 36836
rect 35253 36805 35265 36808
rect 35299 36805 35311 36839
rect 35253 36799 35311 36805
rect 36538 36796 36544 36848
rect 36596 36836 36602 36848
rect 49234 36836 49240 36848
rect 36596 36808 49240 36836
rect 36596 36796 36602 36808
rect 49234 36796 49240 36808
rect 49292 36796 49298 36848
rect 29641 36771 29699 36777
rect 29641 36737 29653 36771
rect 29687 36737 29699 36771
rect 34422 36768 34428 36780
rect 33810 36754 34428 36768
rect 29641 36731 29699 36737
rect 33796 36740 34428 36754
rect 26108 36672 26280 36700
rect 26329 36703 26387 36709
rect 26108 36660 26114 36672
rect 26329 36669 26341 36703
rect 26375 36669 26387 36703
rect 26329 36663 26387 36669
rect 27433 36703 27491 36709
rect 27433 36669 27445 36703
rect 27479 36700 27491 36703
rect 27798 36700 27804 36712
rect 27479 36672 27804 36700
rect 27479 36669 27491 36672
rect 27433 36663 27491 36669
rect 16117 36635 16175 36641
rect 16117 36632 16129 36635
rect 14844 36604 16129 36632
rect 16117 36601 16129 36604
rect 16163 36601 16175 36635
rect 19061 36635 19119 36641
rect 19061 36632 19073 36635
rect 16117 36595 16175 36601
rect 18708 36604 19073 36632
rect 12345 36567 12403 36573
rect 12345 36533 12357 36567
rect 12391 36564 12403 36567
rect 15194 36564 15200 36576
rect 12391 36536 15200 36564
rect 12391 36533 12403 36536
rect 12345 36527 12403 36533
rect 15194 36524 15200 36536
rect 15252 36524 15258 36576
rect 15286 36524 15292 36576
rect 15344 36524 15350 36576
rect 16482 36524 16488 36576
rect 16540 36564 16546 36576
rect 18708 36564 18736 36604
rect 19061 36601 19073 36604
rect 19107 36601 19119 36635
rect 20717 36635 20775 36641
rect 20717 36632 20729 36635
rect 19061 36595 19119 36601
rect 19260 36604 20729 36632
rect 19260 36576 19288 36604
rect 20717 36601 20729 36604
rect 20763 36601 20775 36635
rect 20717 36595 20775 36601
rect 26142 36592 26148 36644
rect 26200 36632 26206 36644
rect 26344 36632 26372 36663
rect 27798 36660 27804 36672
rect 27856 36660 27862 36712
rect 29917 36703 29975 36709
rect 29917 36669 29929 36703
rect 29963 36700 29975 36703
rect 30282 36700 30288 36712
rect 29963 36672 30288 36700
rect 29963 36669 29975 36672
rect 29917 36663 29975 36669
rect 30282 36660 30288 36672
rect 30340 36660 30346 36712
rect 30466 36660 30472 36712
rect 30524 36700 30530 36712
rect 31389 36703 31447 36709
rect 31389 36700 31401 36703
rect 30524 36672 31401 36700
rect 30524 36660 30530 36672
rect 31389 36669 31401 36672
rect 31435 36669 31447 36703
rect 31389 36663 31447 36669
rect 32398 36660 32404 36712
rect 32456 36660 32462 36712
rect 32677 36703 32735 36709
rect 32677 36669 32689 36703
rect 32723 36700 32735 36703
rect 32766 36700 32772 36712
rect 32723 36672 32772 36700
rect 32723 36669 32735 36672
rect 32677 36663 32735 36669
rect 32766 36660 32772 36672
rect 32824 36660 32830 36712
rect 33134 36660 33140 36712
rect 33192 36700 33198 36712
rect 33796 36700 33824 36740
rect 34422 36728 34428 36740
rect 34480 36728 34486 36780
rect 36354 36728 36360 36780
rect 36412 36728 36418 36780
rect 38657 36771 38715 36777
rect 38657 36737 38669 36771
rect 38703 36768 38715 36771
rect 47394 36768 47400 36780
rect 38703 36740 47400 36768
rect 38703 36737 38715 36740
rect 38657 36731 38715 36737
rect 47394 36728 47400 36740
rect 47452 36728 47458 36780
rect 49050 36728 49056 36780
rect 49108 36728 49114 36780
rect 33192 36672 33824 36700
rect 33192 36660 33198 36672
rect 34146 36660 34152 36712
rect 34204 36700 34210 36712
rect 34977 36703 35035 36709
rect 34977 36700 34989 36703
rect 34204 36672 34989 36700
rect 34204 36660 34210 36672
rect 34977 36669 34989 36672
rect 35023 36669 35035 36703
rect 34977 36663 35035 36669
rect 38838 36660 38844 36712
rect 38896 36660 38902 36712
rect 26200 36604 26372 36632
rect 26200 36592 26206 36604
rect 48314 36592 48320 36644
rect 48372 36632 48378 36644
rect 49237 36635 49295 36641
rect 49237 36632 49249 36635
rect 48372 36604 49249 36632
rect 48372 36592 48378 36604
rect 49237 36601 49249 36604
rect 49283 36601 49295 36635
rect 49237 36595 49295 36601
rect 16540 36536 18736 36564
rect 16540 36524 16546 36536
rect 19242 36524 19248 36576
rect 19300 36524 19306 36576
rect 21910 36524 21916 36576
rect 21968 36564 21974 36576
rect 22005 36567 22063 36573
rect 22005 36564 22017 36567
rect 21968 36536 22017 36564
rect 21968 36524 21974 36536
rect 22005 36533 22017 36536
rect 22051 36533 22063 36567
rect 22005 36527 22063 36533
rect 22554 36524 22560 36576
rect 22612 36564 22618 36576
rect 22738 36564 22744 36576
rect 22612 36536 22744 36564
rect 22612 36524 22618 36536
rect 22738 36524 22744 36536
rect 22796 36524 22802 36576
rect 25777 36567 25835 36573
rect 25777 36533 25789 36567
rect 25823 36564 25835 36567
rect 30098 36564 30104 36576
rect 25823 36536 30104 36564
rect 25823 36533 25835 36536
rect 25777 36527 25835 36533
rect 30098 36524 30104 36536
rect 30156 36524 30162 36576
rect 32214 36524 32220 36576
rect 32272 36564 32278 36576
rect 34698 36564 34704 36576
rect 32272 36536 34704 36564
rect 32272 36524 32278 36536
rect 34698 36524 34704 36536
rect 34756 36524 34762 36576
rect 35066 36524 35072 36576
rect 35124 36564 35130 36576
rect 38289 36567 38347 36573
rect 38289 36564 38301 36567
rect 35124 36536 38301 36564
rect 35124 36524 35130 36536
rect 38289 36533 38301 36536
rect 38335 36533 38347 36567
rect 38289 36527 38347 36533
rect 1104 36474 49864 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 32950 36474
rect 33002 36422 33014 36474
rect 33066 36422 33078 36474
rect 33130 36422 33142 36474
rect 33194 36422 33206 36474
rect 33258 36422 42950 36474
rect 43002 36422 43014 36474
rect 43066 36422 43078 36474
rect 43130 36422 43142 36474
rect 43194 36422 43206 36474
rect 43258 36422 49864 36474
rect 1104 36400 49864 36422
rect 1762 36320 1768 36372
rect 1820 36360 1826 36372
rect 8481 36363 8539 36369
rect 8481 36360 8493 36363
rect 1820 36332 8493 36360
rect 1820 36320 1826 36332
rect 8481 36329 8493 36332
rect 8527 36329 8539 36363
rect 8481 36323 8539 36329
rect 9125 36363 9183 36369
rect 9125 36329 9137 36363
rect 9171 36360 9183 36363
rect 11790 36360 11796 36372
rect 9171 36332 11796 36360
rect 9171 36329 9183 36332
rect 9125 36323 9183 36329
rect 11790 36320 11796 36332
rect 11848 36320 11854 36372
rect 13446 36320 13452 36372
rect 13504 36360 13510 36372
rect 14642 36360 14648 36372
rect 13504 36332 14648 36360
rect 13504 36320 13510 36332
rect 14642 36320 14648 36332
rect 14700 36320 14706 36372
rect 15470 36320 15476 36372
rect 15528 36360 15534 36372
rect 15565 36363 15623 36369
rect 15565 36360 15577 36363
rect 15528 36332 15577 36360
rect 15528 36320 15534 36332
rect 15565 36329 15577 36332
rect 15611 36329 15623 36363
rect 15565 36323 15623 36329
rect 17402 36320 17408 36372
rect 17460 36360 17466 36372
rect 18506 36360 18512 36372
rect 17460 36332 18512 36360
rect 17460 36320 17466 36332
rect 18506 36320 18512 36332
rect 18564 36320 18570 36372
rect 19334 36320 19340 36372
rect 19392 36360 19398 36372
rect 21177 36363 21235 36369
rect 21177 36360 21189 36363
rect 19392 36332 21189 36360
rect 19392 36320 19398 36332
rect 21177 36329 21189 36332
rect 21223 36329 21235 36363
rect 23750 36360 23756 36372
rect 21177 36323 21235 36329
rect 22066 36332 23756 36360
rect 12161 36295 12219 36301
rect 12161 36292 12173 36295
rect 2746 36264 12173 36292
rect 2746 36224 2774 36264
rect 12161 36261 12173 36264
rect 12207 36261 12219 36295
rect 12161 36255 12219 36261
rect 17218 36252 17224 36304
rect 17276 36292 17282 36304
rect 18141 36295 18199 36301
rect 18141 36292 18153 36295
rect 17276 36264 18153 36292
rect 17276 36252 17282 36264
rect 18141 36261 18153 36264
rect 18187 36261 18199 36295
rect 18141 36255 18199 36261
rect 20714 36252 20720 36304
rect 20772 36292 20778 36304
rect 22066 36292 22094 36332
rect 23750 36320 23756 36332
rect 23808 36320 23814 36372
rect 23842 36320 23848 36372
rect 23900 36360 23906 36372
rect 24029 36363 24087 36369
rect 24029 36360 24041 36363
rect 23900 36332 24041 36360
rect 23900 36320 23906 36332
rect 24029 36329 24041 36332
rect 24075 36329 24087 36363
rect 24029 36323 24087 36329
rect 24670 36320 24676 36372
rect 24728 36360 24734 36372
rect 26329 36363 26387 36369
rect 26329 36360 26341 36363
rect 24728 36332 26341 36360
rect 24728 36320 24734 36332
rect 26329 36329 26341 36332
rect 26375 36329 26387 36363
rect 26329 36323 26387 36329
rect 27706 36320 27712 36372
rect 27764 36360 27770 36372
rect 32306 36360 32312 36372
rect 27764 36332 32312 36360
rect 27764 36320 27770 36332
rect 32306 36320 32312 36332
rect 32364 36320 32370 36372
rect 33502 36320 33508 36372
rect 33560 36360 33566 36372
rect 36725 36363 36783 36369
rect 36725 36360 36737 36363
rect 33560 36332 36737 36360
rect 33560 36320 33566 36332
rect 36725 36329 36737 36332
rect 36771 36360 36783 36363
rect 38562 36360 38568 36372
rect 36771 36332 38568 36360
rect 36771 36329 36783 36332
rect 36725 36323 36783 36329
rect 38562 36320 38568 36332
rect 38620 36320 38626 36372
rect 49234 36320 49240 36372
rect 49292 36320 49298 36372
rect 20772 36264 22094 36292
rect 20772 36252 20778 36264
rect 28810 36252 28816 36304
rect 28868 36252 28874 36304
rect 29178 36252 29184 36304
rect 29236 36252 29242 36304
rect 31757 36295 31815 36301
rect 31757 36261 31769 36295
rect 31803 36292 31815 36295
rect 31846 36292 31852 36304
rect 31803 36264 31852 36292
rect 31803 36261 31815 36264
rect 31757 36255 31815 36261
rect 31846 36252 31852 36264
rect 31904 36292 31910 36304
rect 32858 36292 32864 36304
rect 31904 36264 32864 36292
rect 31904 36252 31910 36264
rect 32858 36252 32864 36264
rect 32916 36252 32922 36304
rect 1780 36196 2774 36224
rect 1780 36165 1808 36196
rect 9582 36184 9588 36236
rect 9640 36224 9646 36236
rect 9677 36227 9735 36233
rect 9677 36224 9689 36227
rect 9640 36196 9689 36224
rect 9640 36184 9646 36196
rect 9677 36193 9689 36196
rect 9723 36193 9735 36227
rect 9677 36187 9735 36193
rect 12434 36184 12440 36236
rect 12492 36224 12498 36236
rect 13446 36224 13452 36236
rect 12492 36196 13452 36224
rect 12492 36184 12498 36196
rect 13446 36184 13452 36196
rect 13504 36184 13510 36236
rect 13633 36227 13691 36233
rect 13633 36193 13645 36227
rect 13679 36224 13691 36227
rect 14366 36224 14372 36236
rect 13679 36196 14372 36224
rect 13679 36193 13691 36196
rect 13633 36187 13691 36193
rect 14366 36184 14372 36196
rect 14424 36184 14430 36236
rect 15102 36184 15108 36236
rect 15160 36184 15166 36236
rect 16114 36184 16120 36236
rect 16172 36184 16178 36236
rect 16850 36184 16856 36236
rect 16908 36184 16914 36236
rect 16942 36184 16948 36236
rect 17000 36184 17006 36236
rect 18785 36227 18843 36233
rect 18785 36193 18797 36227
rect 18831 36224 18843 36227
rect 18874 36224 18880 36236
rect 18831 36196 18880 36224
rect 18831 36193 18843 36196
rect 18785 36187 18843 36193
rect 18874 36184 18880 36196
rect 18932 36184 18938 36236
rect 19429 36227 19487 36233
rect 19429 36193 19441 36227
rect 19475 36224 19487 36227
rect 20438 36224 20444 36236
rect 19475 36196 20444 36224
rect 19475 36193 19487 36196
rect 19429 36187 19487 36193
rect 20438 36184 20444 36196
rect 20496 36224 20502 36236
rect 22002 36224 22008 36236
rect 20496 36196 22008 36224
rect 20496 36184 20502 36196
rect 22002 36184 22008 36196
rect 22060 36224 22066 36236
rect 22281 36227 22339 36233
rect 22281 36224 22293 36227
rect 22060 36196 22293 36224
rect 22060 36184 22066 36196
rect 22281 36193 22293 36196
rect 22327 36193 22339 36227
rect 22281 36187 22339 36193
rect 24578 36184 24584 36236
rect 24636 36224 24642 36236
rect 27430 36224 27436 36236
rect 24636 36196 27436 36224
rect 24636 36184 24642 36196
rect 27430 36184 27436 36196
rect 27488 36184 27494 36236
rect 27709 36227 27767 36233
rect 27709 36193 27721 36227
rect 27755 36224 27767 36227
rect 28350 36224 28356 36236
rect 27755 36196 28356 36224
rect 27755 36193 27767 36196
rect 27709 36187 27767 36193
rect 28350 36184 28356 36196
rect 28408 36224 28414 36236
rect 28828 36224 28856 36252
rect 28408 36196 28856 36224
rect 28408 36184 28414 36196
rect 29914 36184 29920 36236
rect 29972 36224 29978 36236
rect 30009 36227 30067 36233
rect 30009 36224 30021 36227
rect 29972 36196 30021 36224
rect 29972 36184 29978 36196
rect 30009 36193 30021 36196
rect 30055 36193 30067 36227
rect 30009 36187 30067 36193
rect 30282 36184 30288 36236
rect 30340 36224 30346 36236
rect 32769 36227 32827 36233
rect 32769 36224 32781 36227
rect 30340 36196 32781 36224
rect 30340 36184 30346 36196
rect 32769 36193 32781 36196
rect 32815 36193 32827 36227
rect 37185 36227 37243 36233
rect 37185 36224 37197 36227
rect 32769 36187 32827 36193
rect 34992 36196 37197 36224
rect 1765 36159 1823 36165
rect 1765 36125 1777 36159
rect 1811 36125 1823 36159
rect 1765 36119 1823 36125
rect 9490 36116 9496 36168
rect 9548 36116 9554 36168
rect 11974 36116 11980 36168
rect 12032 36116 12038 36168
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36156 13415 36159
rect 15010 36156 15016 36168
rect 13403 36128 15016 36156
rect 13403 36125 13415 36128
rect 13357 36119 13415 36125
rect 15010 36116 15016 36128
rect 15068 36116 15074 36168
rect 16758 36116 16764 36168
rect 16816 36156 16822 36168
rect 17589 36159 17647 36165
rect 17589 36156 17601 36159
rect 16816 36128 17601 36156
rect 16816 36116 16822 36128
rect 17589 36125 17601 36128
rect 17635 36156 17647 36159
rect 18601 36159 18659 36165
rect 18601 36156 18613 36159
rect 17635 36128 18613 36156
rect 17635 36125 17647 36128
rect 17589 36119 17647 36125
rect 18601 36125 18613 36128
rect 18647 36156 18659 36159
rect 19058 36156 19064 36168
rect 18647 36128 19064 36156
rect 18647 36125 18659 36128
rect 18601 36119 18659 36125
rect 19058 36116 19064 36128
rect 19116 36116 19122 36168
rect 20806 36116 20812 36168
rect 20864 36116 20870 36168
rect 32306 36116 32312 36168
rect 32364 36156 32370 36168
rect 33413 36159 33471 36165
rect 33413 36156 33425 36159
rect 32364 36128 33425 36156
rect 32364 36116 32370 36128
rect 33413 36125 33425 36128
rect 33459 36156 33471 36159
rect 34882 36156 34888 36168
rect 33459 36128 34888 36156
rect 33459 36125 33471 36128
rect 33413 36119 33471 36125
rect 34882 36116 34888 36128
rect 34940 36116 34946 36168
rect 34992 36165 35020 36196
rect 37185 36193 37197 36196
rect 37231 36193 37243 36227
rect 37185 36187 37243 36193
rect 37461 36227 37519 36233
rect 37461 36193 37473 36227
rect 37507 36224 37519 36227
rect 38654 36224 38660 36236
rect 37507 36196 38660 36224
rect 37507 36193 37519 36196
rect 37461 36187 37519 36193
rect 38654 36184 38660 36196
rect 38712 36184 38718 36236
rect 34977 36159 35035 36165
rect 34977 36125 34989 36159
rect 35023 36125 35035 36159
rect 34977 36119 35035 36125
rect 2774 36048 2780 36100
rect 2832 36048 2838 36100
rect 8389 36091 8447 36097
rect 8389 36057 8401 36091
rect 8435 36088 8447 36091
rect 11054 36088 11060 36100
rect 8435 36060 11060 36088
rect 8435 36057 8447 36060
rect 8389 36051 8447 36057
rect 11054 36048 11060 36060
rect 11112 36048 11118 36100
rect 14642 36048 14648 36100
rect 14700 36088 14706 36100
rect 14921 36091 14979 36097
rect 14921 36088 14933 36091
rect 14700 36060 14933 36088
rect 14700 36048 14706 36060
rect 14921 36057 14933 36060
rect 14967 36057 14979 36091
rect 14921 36051 14979 36057
rect 15470 36048 15476 36100
rect 15528 36088 15534 36100
rect 15933 36091 15991 36097
rect 15933 36088 15945 36091
rect 15528 36060 15945 36088
rect 15528 36048 15534 36060
rect 15933 36057 15945 36060
rect 15979 36057 15991 36091
rect 15933 36051 15991 36057
rect 16025 36091 16083 36097
rect 16025 36057 16037 36091
rect 16071 36088 16083 36091
rect 16298 36088 16304 36100
rect 16071 36060 16304 36088
rect 16071 36057 16083 36060
rect 16025 36051 16083 36057
rect 16298 36048 16304 36060
rect 16356 36048 16362 36100
rect 18509 36091 18567 36097
rect 18509 36057 18521 36091
rect 18555 36088 18567 36091
rect 19150 36088 19156 36100
rect 18555 36060 19156 36088
rect 18555 36057 18567 36060
rect 18509 36051 18567 36057
rect 19150 36048 19156 36060
rect 19208 36048 19214 36100
rect 19702 36048 19708 36100
rect 19760 36048 19766 36100
rect 22557 36091 22615 36097
rect 22557 36057 22569 36091
rect 22603 36057 22615 36091
rect 23842 36088 23848 36100
rect 23782 36060 23848 36088
rect 22557 36051 22615 36057
rect 4798 35980 4804 36032
rect 4856 36020 4862 36032
rect 9585 36023 9643 36029
rect 9585 36020 9597 36023
rect 4856 35992 9597 36020
rect 4856 35980 4862 35992
rect 9585 35989 9597 35992
rect 9631 35989 9643 36023
rect 9585 35983 9643 35989
rect 12989 36023 13047 36029
rect 12989 35989 13001 36023
rect 13035 36020 13047 36023
rect 14182 36020 14188 36032
rect 13035 35992 14188 36020
rect 13035 35989 13047 35992
rect 12989 35983 13047 35989
rect 14182 35980 14188 35992
rect 14240 35980 14246 36032
rect 14550 35980 14556 36032
rect 14608 35980 14614 36032
rect 15013 36023 15071 36029
rect 15013 35989 15025 36023
rect 15059 36020 15071 36023
rect 15102 36020 15108 36032
rect 15059 35992 15108 36020
rect 15059 35989 15071 35992
rect 15013 35983 15071 35989
rect 15102 35980 15108 35992
rect 15160 35980 15166 36032
rect 16390 35980 16396 36032
rect 16448 35980 16454 36032
rect 16761 36023 16819 36029
rect 16761 35989 16773 36023
rect 16807 36020 16819 36023
rect 17034 36020 17040 36032
rect 16807 35992 17040 36020
rect 16807 35989 16819 35992
rect 16761 35983 16819 35989
rect 17034 35980 17040 35992
rect 17092 35980 17098 36032
rect 22572 36020 22600 36051
rect 23842 36048 23848 36060
rect 23900 36048 23906 36100
rect 24486 36048 24492 36100
rect 24544 36088 24550 36100
rect 24857 36091 24915 36097
rect 24857 36088 24869 36091
rect 24544 36060 24869 36088
rect 24544 36048 24550 36060
rect 24857 36057 24869 36060
rect 24903 36088 24915 36091
rect 25130 36088 25136 36100
rect 24903 36060 25136 36088
rect 24903 36057 24915 36060
rect 24857 36051 24915 36057
rect 25130 36048 25136 36060
rect 25188 36048 25194 36100
rect 25498 36048 25504 36100
rect 25556 36048 25562 36100
rect 27706 36048 27712 36100
rect 27764 36088 27770 36100
rect 28166 36088 28172 36100
rect 27764 36060 28172 36088
rect 27764 36048 27770 36060
rect 28166 36048 28172 36060
rect 28224 36048 28230 36100
rect 30285 36091 30343 36097
rect 30285 36057 30297 36091
rect 30331 36057 30343 36091
rect 30285 36051 30343 36057
rect 25866 36020 25872 36032
rect 22572 35992 25872 36020
rect 25866 35980 25872 35992
rect 25924 35980 25930 36032
rect 27890 35980 27896 36032
rect 27948 36020 27954 36032
rect 28534 36020 28540 36032
rect 27948 35992 28540 36020
rect 27948 35980 27954 35992
rect 28534 35980 28540 35992
rect 28592 35980 28598 36032
rect 30300 36020 30328 36051
rect 31294 36048 31300 36100
rect 31352 36048 31358 36100
rect 32585 36091 32643 36097
rect 32585 36088 32597 36091
rect 31726 36060 32597 36088
rect 31018 36020 31024 36032
rect 30300 35992 31024 36020
rect 31018 35980 31024 35992
rect 31076 35980 31082 36032
rect 31202 35980 31208 36032
rect 31260 36020 31266 36032
rect 31726 36020 31754 36060
rect 32585 36057 32597 36060
rect 32631 36057 32643 36091
rect 32585 36051 32643 36057
rect 32674 36048 32680 36100
rect 32732 36048 32738 36100
rect 34146 36048 34152 36100
rect 34204 36088 34210 36100
rect 34992 36088 35020 36119
rect 36354 36116 36360 36168
rect 36412 36156 36418 36168
rect 37090 36156 37096 36168
rect 36412 36128 37096 36156
rect 36412 36116 36418 36128
rect 37090 36116 37096 36128
rect 37148 36116 37154 36168
rect 48314 36116 48320 36168
rect 48372 36156 48378 36168
rect 49053 36159 49111 36165
rect 49053 36156 49065 36159
rect 48372 36128 49065 36156
rect 48372 36116 48378 36128
rect 49053 36125 49065 36128
rect 49099 36125 49111 36159
rect 49053 36119 49111 36125
rect 34204 36060 35020 36088
rect 35253 36091 35311 36097
rect 34204 36048 34210 36060
rect 35253 36057 35265 36091
rect 35299 36088 35311 36091
rect 35342 36088 35348 36100
rect 35299 36060 35348 36088
rect 35299 36057 35311 36060
rect 35253 36051 35311 36057
rect 35342 36048 35348 36060
rect 35400 36048 35406 36100
rect 37366 36088 37372 36100
rect 37016 36060 37372 36088
rect 31260 35992 31754 36020
rect 32217 36023 32275 36029
rect 31260 35980 31266 35992
rect 32217 35989 32229 36023
rect 32263 36020 32275 36023
rect 37016 36020 37044 36060
rect 37366 36048 37372 36060
rect 37424 36048 37430 36100
rect 37458 36048 37464 36100
rect 37516 36088 37522 36100
rect 37516 36060 37950 36088
rect 37516 36048 37522 36060
rect 32263 35992 37044 36020
rect 32263 35989 32275 35992
rect 32217 35983 32275 35989
rect 37090 35980 37096 36032
rect 37148 36020 37154 36032
rect 38838 36020 38844 36032
rect 37148 35992 38844 36020
rect 37148 35980 37154 35992
rect 38838 35980 38844 35992
rect 38896 36020 38902 36032
rect 38933 36023 38991 36029
rect 38933 36020 38945 36023
rect 38896 35992 38945 36020
rect 38896 35980 38902 35992
rect 38933 35989 38945 35992
rect 38979 35989 38991 36023
rect 38933 35983 38991 35989
rect 1104 35930 49864 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 27950 35930
rect 28002 35878 28014 35930
rect 28066 35878 28078 35930
rect 28130 35878 28142 35930
rect 28194 35878 28206 35930
rect 28258 35878 37950 35930
rect 38002 35878 38014 35930
rect 38066 35878 38078 35930
rect 38130 35878 38142 35930
rect 38194 35878 38206 35930
rect 38258 35878 47950 35930
rect 48002 35878 48014 35930
rect 48066 35878 48078 35930
rect 48130 35878 48142 35930
rect 48194 35878 48206 35930
rect 48258 35878 49864 35930
rect 1104 35856 49864 35878
rect 3418 35776 3424 35828
rect 3476 35816 3482 35828
rect 9401 35819 9459 35825
rect 9401 35816 9413 35819
rect 3476 35788 9413 35816
rect 3476 35776 3482 35788
rect 9401 35785 9413 35788
rect 9447 35785 9459 35819
rect 9401 35779 9459 35785
rect 12618 35776 12624 35828
rect 12676 35816 12682 35828
rect 12676 35788 14780 35816
rect 12676 35776 12682 35788
rect 9306 35708 9312 35760
rect 9364 35708 9370 35760
rect 14642 35748 14648 35760
rect 14582 35720 14648 35748
rect 14642 35708 14648 35720
rect 14700 35708 14706 35760
rect 14752 35748 14780 35788
rect 14826 35776 14832 35828
rect 14884 35776 14890 35828
rect 15194 35776 15200 35828
rect 15252 35816 15258 35828
rect 15933 35819 15991 35825
rect 15933 35816 15945 35819
rect 15252 35788 15945 35816
rect 15252 35776 15258 35788
rect 15933 35785 15945 35788
rect 15979 35785 15991 35819
rect 15933 35779 15991 35785
rect 16022 35776 16028 35828
rect 16080 35816 16086 35828
rect 17865 35819 17923 35825
rect 17865 35816 17877 35819
rect 16080 35788 17877 35816
rect 16080 35776 16086 35788
rect 17865 35785 17877 35788
rect 17911 35785 17923 35819
rect 17865 35779 17923 35785
rect 17954 35776 17960 35828
rect 18012 35816 18018 35828
rect 19150 35816 19156 35828
rect 18012 35788 19156 35816
rect 18012 35776 18018 35788
rect 19150 35776 19156 35788
rect 19208 35816 19214 35828
rect 20714 35816 20720 35828
rect 19208 35788 20720 35816
rect 19208 35776 19214 35788
rect 20714 35776 20720 35788
rect 20772 35776 20778 35828
rect 23308 35788 31754 35816
rect 15654 35748 15660 35760
rect 14752 35720 15660 35748
rect 15654 35708 15660 35720
rect 15712 35708 15718 35760
rect 15746 35708 15752 35760
rect 15804 35748 15810 35760
rect 15841 35751 15899 35757
rect 15841 35748 15853 35751
rect 15804 35720 15853 35748
rect 15804 35708 15810 35720
rect 15841 35717 15853 35720
rect 15887 35717 15899 35751
rect 15841 35711 15899 35717
rect 17126 35708 17132 35760
rect 17184 35748 17190 35760
rect 17184 35720 18368 35748
rect 17184 35708 17190 35720
rect 17954 35680 17960 35692
rect 15396 35652 17960 35680
rect 9582 35572 9588 35624
rect 9640 35572 9646 35624
rect 13081 35615 13139 35621
rect 13081 35581 13093 35615
rect 13127 35581 13139 35615
rect 13081 35575 13139 35581
rect 13357 35615 13415 35621
rect 13357 35581 13369 35615
rect 13403 35612 13415 35615
rect 13722 35612 13728 35624
rect 13403 35584 13728 35612
rect 13403 35581 13415 35584
rect 13357 35575 13415 35581
rect 8941 35479 8999 35485
rect 8941 35445 8953 35479
rect 8987 35476 8999 35479
rect 10778 35476 10784 35488
rect 8987 35448 10784 35476
rect 8987 35445 8999 35448
rect 8941 35439 8999 35445
rect 10778 35436 10784 35448
rect 10836 35436 10842 35488
rect 13096 35476 13124 35575
rect 13722 35572 13728 35584
rect 13780 35612 13786 35624
rect 15286 35612 15292 35624
rect 13780 35584 15292 35612
rect 13780 35572 13786 35584
rect 15286 35572 15292 35584
rect 15344 35572 15350 35624
rect 14090 35476 14096 35488
rect 13096 35448 14096 35476
rect 14090 35436 14096 35448
rect 14148 35436 14154 35488
rect 14458 35436 14464 35488
rect 14516 35476 14522 35488
rect 15396 35476 15424 35652
rect 17954 35640 17960 35652
rect 18012 35640 18018 35692
rect 18230 35640 18236 35692
rect 18288 35640 18294 35692
rect 18340 35680 18368 35720
rect 19334 35708 19340 35760
rect 19392 35748 19398 35760
rect 19797 35751 19855 35757
rect 19797 35748 19809 35751
rect 19392 35720 19809 35748
rect 19392 35708 19398 35720
rect 19797 35717 19809 35720
rect 19843 35717 19855 35751
rect 19797 35711 19855 35717
rect 20806 35708 20812 35760
rect 20864 35708 20870 35760
rect 22094 35708 22100 35760
rect 22152 35748 22158 35760
rect 23201 35751 23259 35757
rect 23201 35748 23213 35751
rect 22152 35720 23213 35748
rect 22152 35708 22158 35720
rect 23201 35717 23213 35720
rect 23247 35717 23259 35751
rect 23201 35711 23259 35717
rect 18340 35652 18460 35680
rect 16117 35615 16175 35621
rect 16117 35581 16129 35615
rect 16163 35612 16175 35615
rect 17770 35612 17776 35624
rect 16163 35584 17776 35612
rect 16163 35581 16175 35584
rect 16117 35575 16175 35581
rect 17770 35572 17776 35584
rect 17828 35572 17834 35624
rect 18432 35621 18460 35652
rect 22186 35640 22192 35692
rect 22244 35640 22250 35692
rect 23308 35680 23336 35788
rect 23842 35708 23848 35760
rect 23900 35748 23906 35760
rect 28442 35748 28448 35760
rect 23900 35720 24886 35748
rect 28276 35720 28448 35748
rect 23900 35708 23906 35720
rect 28276 35689 28304 35720
rect 28442 35708 28448 35720
rect 28500 35708 28506 35760
rect 28626 35708 28632 35760
rect 28684 35748 28690 35760
rect 28684 35720 29026 35748
rect 28684 35708 28690 35720
rect 30374 35708 30380 35760
rect 30432 35748 30438 35760
rect 31570 35748 31576 35760
rect 30432 35720 31576 35748
rect 30432 35708 30438 35720
rect 31570 35708 31576 35720
rect 31628 35708 31634 35760
rect 31726 35748 31754 35788
rect 32030 35776 32036 35828
rect 32088 35816 32094 35828
rect 33870 35816 33876 35828
rect 32088 35788 33876 35816
rect 32088 35776 32094 35788
rect 33870 35776 33876 35788
rect 33928 35776 33934 35828
rect 34054 35776 34060 35828
rect 34112 35816 34118 35828
rect 35897 35819 35955 35825
rect 34112 35788 35756 35816
rect 34112 35776 34118 35788
rect 32214 35748 32220 35760
rect 31726 35720 32220 35748
rect 32214 35708 32220 35720
rect 32272 35708 32278 35760
rect 32306 35708 32312 35760
rect 32364 35708 32370 35760
rect 34698 35748 34704 35760
rect 34164 35720 34704 35748
rect 22756 35652 23336 35680
rect 28261 35683 28319 35689
rect 18325 35615 18383 35621
rect 18325 35581 18337 35615
rect 18371 35581 18383 35615
rect 18325 35575 18383 35581
rect 18417 35615 18475 35621
rect 18417 35581 18429 35615
rect 18463 35581 18475 35615
rect 18417 35575 18475 35581
rect 17405 35547 17463 35553
rect 17405 35513 17417 35547
rect 17451 35544 17463 35547
rect 18340 35544 18368 35575
rect 19058 35572 19064 35624
rect 19116 35612 19122 35624
rect 19521 35615 19579 35621
rect 19521 35612 19533 35615
rect 19116 35584 19533 35612
rect 19116 35572 19122 35584
rect 19521 35581 19533 35584
rect 19567 35581 19579 35615
rect 19521 35575 19579 35581
rect 22756 35544 22784 35652
rect 28261 35649 28273 35683
rect 28307 35649 28319 35683
rect 28261 35643 28319 35649
rect 30837 35683 30895 35689
rect 30837 35649 30849 35683
rect 30883 35680 30895 35683
rect 34164 35680 34192 35720
rect 34698 35708 34704 35720
rect 34756 35708 34762 35760
rect 30883 35652 34192 35680
rect 35728 35680 35756 35788
rect 35897 35785 35909 35819
rect 35943 35816 35955 35819
rect 35986 35816 35992 35828
rect 35943 35788 35992 35816
rect 35943 35785 35955 35788
rect 35897 35779 35955 35785
rect 35986 35776 35992 35788
rect 36044 35816 36050 35828
rect 36906 35816 36912 35828
rect 36044 35788 36912 35816
rect 36044 35776 36050 35788
rect 36906 35776 36912 35788
rect 36964 35776 36970 35828
rect 38197 35683 38255 35689
rect 38197 35680 38209 35683
rect 30883 35649 30895 35652
rect 30837 35643 30895 35649
rect 23293 35615 23351 35621
rect 23293 35581 23305 35615
rect 23339 35581 23351 35615
rect 23293 35575 23351 35581
rect 17451 35516 18368 35544
rect 17451 35513 17463 35516
rect 17405 35507 17463 35513
rect 14516 35448 15424 35476
rect 15473 35479 15531 35485
rect 14516 35436 14522 35448
rect 15473 35445 15485 35479
rect 15519 35476 15531 35479
rect 16114 35476 16120 35488
rect 15519 35448 16120 35476
rect 15519 35445 15531 35448
rect 15473 35439 15531 35445
rect 16114 35436 16120 35448
rect 16172 35436 16178 35488
rect 18340 35476 18368 35516
rect 20824 35516 22784 35544
rect 22833 35547 22891 35553
rect 20824 35476 20852 35516
rect 22833 35513 22845 35547
rect 22879 35513 22891 35547
rect 22833 35507 22891 35513
rect 18340 35448 20852 35476
rect 21266 35436 21272 35488
rect 21324 35436 21330 35488
rect 21450 35436 21456 35488
rect 21508 35476 21514 35488
rect 22848 35476 22876 35507
rect 21508 35448 22876 35476
rect 23308 35476 23336 35575
rect 23382 35572 23388 35624
rect 23440 35572 23446 35624
rect 24121 35615 24179 35621
rect 24121 35581 24133 35615
rect 24167 35612 24179 35615
rect 24397 35615 24455 35621
rect 24167 35584 24256 35612
rect 24167 35581 24179 35584
rect 24121 35575 24179 35581
rect 23382 35476 23388 35488
rect 23308 35448 23388 35476
rect 21508 35436 21514 35448
rect 23382 35436 23388 35448
rect 23440 35436 23446 35488
rect 24228 35476 24256 35584
rect 24397 35581 24409 35615
rect 24443 35612 24455 35615
rect 24946 35612 24952 35624
rect 24443 35584 24952 35612
rect 24443 35581 24455 35584
rect 24397 35575 24455 35581
rect 24946 35572 24952 35584
rect 25004 35572 25010 35624
rect 25866 35572 25872 35624
rect 25924 35572 25930 35624
rect 28537 35615 28595 35621
rect 28537 35581 28549 35615
rect 28583 35612 28595 35615
rect 29086 35612 29092 35624
rect 28583 35584 29092 35612
rect 28583 35581 28595 35584
rect 28537 35575 28595 35581
rect 29086 35572 29092 35584
rect 29144 35572 29150 35624
rect 30190 35572 30196 35624
rect 30248 35612 30254 35624
rect 30929 35615 30987 35621
rect 30929 35612 30941 35615
rect 30248 35584 30941 35612
rect 30248 35572 30254 35584
rect 30929 35581 30941 35584
rect 30975 35581 30987 35615
rect 30929 35575 30987 35581
rect 31018 35572 31024 35624
rect 31076 35612 31082 35624
rect 31478 35612 31484 35624
rect 31076 35584 31484 35612
rect 31076 35572 31082 35584
rect 31478 35572 31484 35584
rect 31536 35572 31542 35624
rect 32490 35572 32496 35624
rect 32548 35612 32554 35624
rect 33045 35615 33103 35621
rect 33045 35612 33057 35615
rect 32548 35584 33057 35612
rect 32548 35572 32554 35584
rect 33045 35581 33057 35584
rect 33091 35581 33103 35615
rect 33045 35575 33103 35581
rect 33686 35572 33692 35624
rect 33744 35612 33750 35624
rect 33744 35584 34100 35612
rect 33744 35572 33750 35584
rect 30009 35547 30067 35553
rect 30009 35513 30021 35547
rect 30055 35544 30067 35547
rect 30282 35544 30288 35556
rect 30055 35516 30288 35544
rect 30055 35513 30067 35516
rect 30009 35507 30067 35513
rect 30282 35504 30288 35516
rect 30340 35504 30346 35556
rect 31110 35504 31116 35556
rect 31168 35544 31174 35556
rect 33962 35544 33968 35556
rect 31168 35516 33968 35544
rect 31168 35504 31174 35516
rect 33962 35504 33968 35516
rect 34020 35504 34026 35556
rect 34072 35544 34100 35584
rect 34146 35572 34152 35624
rect 34204 35572 34210 35624
rect 34425 35615 34483 35621
rect 34425 35612 34437 35615
rect 34256 35584 34437 35612
rect 34256 35544 34284 35584
rect 34425 35581 34437 35584
rect 34471 35612 34483 35615
rect 35158 35612 35164 35624
rect 34471 35584 35164 35612
rect 34471 35581 34483 35584
rect 34425 35575 34483 35581
rect 35158 35572 35164 35584
rect 35216 35572 35222 35624
rect 35544 35612 35572 35666
rect 35728 35652 38209 35680
rect 38197 35649 38209 35652
rect 38243 35649 38255 35683
rect 38197 35643 38255 35649
rect 36354 35612 36360 35624
rect 35544 35584 36360 35612
rect 34072 35516 34284 35544
rect 24578 35476 24584 35488
rect 24228 35448 24584 35476
rect 24578 35436 24584 35448
rect 24636 35436 24642 35488
rect 25038 35436 25044 35488
rect 25096 35476 25102 35488
rect 27246 35476 27252 35488
rect 25096 35448 27252 35476
rect 25096 35436 25102 35448
rect 27246 35436 27252 35448
rect 27304 35436 27310 35488
rect 30469 35479 30527 35485
rect 30469 35445 30481 35479
rect 30515 35476 30527 35479
rect 33778 35476 33784 35488
rect 30515 35448 33784 35476
rect 30515 35445 30527 35448
rect 30469 35439 30527 35445
rect 33778 35436 33784 35448
rect 33836 35436 33842 35488
rect 34422 35436 34428 35488
rect 34480 35476 34486 35488
rect 35544 35476 35572 35584
rect 36354 35572 36360 35584
rect 36412 35572 36418 35624
rect 34480 35448 35572 35476
rect 38013 35479 38071 35485
rect 34480 35436 34486 35448
rect 38013 35445 38025 35479
rect 38059 35476 38071 35479
rect 39942 35476 39948 35488
rect 38059 35448 39948 35476
rect 38059 35445 38071 35448
rect 38013 35439 38071 35445
rect 39942 35436 39948 35448
rect 40000 35436 40006 35488
rect 1104 35386 49864 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 32950 35386
rect 33002 35334 33014 35386
rect 33066 35334 33078 35386
rect 33130 35334 33142 35386
rect 33194 35334 33206 35386
rect 33258 35334 42950 35386
rect 43002 35334 43014 35386
rect 43066 35334 43078 35386
rect 43130 35334 43142 35386
rect 43194 35334 43206 35386
rect 43258 35334 49864 35386
rect 1104 35312 49864 35334
rect 16669 35275 16727 35281
rect 16669 35272 16681 35275
rect 14016 35244 16681 35272
rect 1302 35096 1308 35148
rect 1360 35136 1366 35148
rect 2041 35139 2099 35145
rect 2041 35136 2053 35139
rect 1360 35108 2053 35136
rect 1360 35096 1366 35108
rect 2041 35105 2053 35108
rect 2087 35105 2099 35139
rect 11793 35139 11851 35145
rect 11793 35136 11805 35139
rect 2041 35099 2099 35105
rect 2746 35108 11805 35136
rect 1765 35071 1823 35077
rect 1765 35037 1777 35071
rect 1811 35068 1823 35071
rect 2746 35068 2774 35108
rect 11793 35105 11805 35108
rect 11839 35105 11851 35139
rect 11793 35099 11851 35105
rect 12618 35096 12624 35148
rect 12676 35136 12682 35148
rect 13538 35136 13544 35148
rect 12676 35108 13544 35136
rect 12676 35096 12682 35108
rect 13538 35096 13544 35108
rect 13596 35096 13602 35148
rect 1811 35040 2774 35068
rect 1811 35037 1823 35040
rect 1765 35031 1823 35037
rect 10870 35028 10876 35080
rect 10928 35028 10934 35080
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35068 13415 35071
rect 14016 35068 14044 35244
rect 16669 35241 16681 35244
rect 16715 35241 16727 35275
rect 16669 35235 16727 35241
rect 18782 35232 18788 35284
rect 18840 35272 18846 35284
rect 21450 35272 21456 35284
rect 18840 35244 21456 35272
rect 18840 35232 18846 35244
rect 21450 35232 21456 35244
rect 21508 35232 21514 35284
rect 22370 35232 22376 35284
rect 22428 35232 22434 35284
rect 23293 35275 23351 35281
rect 23293 35241 23305 35275
rect 23339 35272 23351 35275
rect 23658 35272 23664 35284
rect 23339 35244 23664 35272
rect 23339 35241 23351 35244
rect 23293 35235 23351 35241
rect 23658 35232 23664 35244
rect 23716 35232 23722 35284
rect 24946 35232 24952 35284
rect 25004 35272 25010 35284
rect 26421 35275 26479 35281
rect 26421 35272 26433 35275
rect 25004 35244 26433 35272
rect 25004 35232 25010 35244
rect 26421 35241 26433 35244
rect 26467 35241 26479 35275
rect 26421 35235 26479 35241
rect 29086 35232 29092 35284
rect 29144 35272 29150 35284
rect 30282 35272 30288 35284
rect 29144 35244 30288 35272
rect 29144 35232 29150 35244
rect 30282 35232 30288 35244
rect 30340 35232 30346 35284
rect 30929 35275 30987 35281
rect 30929 35241 30941 35275
rect 30975 35272 30987 35275
rect 31110 35272 31116 35284
rect 30975 35244 31116 35272
rect 30975 35241 30987 35244
rect 30929 35235 30987 35241
rect 31110 35232 31116 35244
rect 31168 35232 31174 35284
rect 33413 35275 33471 35281
rect 31220 35244 32720 35272
rect 15654 35164 15660 35216
rect 15712 35204 15718 35216
rect 16025 35207 16083 35213
rect 16025 35204 16037 35207
rect 15712 35176 16037 35204
rect 15712 35164 15718 35176
rect 16025 35173 16037 35176
rect 16071 35173 16083 35207
rect 16025 35167 16083 35173
rect 16206 35164 16212 35216
rect 16264 35204 16270 35216
rect 27525 35207 27583 35213
rect 16264 35176 18552 35204
rect 16264 35164 16270 35176
rect 14090 35096 14096 35148
rect 14148 35136 14154 35148
rect 14277 35139 14335 35145
rect 14277 35136 14289 35139
rect 14148 35108 14289 35136
rect 14148 35096 14154 35108
rect 14277 35105 14289 35108
rect 14323 35136 14335 35139
rect 15286 35136 15292 35148
rect 14323 35108 15292 35136
rect 14323 35105 14335 35108
rect 14277 35099 14335 35105
rect 15286 35096 15292 35108
rect 15344 35096 15350 35148
rect 16390 35096 16396 35148
rect 16448 35136 16454 35148
rect 17129 35139 17187 35145
rect 17129 35136 17141 35139
rect 16448 35108 17141 35136
rect 16448 35096 16454 35108
rect 17129 35105 17141 35108
rect 17175 35105 17187 35139
rect 17129 35099 17187 35105
rect 17313 35139 17371 35145
rect 17313 35105 17325 35139
rect 17359 35136 17371 35139
rect 17494 35136 17500 35148
rect 17359 35108 17500 35136
rect 17359 35105 17371 35108
rect 17313 35099 17371 35105
rect 13403 35040 14044 35068
rect 13403 35037 13415 35040
rect 13357 35031 13415 35037
rect 15838 35028 15844 35080
rect 15896 35068 15902 35080
rect 17328 35068 17356 35099
rect 17494 35096 17500 35108
rect 17552 35096 17558 35148
rect 18322 35096 18328 35148
rect 18380 35096 18386 35148
rect 18524 35145 18552 35176
rect 23768 35176 24808 35204
rect 23768 35148 23796 35176
rect 18509 35139 18567 35145
rect 18509 35105 18521 35139
rect 18555 35136 18567 35139
rect 19610 35136 19616 35148
rect 18555 35108 19616 35136
rect 18555 35105 18567 35108
rect 18509 35099 18567 35105
rect 19610 35096 19616 35108
rect 19668 35136 19674 35148
rect 19981 35139 20039 35145
rect 19981 35136 19993 35139
rect 19668 35108 19993 35136
rect 19668 35096 19674 35108
rect 19981 35105 19993 35108
rect 20027 35105 20039 35139
rect 19981 35099 20039 35105
rect 20438 35096 20444 35148
rect 20496 35136 20502 35148
rect 20625 35139 20683 35145
rect 20625 35136 20637 35139
rect 20496 35108 20637 35136
rect 20496 35096 20502 35108
rect 20625 35105 20637 35108
rect 20671 35105 20683 35139
rect 20625 35099 20683 35105
rect 20901 35139 20959 35145
rect 20901 35105 20913 35139
rect 20947 35136 20959 35139
rect 21266 35136 21272 35148
rect 20947 35108 21272 35136
rect 20947 35105 20959 35108
rect 20901 35099 20959 35105
rect 21266 35096 21272 35108
rect 21324 35136 21330 35148
rect 22554 35136 22560 35148
rect 21324 35108 22560 35136
rect 21324 35096 21330 35108
rect 22554 35096 22560 35108
rect 22612 35096 22618 35148
rect 23750 35096 23756 35148
rect 23808 35096 23814 35148
rect 23937 35139 23995 35145
rect 23937 35105 23949 35139
rect 23983 35136 23995 35139
rect 24486 35136 24492 35148
rect 23983 35108 24492 35136
rect 23983 35105 23995 35108
rect 23937 35099 23995 35105
rect 24486 35096 24492 35108
rect 24544 35096 24550 35148
rect 24578 35096 24584 35148
rect 24636 35136 24642 35148
rect 24673 35139 24731 35145
rect 24673 35136 24685 35139
rect 24636 35108 24685 35136
rect 24636 35096 24642 35108
rect 24673 35105 24685 35108
rect 24719 35105 24731 35139
rect 24780 35136 24808 35176
rect 27525 35173 27537 35207
rect 27571 35204 27583 35207
rect 29270 35204 29276 35216
rect 27571 35176 29276 35204
rect 27571 35173 27583 35176
rect 27525 35167 27583 35173
rect 29270 35164 29276 35176
rect 29328 35164 29334 35216
rect 29733 35207 29791 35213
rect 29733 35173 29745 35207
rect 29779 35204 29791 35207
rect 31018 35204 31024 35216
rect 29779 35176 31024 35204
rect 29779 35173 29791 35176
rect 29733 35167 29791 35173
rect 31018 35164 31024 35176
rect 31076 35164 31082 35216
rect 24780 35108 27936 35136
rect 24673 35099 24731 35105
rect 15896 35040 17356 35068
rect 15896 35028 15902 35040
rect 17862 35028 17868 35080
rect 17920 35068 17926 35080
rect 18233 35071 18291 35077
rect 18233 35068 18245 35071
rect 17920 35040 18245 35068
rect 17920 35028 17926 35040
rect 18233 35037 18245 35040
rect 18279 35037 18291 35071
rect 18233 35031 18291 35037
rect 19797 35071 19855 35077
rect 19797 35037 19809 35071
rect 19843 35068 19855 35071
rect 20346 35068 20352 35080
rect 19843 35040 20352 35068
rect 19843 35037 19855 35040
rect 19797 35031 19855 35037
rect 20346 35028 20352 35040
rect 20404 35028 20410 35080
rect 27908 35077 27936 35108
rect 27982 35096 27988 35148
rect 28040 35096 28046 35148
rect 28169 35139 28227 35145
rect 28169 35105 28181 35139
rect 28215 35136 28227 35139
rect 28215 35108 28948 35136
rect 28215 35105 28227 35108
rect 28169 35099 28227 35105
rect 27893 35071 27951 35077
rect 27893 35037 27905 35071
rect 27939 35037 27951 35071
rect 27893 35031 27951 35037
rect 11609 35003 11667 35009
rect 11609 34969 11621 35003
rect 11655 35000 11667 35003
rect 14458 35000 14464 35012
rect 11655 34972 14464 35000
rect 11655 34969 11667 34972
rect 11609 34963 11667 34969
rect 14458 34960 14464 34972
rect 14516 34960 14522 35012
rect 14553 35003 14611 35009
rect 14553 34969 14565 35003
rect 14599 35000 14611 35003
rect 14826 35000 14832 35012
rect 14599 34972 14832 35000
rect 14599 34969 14611 34972
rect 14553 34963 14611 34969
rect 14826 34960 14832 34972
rect 14884 34960 14890 35012
rect 16022 35000 16028 35012
rect 15778 34972 16028 35000
rect 16022 34960 16028 34972
rect 16080 34960 16086 35012
rect 17037 35003 17095 35009
rect 17037 34969 17049 35003
rect 17083 35000 17095 35003
rect 20530 35000 20536 35012
rect 17083 34972 20536 35000
rect 17083 34969 17095 34972
rect 17037 34963 17095 34969
rect 20530 34960 20536 34972
rect 20588 34960 20594 35012
rect 20806 34960 20812 35012
rect 20864 35000 20870 35012
rect 23661 35003 23719 35009
rect 20864 34972 21390 35000
rect 20864 34960 20870 34972
rect 23661 34969 23673 35003
rect 23707 35000 23719 35003
rect 24949 35003 25007 35009
rect 23707 34972 24900 35000
rect 23707 34969 23719 34972
rect 23661 34963 23719 34969
rect 10962 34892 10968 34944
rect 11020 34892 11026 34944
rect 12986 34892 12992 34944
rect 13044 34892 13050 34944
rect 13446 34892 13452 34944
rect 13504 34892 13510 34944
rect 17862 34892 17868 34944
rect 17920 34892 17926 34944
rect 18414 34892 18420 34944
rect 18472 34932 18478 34944
rect 19429 34935 19487 34941
rect 19429 34932 19441 34935
rect 18472 34904 19441 34932
rect 18472 34892 18478 34904
rect 19429 34901 19441 34904
rect 19475 34901 19487 34935
rect 19429 34895 19487 34901
rect 19886 34892 19892 34944
rect 19944 34892 19950 34944
rect 20438 34892 20444 34944
rect 20496 34932 20502 34944
rect 22462 34932 22468 34944
rect 20496 34904 22468 34932
rect 20496 34892 20502 34904
rect 22462 34892 22468 34904
rect 22520 34892 22526 34944
rect 24872 34932 24900 34972
rect 24949 34969 24961 35003
rect 24995 35000 25007 35003
rect 25038 35000 25044 35012
rect 24995 34972 25044 35000
rect 24995 34969 25007 34972
rect 24949 34963 25007 34969
rect 25038 34960 25044 34972
rect 25096 34960 25102 35012
rect 25682 34960 25688 35012
rect 25740 34960 25746 35012
rect 28920 35000 28948 35108
rect 29178 35096 29184 35148
rect 29236 35136 29242 35148
rect 29236 35108 30236 35136
rect 29236 35096 29242 35108
rect 28997 35071 29055 35077
rect 28997 35037 29009 35071
rect 29043 35068 29055 35071
rect 30101 35071 30159 35077
rect 30101 35068 30113 35071
rect 29043 35040 30113 35068
rect 29043 35037 29055 35040
rect 28997 35031 29055 35037
rect 30101 35037 30113 35040
rect 30147 35037 30159 35071
rect 30208 35068 30236 35108
rect 30282 35096 30288 35148
rect 30340 35096 30346 35148
rect 31220 35068 31248 35244
rect 32125 35207 32183 35213
rect 32125 35173 32137 35207
rect 32171 35173 32183 35207
rect 32125 35167 32183 35173
rect 31573 35139 31631 35145
rect 31573 35105 31585 35139
rect 31619 35105 31631 35139
rect 31573 35099 31631 35105
rect 30208 35040 31248 35068
rect 31588 35068 31616 35099
rect 32030 35068 32036 35080
rect 31588 35040 32036 35068
rect 30101 35031 30159 35037
rect 32030 35028 32036 35040
rect 32088 35028 32094 35080
rect 32140 35068 32168 35167
rect 32582 35096 32588 35148
rect 32640 35096 32646 35148
rect 32692 35145 32720 35244
rect 33413 35241 33425 35275
rect 33459 35272 33471 35275
rect 37182 35272 37188 35284
rect 33459 35244 37188 35272
rect 33459 35241 33471 35244
rect 33413 35235 33471 35241
rect 37182 35232 37188 35244
rect 37240 35232 37246 35284
rect 34790 35204 34796 35216
rect 32784 35176 34796 35204
rect 32677 35139 32735 35145
rect 32677 35105 32689 35139
rect 32723 35105 32735 35139
rect 32677 35099 32735 35105
rect 32784 35068 32812 35176
rect 34790 35164 34796 35176
rect 34848 35164 34854 35216
rect 32858 35096 32864 35148
rect 32916 35136 32922 35148
rect 33965 35139 34023 35145
rect 33965 35136 33977 35139
rect 32916 35108 33977 35136
rect 32916 35096 32922 35108
rect 33965 35105 33977 35108
rect 34011 35105 34023 35139
rect 33965 35099 34023 35105
rect 35158 35096 35164 35148
rect 35216 35136 35222 35148
rect 36633 35139 36691 35145
rect 36633 35136 36645 35139
rect 35216 35108 36645 35136
rect 35216 35096 35222 35108
rect 36633 35105 36645 35108
rect 36679 35105 36691 35139
rect 36633 35099 36691 35105
rect 32140 35040 32812 35068
rect 33778 35028 33784 35080
rect 33836 35028 33842 35080
rect 34146 35028 34152 35080
rect 34204 35068 34210 35080
rect 34422 35068 34428 35080
rect 34204 35040 34428 35068
rect 34204 35028 34210 35040
rect 34422 35028 34428 35040
rect 34480 35068 34486 35080
rect 34885 35071 34943 35077
rect 34885 35068 34897 35071
rect 34480 35040 34897 35068
rect 34480 35028 34486 35040
rect 34885 35037 34897 35040
rect 34931 35037 34943 35071
rect 34885 35031 34943 35037
rect 36262 35028 36268 35080
rect 36320 35028 36326 35080
rect 39482 35028 39488 35080
rect 39540 35068 39546 35080
rect 40221 35071 40279 35077
rect 40221 35068 40233 35071
rect 39540 35040 40233 35068
rect 39540 35028 39546 35040
rect 40221 35037 40233 35040
rect 40267 35037 40279 35071
rect 40221 35031 40279 35037
rect 49050 35028 49056 35080
rect 49108 35028 49114 35080
rect 30374 35000 30380 35012
rect 28920 34972 30380 35000
rect 30374 34960 30380 34972
rect 30432 34960 30438 35012
rect 31297 35003 31355 35009
rect 31297 34969 31309 35003
rect 31343 35000 31355 35003
rect 33686 35000 33692 35012
rect 31343 34972 33692 35000
rect 31343 34969 31355 34972
rect 31297 34963 31355 34969
rect 33686 34960 33692 34972
rect 33744 34960 33750 35012
rect 34238 34960 34244 35012
rect 34296 35000 34302 35012
rect 35161 35003 35219 35009
rect 35161 35000 35173 35003
rect 34296 34972 35173 35000
rect 34296 34960 34302 34972
rect 35161 34969 35173 34972
rect 35207 34969 35219 35003
rect 35161 34963 35219 34969
rect 25958 34932 25964 34944
rect 24872 34904 25964 34932
rect 25958 34892 25964 34904
rect 26016 34892 26022 34944
rect 29454 34892 29460 34944
rect 29512 34932 29518 34944
rect 30193 34935 30251 34941
rect 30193 34932 30205 34935
rect 29512 34904 30205 34932
rect 29512 34892 29518 34904
rect 30193 34901 30205 34904
rect 30239 34901 30251 34935
rect 30193 34895 30251 34901
rect 31389 34935 31447 34941
rect 31389 34901 31401 34935
rect 31435 34932 31447 34935
rect 31478 34932 31484 34944
rect 31435 34904 31484 34932
rect 31435 34901 31447 34904
rect 31389 34895 31447 34901
rect 31478 34892 31484 34904
rect 31536 34892 31542 34944
rect 32214 34892 32220 34944
rect 32272 34932 32278 34944
rect 32493 34935 32551 34941
rect 32493 34932 32505 34935
rect 32272 34904 32505 34932
rect 32272 34892 32278 34904
rect 32493 34901 32505 34904
rect 32539 34901 32551 34935
rect 32493 34895 32551 34901
rect 33873 34935 33931 34941
rect 33873 34901 33885 34935
rect 33919 34932 33931 34935
rect 34974 34932 34980 34944
rect 33919 34904 34980 34932
rect 33919 34901 33931 34904
rect 33873 34895 33931 34901
rect 34974 34892 34980 34904
rect 35032 34892 35038 34944
rect 35176 34932 35204 34963
rect 37090 34932 37096 34944
rect 35176 34904 37096 34932
rect 37090 34892 37096 34904
rect 37148 34892 37154 34944
rect 40037 34935 40095 34941
rect 40037 34901 40049 34935
rect 40083 34932 40095 34935
rect 42610 34932 42616 34944
rect 40083 34904 42616 34932
rect 40083 34901 40095 34904
rect 40037 34895 40095 34901
rect 42610 34892 42616 34904
rect 42668 34892 42674 34944
rect 48314 34892 48320 34944
rect 48372 34932 48378 34944
rect 49237 34935 49295 34941
rect 49237 34932 49249 34935
rect 48372 34904 49249 34932
rect 48372 34892 48378 34904
rect 49237 34901 49249 34904
rect 49283 34901 49295 34935
rect 49237 34895 49295 34901
rect 1104 34842 49864 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 27950 34842
rect 28002 34790 28014 34842
rect 28066 34790 28078 34842
rect 28130 34790 28142 34842
rect 28194 34790 28206 34842
rect 28258 34790 37950 34842
rect 38002 34790 38014 34842
rect 38066 34790 38078 34842
rect 38130 34790 38142 34842
rect 38194 34790 38206 34842
rect 38258 34790 47950 34842
rect 48002 34790 48014 34842
rect 48066 34790 48078 34842
rect 48130 34790 48142 34842
rect 48194 34790 48206 34842
rect 48258 34790 49864 34842
rect 1104 34768 49864 34790
rect 13446 34688 13452 34740
rect 13504 34728 13510 34740
rect 14277 34731 14335 34737
rect 14277 34728 14289 34731
rect 13504 34700 14289 34728
rect 13504 34688 13510 34700
rect 14277 34697 14289 34700
rect 14323 34697 14335 34731
rect 14277 34691 14335 34697
rect 14550 34688 14556 34740
rect 14608 34728 14614 34740
rect 14645 34731 14703 34737
rect 14645 34728 14657 34731
rect 14608 34700 14657 34728
rect 14608 34688 14614 34700
rect 14645 34697 14657 34700
rect 14691 34697 14703 34731
rect 14645 34691 14703 34697
rect 14734 34688 14740 34740
rect 14792 34688 14798 34740
rect 15378 34688 15384 34740
rect 15436 34728 15442 34740
rect 15933 34731 15991 34737
rect 15933 34728 15945 34731
rect 15436 34700 15945 34728
rect 15436 34688 15442 34700
rect 15933 34697 15945 34700
rect 15979 34697 15991 34731
rect 23198 34728 23204 34740
rect 15933 34691 15991 34697
rect 16960 34700 23204 34728
rect 12986 34620 12992 34672
rect 13044 34660 13050 34672
rect 13541 34663 13599 34669
rect 13541 34660 13553 34663
rect 13044 34632 13553 34660
rect 13044 34620 13050 34632
rect 13541 34629 13553 34632
rect 13587 34629 13599 34663
rect 13541 34623 13599 34629
rect 13906 34620 13912 34672
rect 13964 34660 13970 34672
rect 16206 34660 16212 34672
rect 13964 34632 16212 34660
rect 13964 34620 13970 34632
rect 16206 34620 16212 34632
rect 16264 34620 16270 34672
rect 16960 34669 16988 34700
rect 23198 34688 23204 34700
rect 23256 34688 23262 34740
rect 23658 34688 23664 34740
rect 23716 34728 23722 34740
rect 23753 34731 23811 34737
rect 23753 34728 23765 34731
rect 23716 34700 23765 34728
rect 23716 34688 23722 34700
rect 23753 34697 23765 34700
rect 23799 34728 23811 34731
rect 24026 34728 24032 34740
rect 23799 34700 24032 34728
rect 23799 34697 23811 34700
rect 23753 34691 23811 34697
rect 24026 34688 24032 34700
rect 24084 34688 24090 34740
rect 24394 34688 24400 34740
rect 24452 34728 24458 34740
rect 24452 34700 24808 34728
rect 24452 34688 24458 34700
rect 16945 34663 17003 34669
rect 16945 34629 16957 34663
rect 16991 34629 17003 34663
rect 20714 34660 20720 34672
rect 20562 34632 20720 34660
rect 16945 34623 17003 34629
rect 20714 34620 20720 34632
rect 20772 34620 20778 34672
rect 22281 34663 22339 34669
rect 22281 34629 22293 34663
rect 22327 34660 22339 34663
rect 22370 34660 22376 34672
rect 22327 34632 22376 34660
rect 22327 34629 22339 34632
rect 22281 34623 22339 34629
rect 22370 34620 22376 34632
rect 22428 34620 22434 34672
rect 22922 34620 22928 34672
rect 22980 34620 22986 34672
rect 24670 34620 24676 34672
rect 24728 34620 24734 34672
rect 24780 34660 24808 34700
rect 25590 34688 25596 34740
rect 25648 34728 25654 34740
rect 26145 34731 26203 34737
rect 26145 34728 26157 34731
rect 25648 34700 26157 34728
rect 25648 34688 25654 34700
rect 26145 34697 26157 34700
rect 26191 34697 26203 34731
rect 27706 34728 27712 34740
rect 26145 34691 26203 34697
rect 27080 34700 27712 34728
rect 24780 34632 25162 34660
rect 1765 34595 1823 34601
rect 1765 34561 1777 34595
rect 1811 34592 1823 34595
rect 10962 34592 10968 34604
rect 1811 34564 10968 34592
rect 1811 34561 1823 34564
rect 1765 34555 1823 34561
rect 10962 34552 10968 34564
rect 11020 34552 11026 34604
rect 13449 34595 13507 34601
rect 13449 34561 13461 34595
rect 13495 34592 13507 34595
rect 14366 34592 14372 34604
rect 13495 34564 14372 34592
rect 13495 34561 13507 34564
rect 13449 34555 13507 34561
rect 14366 34552 14372 34564
rect 14424 34552 14430 34604
rect 16025 34595 16083 34601
rect 16025 34561 16037 34595
rect 16071 34592 16083 34595
rect 16298 34592 16304 34604
rect 16071 34564 16304 34592
rect 16071 34561 16083 34564
rect 16025 34555 16083 34561
rect 16298 34552 16304 34564
rect 16356 34552 16362 34604
rect 16666 34552 16672 34604
rect 16724 34592 16730 34604
rect 17129 34595 17187 34601
rect 17129 34592 17141 34595
rect 16724 34564 17141 34592
rect 16724 34552 16730 34564
rect 17129 34561 17141 34564
rect 17175 34561 17187 34595
rect 17129 34555 17187 34561
rect 17494 34552 17500 34604
rect 17552 34592 17558 34604
rect 17552 34564 18000 34592
rect 17552 34552 17558 34564
rect 2038 34484 2044 34536
rect 2096 34484 2102 34536
rect 9582 34484 9588 34536
rect 9640 34524 9646 34536
rect 9640 34496 13584 34524
rect 9640 34484 9646 34496
rect 13556 34456 13584 34496
rect 13630 34484 13636 34536
rect 13688 34484 13694 34536
rect 14826 34484 14832 34536
rect 14884 34524 14890 34536
rect 14921 34527 14979 34533
rect 14921 34524 14933 34527
rect 14884 34496 14933 34524
rect 14884 34484 14890 34496
rect 14921 34493 14933 34496
rect 14967 34524 14979 34527
rect 15838 34524 15844 34536
rect 14967 34496 15844 34524
rect 14967 34493 14979 34496
rect 14921 34487 14979 34493
rect 15838 34484 15844 34496
rect 15896 34484 15902 34536
rect 16209 34527 16267 34533
rect 16209 34493 16221 34527
rect 16255 34493 16267 34527
rect 16209 34487 16267 34493
rect 13556 34428 14596 34456
rect 14568 34400 14596 34428
rect 15562 34416 15568 34468
rect 15620 34416 15626 34468
rect 16224 34456 16252 34487
rect 16390 34484 16396 34536
rect 16448 34524 16454 34536
rect 16448 34496 17908 34524
rect 16448 34484 16454 34496
rect 17880 34465 17908 34496
rect 17865 34459 17923 34465
rect 16224 34428 16344 34456
rect 13081 34391 13139 34397
rect 13081 34357 13093 34391
rect 13127 34388 13139 34391
rect 13354 34388 13360 34400
rect 13127 34360 13360 34388
rect 13127 34357 13139 34360
rect 13081 34351 13139 34357
rect 13354 34348 13360 34360
rect 13412 34348 13418 34400
rect 14550 34348 14556 34400
rect 14608 34388 14614 34400
rect 16316 34388 16344 34428
rect 17865 34425 17877 34459
rect 17911 34425 17923 34459
rect 17972 34456 18000 34564
rect 18230 34552 18236 34604
rect 18288 34552 18294 34604
rect 18325 34595 18383 34601
rect 18325 34561 18337 34595
rect 18371 34592 18383 34595
rect 18371 34564 18828 34592
rect 18371 34561 18383 34564
rect 18325 34555 18383 34561
rect 18417 34527 18475 34533
rect 18417 34493 18429 34527
rect 18463 34493 18475 34527
rect 18800 34524 18828 34564
rect 19058 34552 19064 34604
rect 19116 34552 19122 34604
rect 25682 34552 25688 34604
rect 25740 34592 25746 34604
rect 27080 34592 27108 34700
rect 27706 34688 27712 34700
rect 27764 34688 27770 34740
rect 27798 34688 27804 34740
rect 27856 34728 27862 34740
rect 28905 34731 28963 34737
rect 28905 34728 28917 34731
rect 27856 34700 28917 34728
rect 27856 34688 27862 34700
rect 28905 34697 28917 34700
rect 28951 34728 28963 34731
rect 30374 34728 30380 34740
rect 28951 34700 30380 34728
rect 28951 34697 28963 34700
rect 28905 34691 28963 34697
rect 30374 34688 30380 34700
rect 30432 34688 30438 34740
rect 32769 34731 32827 34737
rect 32769 34728 32781 34731
rect 30484 34700 31754 34728
rect 27430 34660 27436 34672
rect 27172 34632 27436 34660
rect 27172 34604 27200 34632
rect 27430 34620 27436 34632
rect 27488 34620 27494 34672
rect 27724 34660 27752 34688
rect 27890 34660 27896 34672
rect 27724 34632 27896 34660
rect 27890 34620 27896 34632
rect 27948 34620 27954 34672
rect 30484 34660 30512 34700
rect 28736 34632 30512 34660
rect 25740 34564 27108 34592
rect 25740 34552 25746 34564
rect 27154 34552 27160 34604
rect 27212 34552 27218 34604
rect 19334 34524 19340 34536
rect 18800 34496 19340 34524
rect 18417 34487 18475 34493
rect 18432 34456 18460 34487
rect 19334 34484 19340 34496
rect 19392 34484 19398 34536
rect 19702 34484 19708 34536
rect 19760 34524 19766 34536
rect 20622 34524 20628 34536
rect 19760 34496 20628 34524
rect 19760 34484 19766 34496
rect 20622 34484 20628 34496
rect 20680 34524 20686 34536
rect 20809 34527 20867 34533
rect 20809 34524 20821 34527
rect 20680 34496 20821 34524
rect 20680 34484 20686 34496
rect 20809 34493 20821 34496
rect 20855 34493 20867 34527
rect 20809 34487 20867 34493
rect 22002 34484 22008 34536
rect 22060 34524 22066 34536
rect 24397 34527 24455 34533
rect 24397 34524 24409 34527
rect 22060 34496 24409 34524
rect 22060 34484 22066 34496
rect 24397 34493 24409 34496
rect 24443 34493 24455 34527
rect 24397 34487 24455 34493
rect 26326 34484 26332 34536
rect 26384 34524 26390 34536
rect 28736 34524 28764 34632
rect 31202 34620 31208 34672
rect 31260 34620 31266 34672
rect 29914 34552 29920 34604
rect 29972 34552 29978 34604
rect 31726 34592 31754 34700
rect 32140 34700 32781 34728
rect 32140 34604 32168 34700
rect 32769 34697 32781 34700
rect 32815 34697 32827 34731
rect 32769 34691 32827 34697
rect 32858 34688 32864 34740
rect 32916 34728 32922 34740
rect 36630 34728 36636 34740
rect 32916 34700 36636 34728
rect 32916 34688 32922 34700
rect 36630 34688 36636 34700
rect 36688 34688 36694 34740
rect 37550 34688 37556 34740
rect 37608 34728 37614 34740
rect 38289 34731 38347 34737
rect 38289 34728 38301 34731
rect 37608 34700 38301 34728
rect 37608 34688 37614 34700
rect 38289 34697 38301 34700
rect 38335 34697 38347 34731
rect 38289 34691 38347 34697
rect 41141 34731 41199 34737
rect 41141 34697 41153 34731
rect 41187 34728 41199 34731
rect 44174 34728 44180 34740
rect 41187 34700 44180 34728
rect 41187 34697 41199 34700
rect 41141 34691 41199 34697
rect 44174 34688 44180 34700
rect 44232 34688 44238 34740
rect 47394 34688 47400 34740
rect 47452 34728 47458 34740
rect 49145 34731 49203 34737
rect 49145 34728 49157 34731
rect 47452 34700 49157 34728
rect 47452 34688 47458 34700
rect 49145 34697 49157 34700
rect 49191 34697 49203 34731
rect 49145 34691 49203 34697
rect 34054 34660 34060 34672
rect 32324 34632 34060 34660
rect 32122 34592 32128 34604
rect 31726 34564 32128 34592
rect 32122 34552 32128 34564
rect 32180 34552 32186 34604
rect 26384 34496 28764 34524
rect 26384 34484 26390 34496
rect 28810 34484 28816 34536
rect 28868 34524 28874 34536
rect 28868 34496 31524 34524
rect 28868 34484 28874 34496
rect 17972 34428 18460 34456
rect 17865 34419 17923 34425
rect 18874 34388 18880 34400
rect 14608 34360 18880 34388
rect 14608 34348 14614 34360
rect 18874 34348 18880 34360
rect 18932 34348 18938 34400
rect 19324 34391 19382 34397
rect 19324 34357 19336 34391
rect 19370 34388 19382 34391
rect 19518 34388 19524 34400
rect 19370 34360 19524 34388
rect 19370 34357 19382 34360
rect 19324 34351 19382 34357
rect 19518 34348 19524 34360
rect 19576 34388 19582 34400
rect 21634 34388 21640 34400
rect 19576 34360 21640 34388
rect 19576 34348 19582 34360
rect 21634 34348 21640 34360
rect 21692 34348 21698 34400
rect 22094 34348 22100 34400
rect 22152 34388 22158 34400
rect 22922 34388 22928 34400
rect 22152 34360 22928 34388
rect 22152 34348 22158 34360
rect 22922 34348 22928 34360
rect 22980 34388 22986 34400
rect 23842 34388 23848 34400
rect 22980 34360 23848 34388
rect 22980 34348 22986 34360
rect 23842 34348 23848 34360
rect 23900 34388 23906 34400
rect 24394 34388 24400 34400
rect 23900 34360 24400 34388
rect 23900 34348 23906 34360
rect 24394 34348 24400 34360
rect 24452 34348 24458 34400
rect 27420 34391 27478 34397
rect 27420 34357 27432 34391
rect 27466 34388 27478 34391
rect 29362 34388 29368 34400
rect 27466 34360 29368 34388
rect 27466 34357 27478 34360
rect 27420 34351 27478 34357
rect 29362 34348 29368 34360
rect 29420 34348 29426 34400
rect 29822 34348 29828 34400
rect 29880 34388 29886 34400
rect 30174 34391 30232 34397
rect 30174 34388 30186 34391
rect 29880 34360 30186 34388
rect 29880 34348 29886 34360
rect 30174 34357 30186 34360
rect 30220 34357 30232 34391
rect 31496 34388 31524 34496
rect 31662 34484 31668 34536
rect 31720 34484 31726 34536
rect 32214 34524 32220 34536
rect 31772 34496 32220 34524
rect 31570 34416 31576 34468
rect 31628 34456 31634 34468
rect 31772 34456 31800 34496
rect 32214 34484 32220 34496
rect 32272 34484 32278 34536
rect 32324 34456 32352 34632
rect 34054 34620 34060 34632
rect 34112 34620 34118 34672
rect 36262 34660 36268 34672
rect 36018 34632 36268 34660
rect 36262 34620 36268 34632
rect 36320 34620 36326 34672
rect 32677 34595 32735 34601
rect 32677 34561 32689 34595
rect 32723 34592 32735 34595
rect 34330 34592 34336 34604
rect 32723 34564 34336 34592
rect 32723 34561 32735 34564
rect 32677 34555 32735 34561
rect 34330 34552 34336 34564
rect 34388 34552 34394 34604
rect 38197 34595 38255 34601
rect 38197 34561 38209 34595
rect 38243 34592 38255 34595
rect 38562 34592 38568 34604
rect 38243 34564 38568 34592
rect 38243 34561 38255 34564
rect 38197 34555 38255 34561
rect 38562 34552 38568 34564
rect 38620 34552 38626 34604
rect 41322 34552 41328 34604
rect 41380 34552 41386 34604
rect 49326 34552 49332 34604
rect 49384 34552 49390 34604
rect 32766 34524 32772 34536
rect 31628 34428 31800 34456
rect 31864 34428 32352 34456
rect 32416 34496 32772 34524
rect 31628 34416 31634 34428
rect 31864 34388 31892 34428
rect 31496 34360 31892 34388
rect 32309 34391 32367 34397
rect 30174 34351 30232 34357
rect 32309 34357 32321 34391
rect 32355 34388 32367 34391
rect 32416 34388 32444 34496
rect 32766 34484 32772 34496
rect 32824 34484 32830 34536
rect 32953 34527 33011 34533
rect 32953 34493 32965 34527
rect 32999 34524 33011 34527
rect 33502 34524 33508 34536
rect 32999 34496 33508 34524
rect 32999 34493 33011 34496
rect 32953 34487 33011 34493
rect 33502 34484 33508 34496
rect 33560 34484 33566 34536
rect 34422 34484 34428 34536
rect 34480 34524 34486 34536
rect 34517 34527 34575 34533
rect 34517 34524 34529 34527
rect 34480 34496 34529 34524
rect 34480 34484 34486 34496
rect 34517 34493 34529 34496
rect 34563 34493 34575 34527
rect 34517 34487 34575 34493
rect 35802 34484 35808 34536
rect 35860 34524 35866 34536
rect 38381 34527 38439 34533
rect 35860 34496 37872 34524
rect 35860 34484 35866 34496
rect 32582 34416 32588 34468
rect 32640 34456 32646 34468
rect 34440 34456 34468 34484
rect 37844 34465 37872 34496
rect 38381 34493 38393 34527
rect 38427 34493 38439 34527
rect 38381 34487 38439 34493
rect 32640 34428 34468 34456
rect 37829 34459 37887 34465
rect 32640 34416 32646 34428
rect 37829 34425 37841 34459
rect 37875 34425 37887 34459
rect 37829 34419 37887 34425
rect 32355 34360 32444 34388
rect 32355 34357 32367 34360
rect 32309 34351 32367 34357
rect 33686 34348 33692 34400
rect 33744 34348 33750 34400
rect 34780 34391 34838 34397
rect 34780 34357 34792 34391
rect 34826 34388 34838 34391
rect 35986 34388 35992 34400
rect 34826 34360 35992 34388
rect 34826 34357 34838 34360
rect 34780 34351 34838 34357
rect 35986 34348 35992 34360
rect 36044 34348 36050 34400
rect 36262 34348 36268 34400
rect 36320 34388 36326 34400
rect 38396 34388 38424 34487
rect 36320 34360 38424 34388
rect 36320 34348 36326 34360
rect 1104 34298 49864 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 32950 34298
rect 33002 34246 33014 34298
rect 33066 34246 33078 34298
rect 33130 34246 33142 34298
rect 33194 34246 33206 34298
rect 33258 34246 42950 34298
rect 43002 34246 43014 34298
rect 43066 34246 43078 34298
rect 43130 34246 43142 34298
rect 43194 34246 43206 34298
rect 43258 34246 49864 34298
rect 1104 34224 49864 34246
rect 14274 34144 14280 34196
rect 14332 34144 14338 34196
rect 15488 34156 17080 34184
rect 10778 34008 10784 34060
rect 10836 34048 10842 34060
rect 11885 34051 11943 34057
rect 11885 34048 11897 34051
rect 10836 34020 11897 34048
rect 10836 34008 10842 34020
rect 11885 34017 11897 34020
rect 11931 34017 11943 34051
rect 11885 34011 11943 34017
rect 12069 34051 12127 34057
rect 12069 34017 12081 34051
rect 12115 34048 12127 34051
rect 12526 34048 12532 34060
rect 12115 34020 12532 34048
rect 12115 34017 12127 34020
rect 12069 34011 12127 34017
rect 12526 34008 12532 34020
rect 12584 34008 12590 34060
rect 14921 34051 14979 34057
rect 14921 34017 14933 34051
rect 14967 34048 14979 34051
rect 14967 34020 15148 34048
rect 14967 34017 14979 34020
rect 14921 34011 14979 34017
rect 11790 33940 11796 33992
rect 11848 33940 11854 33992
rect 13725 33983 13783 33989
rect 13725 33949 13737 33983
rect 13771 33980 13783 33983
rect 14645 33983 14703 33989
rect 14645 33980 14657 33983
rect 13771 33952 14657 33980
rect 13771 33949 13783 33952
rect 13725 33943 13783 33949
rect 14645 33949 14657 33952
rect 14691 33949 14703 33983
rect 14645 33943 14703 33949
rect 15120 33912 15148 34020
rect 15286 34008 15292 34060
rect 15344 34048 15350 34060
rect 15488 34057 15516 34156
rect 17052 34116 17080 34156
rect 17126 34144 17132 34196
rect 17184 34184 17190 34196
rect 17221 34187 17279 34193
rect 17221 34184 17233 34187
rect 17184 34156 17233 34184
rect 17184 34144 17190 34156
rect 17221 34153 17233 34156
rect 17267 34153 17279 34187
rect 19058 34184 19064 34196
rect 17221 34147 17279 34153
rect 17604 34156 19064 34184
rect 17604 34116 17632 34156
rect 19058 34144 19064 34156
rect 19116 34184 19122 34196
rect 19242 34184 19248 34196
rect 19116 34156 19248 34184
rect 19116 34144 19122 34156
rect 19242 34144 19248 34156
rect 19300 34144 19306 34196
rect 20244 34187 20302 34193
rect 20244 34153 20256 34187
rect 20290 34184 20302 34187
rect 21450 34184 21456 34196
rect 20290 34156 21456 34184
rect 20290 34153 20302 34156
rect 20244 34147 20302 34153
rect 21450 34144 21456 34156
rect 21508 34144 21514 34196
rect 21634 34144 21640 34196
rect 21692 34184 21698 34196
rect 21729 34187 21787 34193
rect 21729 34184 21741 34187
rect 21692 34156 21741 34184
rect 21692 34144 21698 34156
rect 21729 34153 21741 34156
rect 21775 34153 21787 34187
rect 21729 34147 21787 34153
rect 23566 34144 23572 34196
rect 23624 34184 23630 34196
rect 24581 34187 24639 34193
rect 24581 34184 24593 34187
rect 23624 34156 24593 34184
rect 23624 34144 23630 34156
rect 24581 34153 24593 34156
rect 24627 34153 24639 34187
rect 24581 34147 24639 34153
rect 25958 34144 25964 34196
rect 26016 34144 26022 34196
rect 28077 34187 28135 34193
rect 28077 34153 28089 34187
rect 28123 34184 28135 34187
rect 28902 34184 28908 34196
rect 28123 34156 28908 34184
rect 28123 34153 28135 34156
rect 28077 34147 28135 34153
rect 28902 34144 28908 34156
rect 28960 34144 28966 34196
rect 31726 34156 34284 34184
rect 17052 34088 17632 34116
rect 17678 34076 17684 34128
rect 17736 34116 17742 34128
rect 17736 34088 18736 34116
rect 17736 34076 17742 34088
rect 15473 34051 15531 34057
rect 15473 34048 15485 34051
rect 15344 34020 15485 34048
rect 15344 34008 15350 34020
rect 15473 34017 15485 34020
rect 15519 34017 15531 34051
rect 15473 34011 15531 34017
rect 17586 34008 17592 34060
rect 17644 34048 17650 34060
rect 18708 34057 18736 34088
rect 24118 34076 24124 34128
rect 24176 34116 24182 34128
rect 29733 34119 29791 34125
rect 29733 34116 29745 34119
rect 24176 34088 29745 34116
rect 24176 34076 24182 34088
rect 29733 34085 29745 34088
rect 29779 34085 29791 34119
rect 31726 34116 31754 34156
rect 29733 34079 29791 34085
rect 30208 34088 31754 34116
rect 34256 34116 34284 34156
rect 34330 34144 34336 34196
rect 34388 34184 34394 34196
rect 35713 34187 35771 34193
rect 35713 34184 35725 34187
rect 34388 34156 35725 34184
rect 34388 34144 34394 34156
rect 35713 34153 35725 34156
rect 35759 34153 35771 34187
rect 35713 34147 35771 34153
rect 34606 34116 34612 34128
rect 34256 34088 34612 34116
rect 18601 34051 18659 34057
rect 18601 34048 18613 34051
rect 17644 34020 18613 34048
rect 17644 34008 17650 34020
rect 18601 34017 18613 34020
rect 18647 34017 18659 34051
rect 18601 34011 18659 34017
rect 18693 34051 18751 34057
rect 18693 34017 18705 34051
rect 18739 34017 18751 34051
rect 18693 34011 18751 34017
rect 19981 34051 20039 34057
rect 19981 34017 19993 34051
rect 20027 34048 20039 34051
rect 25133 34051 25191 34057
rect 20027 34020 21588 34048
rect 20027 34017 20039 34020
rect 19981 34011 20039 34017
rect 18509 33983 18567 33989
rect 18509 33949 18521 33983
rect 18555 33980 18567 33983
rect 18782 33980 18788 33992
rect 18555 33952 18788 33980
rect 18555 33949 18567 33952
rect 18509 33943 18567 33949
rect 18782 33940 18788 33952
rect 18840 33940 18846 33992
rect 21560 33980 21588 34020
rect 25133 34017 25145 34051
rect 25179 34048 25191 34051
rect 25866 34048 25872 34060
rect 25179 34020 25872 34048
rect 25179 34017 25191 34020
rect 25133 34011 25191 34017
rect 25866 34008 25872 34020
rect 25924 34008 25930 34060
rect 28721 34051 28779 34057
rect 28721 34017 28733 34051
rect 28767 34048 28779 34051
rect 30006 34048 30012 34060
rect 28767 34020 30012 34048
rect 28767 34017 28779 34020
rect 28721 34011 28779 34017
rect 30006 34008 30012 34020
rect 30064 34008 30070 34060
rect 30208 34057 30236 34088
rect 34606 34076 34612 34088
rect 34664 34076 34670 34128
rect 34698 34076 34704 34128
rect 34756 34116 34762 34128
rect 35069 34119 35127 34125
rect 35069 34116 35081 34119
rect 34756 34088 35081 34116
rect 34756 34076 34762 34088
rect 35069 34085 35081 34088
rect 35115 34085 35127 34119
rect 35069 34079 35127 34085
rect 30193 34051 30251 34057
rect 30193 34017 30205 34051
rect 30239 34017 30251 34051
rect 30193 34011 30251 34017
rect 30285 34051 30343 34057
rect 30285 34017 30297 34051
rect 30331 34048 30343 34051
rect 31110 34048 31116 34060
rect 30331 34020 31116 34048
rect 30331 34017 30343 34020
rect 30285 34011 30343 34017
rect 31110 34008 31116 34020
rect 31168 34008 31174 34060
rect 31573 34051 31631 34057
rect 31573 34017 31585 34051
rect 31619 34048 31631 34051
rect 32398 34048 32404 34060
rect 31619 34020 32404 34048
rect 31619 34017 31631 34020
rect 31573 34011 31631 34017
rect 32398 34008 32404 34020
rect 32456 34008 32462 34060
rect 32861 34051 32919 34057
rect 32861 34017 32873 34051
rect 32907 34048 32919 34051
rect 33318 34048 33324 34060
rect 32907 34020 33324 34048
rect 32907 34017 32919 34020
rect 32861 34011 32919 34017
rect 33318 34008 33324 34020
rect 33376 34048 33382 34060
rect 34330 34048 34336 34060
rect 33376 34020 34336 34048
rect 33376 34008 33382 34020
rect 34330 34008 34336 34020
rect 34388 34008 34394 34060
rect 22002 33980 22008 33992
rect 21560 33952 22008 33980
rect 22002 33940 22008 33952
rect 22060 33980 22066 33992
rect 22925 33983 22983 33989
rect 22925 33980 22937 33983
rect 22060 33952 22937 33980
rect 22060 33940 22066 33952
rect 22925 33949 22937 33952
rect 22971 33949 22983 33983
rect 22925 33943 22983 33949
rect 23753 33983 23811 33989
rect 23753 33949 23765 33983
rect 23799 33980 23811 33983
rect 24949 33983 25007 33989
rect 24949 33980 24961 33983
rect 23799 33952 24961 33980
rect 23799 33949 23811 33952
rect 23753 33943 23811 33949
rect 24949 33949 24961 33952
rect 24995 33949 25007 33983
rect 24949 33943 25007 33949
rect 25041 33983 25099 33989
rect 25041 33949 25053 33983
rect 25087 33980 25099 33983
rect 25222 33980 25228 33992
rect 25087 33952 25228 33980
rect 25087 33949 25099 33952
rect 25041 33943 25099 33949
rect 25222 33940 25228 33952
rect 25280 33940 25286 33992
rect 27614 33940 27620 33992
rect 27672 33940 27678 33992
rect 27706 33940 27712 33992
rect 27764 33980 27770 33992
rect 28537 33983 28595 33989
rect 28537 33980 28549 33983
rect 27764 33952 28549 33980
rect 27764 33940 27770 33952
rect 28537 33949 28549 33952
rect 28583 33949 28595 33983
rect 28537 33943 28595 33949
rect 28810 33940 28816 33992
rect 28868 33980 28874 33992
rect 30101 33983 30159 33989
rect 30101 33980 30113 33983
rect 28868 33952 30113 33980
rect 28868 33940 28874 33952
rect 30101 33949 30113 33952
rect 30147 33949 30159 33983
rect 30101 33943 30159 33949
rect 31297 33983 31355 33989
rect 31297 33949 31309 33983
rect 31343 33980 31355 33983
rect 31343 33952 31754 33980
rect 31343 33949 31355 33952
rect 31297 33943 31355 33949
rect 15749 33915 15807 33921
rect 15749 33912 15761 33915
rect 11440 33884 12434 33912
rect 15120 33884 15761 33912
rect 11440 33853 11468 33884
rect 11425 33847 11483 33853
rect 11425 33813 11437 33847
rect 11471 33813 11483 33847
rect 12406 33844 12434 33884
rect 15749 33881 15761 33884
rect 15795 33881 15807 33915
rect 15749 33875 15807 33881
rect 14458 33844 14464 33856
rect 12406 33816 14464 33844
rect 11425 33807 11483 33813
rect 14458 33804 14464 33816
rect 14516 33804 14522 33856
rect 14737 33847 14795 33853
rect 14737 33813 14749 33847
rect 14783 33844 14795 33847
rect 15378 33844 15384 33856
rect 14783 33816 15384 33844
rect 14783 33813 14795 33816
rect 14737 33807 14795 33813
rect 15378 33804 15384 33816
rect 15436 33804 15442 33856
rect 15764 33844 15792 33875
rect 16022 33872 16028 33924
rect 16080 33912 16086 33924
rect 20162 33912 20168 33924
rect 16080 33884 16238 33912
rect 18616 33884 20168 33912
rect 16080 33872 16086 33884
rect 16574 33844 16580 33856
rect 15764 33816 16580 33844
rect 16574 33804 16580 33816
rect 16632 33804 16638 33856
rect 18141 33847 18199 33853
rect 18141 33813 18153 33847
rect 18187 33844 18199 33847
rect 18616 33844 18644 33884
rect 20162 33872 20168 33884
rect 20220 33872 20226 33924
rect 20714 33872 20720 33924
rect 20772 33872 20778 33924
rect 22189 33915 22247 33921
rect 22189 33912 22201 33915
rect 22066 33884 22201 33912
rect 18187 33816 18644 33844
rect 18187 33813 18199 33816
rect 18141 33807 18199 33813
rect 18782 33804 18788 33856
rect 18840 33844 18846 33856
rect 22066 33844 22094 33884
rect 22189 33881 22201 33884
rect 22235 33881 22247 33915
rect 22189 33875 22247 33881
rect 28445 33915 28503 33921
rect 28445 33881 28457 33915
rect 28491 33912 28503 33915
rect 29546 33912 29552 33924
rect 28491 33884 29552 33912
rect 28491 33881 28503 33884
rect 28445 33875 28503 33881
rect 29546 33872 29552 33884
rect 29604 33872 29610 33924
rect 31726 33912 31754 33952
rect 32490 33940 32496 33992
rect 32548 33980 32554 33992
rect 32585 33983 32643 33989
rect 32585 33980 32597 33983
rect 32548 33952 32597 33980
rect 32548 33940 32554 33952
rect 32585 33949 32597 33952
rect 32631 33949 32643 33983
rect 32585 33943 32643 33949
rect 34146 33940 34152 33992
rect 34204 33980 34210 33992
rect 36078 33980 36084 33992
rect 34204 33952 36084 33980
rect 34204 33940 34210 33952
rect 36078 33940 36084 33952
rect 36136 33940 36142 33992
rect 32398 33912 32404 33924
rect 30944 33884 31524 33912
rect 31726 33884 32404 33912
rect 18840 33816 22094 33844
rect 18840 33804 18846 33816
rect 30098 33804 30104 33856
rect 30156 33844 30162 33856
rect 30834 33844 30840 33856
rect 30156 33816 30840 33844
rect 30156 33804 30162 33816
rect 30834 33804 30840 33816
rect 30892 33804 30898 33856
rect 30944 33853 30972 33884
rect 30929 33847 30987 33853
rect 30929 33813 30941 33847
rect 30975 33813 30987 33847
rect 30929 33807 30987 33813
rect 31018 33804 31024 33856
rect 31076 33844 31082 33856
rect 31389 33847 31447 33853
rect 31389 33844 31401 33847
rect 31076 33816 31401 33844
rect 31076 33804 31082 33816
rect 31389 33813 31401 33816
rect 31435 33813 31447 33847
rect 31496 33844 31524 33884
rect 32398 33872 32404 33884
rect 32456 33872 32462 33924
rect 33134 33872 33140 33924
rect 33192 33912 33198 33924
rect 33192 33884 33350 33912
rect 33192 33872 33198 33884
rect 33042 33844 33048 33856
rect 31496 33816 33048 33844
rect 31389 33807 31447 33813
rect 33042 33804 33048 33816
rect 33100 33804 33106 33856
rect 33226 33804 33232 33856
rect 33284 33844 33290 33856
rect 34333 33847 34391 33853
rect 34333 33844 34345 33847
rect 33284 33816 34345 33844
rect 33284 33804 33290 33816
rect 34333 33813 34345 33816
rect 34379 33844 34391 33847
rect 35526 33844 35532 33856
rect 34379 33816 35532 33844
rect 34379 33813 34391 33816
rect 34333 33807 34391 33813
rect 35526 33804 35532 33816
rect 35584 33804 35590 33856
rect 1104 33754 49864 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 27950 33754
rect 28002 33702 28014 33754
rect 28066 33702 28078 33754
rect 28130 33702 28142 33754
rect 28194 33702 28206 33754
rect 28258 33702 37950 33754
rect 38002 33702 38014 33754
rect 38066 33702 38078 33754
rect 38130 33702 38142 33754
rect 38194 33702 38206 33754
rect 38258 33702 47950 33754
rect 48002 33702 48014 33754
rect 48066 33702 48078 33754
rect 48130 33702 48142 33754
rect 48194 33702 48206 33754
rect 48258 33702 49864 33754
rect 1104 33680 49864 33702
rect 14366 33600 14372 33652
rect 14424 33600 14430 33652
rect 14737 33643 14795 33649
rect 14737 33609 14749 33643
rect 14783 33640 14795 33643
rect 16390 33640 16396 33652
rect 14783 33612 16396 33640
rect 14783 33609 14795 33612
rect 14737 33603 14795 33609
rect 16390 33600 16396 33612
rect 16448 33600 16454 33652
rect 17773 33643 17831 33649
rect 17773 33609 17785 33643
rect 17819 33640 17831 33643
rect 17862 33640 17868 33652
rect 17819 33612 17868 33640
rect 17819 33609 17831 33612
rect 17773 33603 17831 33609
rect 17862 33600 17868 33612
rect 17920 33600 17926 33652
rect 20530 33600 20536 33652
rect 20588 33640 20594 33652
rect 20717 33643 20775 33649
rect 20717 33640 20729 33643
rect 20588 33612 20729 33640
rect 20588 33600 20594 33612
rect 20717 33609 20729 33612
rect 20763 33609 20775 33643
rect 20717 33603 20775 33609
rect 21082 33600 21088 33652
rect 21140 33600 21146 33652
rect 22094 33600 22100 33652
rect 22152 33640 22158 33652
rect 22152 33612 22692 33640
rect 22152 33600 22158 33612
rect 14182 33532 14188 33584
rect 14240 33572 14246 33584
rect 16025 33575 16083 33581
rect 16025 33572 16037 33575
rect 14240 33544 16037 33572
rect 14240 33532 14246 33544
rect 16025 33541 16037 33544
rect 16071 33541 16083 33575
rect 16025 33535 16083 33541
rect 17678 33532 17684 33584
rect 17736 33572 17742 33584
rect 17736 33544 18552 33572
rect 17736 33532 17742 33544
rect 1765 33507 1823 33513
rect 1765 33473 1777 33507
rect 1811 33504 1823 33507
rect 8570 33504 8576 33516
rect 1811 33476 8576 33504
rect 1811 33473 1823 33476
rect 1765 33467 1823 33473
rect 8570 33464 8576 33476
rect 8628 33464 8634 33516
rect 13538 33464 13544 33516
rect 13596 33504 13602 33516
rect 15933 33507 15991 33513
rect 13596 33476 14964 33504
rect 13596 33464 13602 33476
rect 1302 33396 1308 33448
rect 1360 33436 1366 33448
rect 2041 33439 2099 33445
rect 2041 33436 2053 33439
rect 1360 33408 2053 33436
rect 1360 33396 1366 33408
rect 2041 33405 2053 33408
rect 2087 33405 2099 33439
rect 2041 33399 2099 33405
rect 14642 33396 14648 33448
rect 14700 33436 14706 33448
rect 14936 33445 14964 33476
rect 15933 33473 15945 33507
rect 15979 33504 15991 33507
rect 16482 33504 16488 33516
rect 15979 33476 16488 33504
rect 15979 33473 15991 33476
rect 15933 33467 15991 33473
rect 16482 33464 16488 33476
rect 16540 33464 16546 33516
rect 17865 33507 17923 33513
rect 17865 33473 17877 33507
rect 17911 33504 17923 33507
rect 18414 33504 18420 33516
rect 17911 33476 18420 33504
rect 17911 33473 17923 33476
rect 17865 33467 17923 33473
rect 18414 33464 18420 33476
rect 18472 33464 18478 33516
rect 18524 33504 18552 33544
rect 18598 33532 18604 33584
rect 18656 33572 18662 33584
rect 18782 33572 18788 33584
rect 18656 33544 18788 33572
rect 18656 33532 18662 33544
rect 18782 33532 18788 33544
rect 18840 33532 18846 33584
rect 19058 33532 19064 33584
rect 19116 33572 19122 33584
rect 19242 33572 19248 33584
rect 19116 33544 19248 33572
rect 19116 33532 19122 33544
rect 19242 33532 19248 33544
rect 19300 33572 19306 33584
rect 19337 33575 19395 33581
rect 19337 33572 19349 33575
rect 19300 33544 19349 33572
rect 19300 33532 19306 33544
rect 19337 33541 19349 33544
rect 19383 33541 19395 33575
rect 19337 33535 19395 33541
rect 21177 33575 21235 33581
rect 21177 33541 21189 33575
rect 21223 33572 21235 33575
rect 21266 33572 21272 33584
rect 21223 33544 21272 33572
rect 21223 33541 21235 33544
rect 21177 33535 21235 33541
rect 21266 33532 21272 33544
rect 21324 33532 21330 33584
rect 21358 33532 21364 33584
rect 21416 33572 21422 33584
rect 22278 33572 22284 33584
rect 21416 33544 22284 33572
rect 21416 33532 21422 33544
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 22664 33572 22692 33612
rect 23934 33600 23940 33652
rect 23992 33640 23998 33652
rect 26053 33643 26111 33649
rect 26053 33640 26065 33643
rect 23992 33612 26065 33640
rect 23992 33600 23998 33612
rect 26053 33609 26065 33612
rect 26099 33609 26111 33643
rect 31110 33640 31116 33652
rect 26053 33603 26111 33609
rect 27448 33612 31116 33640
rect 24578 33572 24584 33584
rect 22664 33544 22770 33572
rect 24320 33544 24584 33572
rect 20990 33504 20996 33516
rect 18524 33476 20996 33504
rect 20990 33464 20996 33476
rect 21048 33464 21054 33516
rect 24320 33513 24348 33544
rect 24578 33532 24584 33544
rect 24636 33532 24642 33584
rect 24670 33532 24676 33584
rect 24728 33572 24734 33584
rect 27448 33581 27476 33612
rect 31110 33600 31116 33612
rect 31168 33600 31174 33652
rect 31202 33600 31208 33652
rect 31260 33640 31266 33652
rect 33134 33640 33140 33652
rect 31260 33612 33140 33640
rect 31260 33600 31266 33612
rect 33134 33600 33140 33612
rect 33192 33640 33198 33652
rect 33192 33612 33456 33640
rect 33192 33600 33198 33612
rect 27433 33575 27491 33581
rect 24728 33544 25070 33572
rect 24728 33532 24734 33544
rect 27433 33541 27445 33575
rect 27479 33541 27491 33575
rect 27433 33535 27491 33541
rect 27890 33532 27896 33584
rect 27948 33532 27954 33584
rect 30742 33532 30748 33584
rect 30800 33532 30806 33584
rect 33428 33572 33456 33612
rect 33686 33600 33692 33652
rect 33744 33640 33750 33652
rect 36262 33640 36268 33652
rect 33744 33612 36268 33640
rect 33744 33600 33750 33612
rect 36262 33600 36268 33612
rect 36320 33600 36326 33652
rect 33778 33572 33784 33584
rect 33428 33544 33784 33572
rect 33778 33532 33784 33544
rect 33836 33532 33842 33584
rect 24305 33507 24363 33513
rect 24305 33473 24317 33507
rect 24351 33473 24363 33507
rect 24305 33467 24363 33473
rect 27154 33464 27160 33516
rect 27212 33464 27218 33516
rect 29546 33464 29552 33516
rect 29604 33464 29610 33516
rect 29730 33464 29736 33516
rect 29788 33504 29794 33516
rect 30006 33504 30012 33516
rect 29788 33476 30012 33504
rect 29788 33464 29794 33476
rect 30006 33464 30012 33476
rect 30064 33464 30070 33516
rect 32398 33464 32404 33516
rect 32456 33504 32462 33516
rect 32493 33507 32551 33513
rect 32493 33504 32505 33507
rect 32456 33476 32505 33504
rect 32456 33464 32462 33476
rect 32493 33473 32505 33476
rect 32539 33473 32551 33507
rect 32493 33467 32551 33473
rect 39666 33464 39672 33516
rect 39724 33464 39730 33516
rect 39850 33464 39856 33516
rect 39908 33504 39914 33516
rect 41049 33507 41107 33513
rect 41049 33504 41061 33507
rect 39908 33476 41061 33504
rect 39908 33464 39914 33476
rect 41049 33473 41061 33476
rect 41095 33473 41107 33507
rect 41049 33467 41107 33473
rect 49142 33464 49148 33516
rect 49200 33464 49206 33516
rect 14829 33439 14887 33445
rect 14829 33436 14841 33439
rect 14700 33408 14841 33436
rect 14700 33396 14706 33408
rect 14829 33405 14841 33408
rect 14875 33405 14887 33439
rect 14829 33399 14887 33405
rect 14921 33439 14979 33445
rect 14921 33405 14933 33439
rect 14967 33405 14979 33439
rect 14921 33399 14979 33405
rect 16209 33439 16267 33445
rect 16209 33405 16221 33439
rect 16255 33436 16267 33439
rect 17678 33436 17684 33448
rect 16255 33408 17684 33436
rect 16255 33405 16267 33408
rect 16209 33399 16267 33405
rect 17678 33396 17684 33408
rect 17736 33396 17742 33448
rect 17770 33396 17776 33448
rect 17828 33436 17834 33448
rect 17957 33439 18015 33445
rect 17957 33436 17969 33439
rect 17828 33408 17969 33436
rect 17828 33396 17834 33408
rect 17957 33405 17969 33408
rect 18003 33436 18015 33439
rect 18782 33436 18788 33448
rect 18003 33408 18788 33436
rect 18003 33405 18015 33408
rect 17957 33399 18015 33405
rect 18782 33396 18788 33408
rect 18840 33396 18846 33448
rect 21269 33439 21327 33445
rect 21269 33405 21281 33439
rect 21315 33405 21327 33439
rect 21269 33399 21327 33405
rect 15565 33371 15623 33377
rect 15565 33337 15577 33371
rect 15611 33368 15623 33371
rect 19242 33368 19248 33380
rect 15611 33340 19248 33368
rect 15611 33337 15623 33340
rect 15565 33331 15623 33337
rect 19242 33328 19248 33340
rect 19300 33328 19306 33380
rect 17402 33260 17408 33312
rect 17460 33260 17466 33312
rect 17862 33260 17868 33312
rect 17920 33300 17926 33312
rect 21284 33300 21312 33399
rect 21358 33396 21364 33448
rect 21416 33436 21422 33448
rect 22002 33436 22008 33448
rect 21416 33408 22008 33436
rect 21416 33396 21422 33408
rect 22002 33396 22008 33408
rect 22060 33396 22066 33448
rect 22278 33396 22284 33448
rect 22336 33436 22342 33448
rect 24026 33436 24032 33448
rect 22336 33408 24032 33436
rect 22336 33396 22342 33408
rect 24026 33396 24032 33408
rect 24084 33396 24090 33448
rect 24581 33439 24639 33445
rect 24581 33405 24593 33439
rect 24627 33436 24639 33439
rect 25222 33436 25228 33448
rect 24627 33408 25228 33436
rect 24627 33405 24639 33408
rect 24581 33399 24639 33405
rect 25222 33396 25228 33408
rect 25280 33436 25286 33448
rect 25590 33436 25596 33448
rect 25280 33408 25596 33436
rect 25280 33396 25286 33408
rect 25590 33396 25596 33408
rect 25648 33396 25654 33448
rect 30285 33439 30343 33445
rect 30285 33405 30297 33439
rect 30331 33436 30343 33439
rect 31662 33436 31668 33448
rect 30331 33408 31668 33436
rect 30331 33405 30343 33408
rect 30285 33399 30343 33405
rect 31662 33396 31668 33408
rect 31720 33396 31726 33448
rect 32582 33396 32588 33448
rect 32640 33436 32646 33448
rect 33045 33439 33103 33445
rect 33045 33436 33057 33439
rect 32640 33408 33057 33436
rect 32640 33396 32646 33408
rect 33045 33405 33057 33408
rect 33091 33405 33103 33439
rect 33045 33399 33103 33405
rect 33321 33439 33379 33445
rect 33321 33405 33333 33439
rect 33367 33436 33379 33439
rect 33686 33436 33692 33448
rect 33367 33408 33692 33436
rect 33367 33405 33379 33408
rect 33321 33399 33379 33405
rect 33686 33396 33692 33408
rect 33744 33396 33750 33448
rect 34054 33396 34060 33448
rect 34112 33436 34118 33448
rect 49329 33439 49387 33445
rect 49329 33436 49341 33439
rect 34112 33408 49341 33436
rect 34112 33396 34118 33408
rect 49329 33405 49341 33408
rect 49375 33405 49387 33439
rect 49329 33399 49387 33405
rect 34330 33328 34336 33380
rect 34388 33368 34394 33380
rect 34793 33371 34851 33377
rect 34793 33368 34805 33371
rect 34388 33340 34805 33368
rect 34388 33328 34394 33340
rect 34793 33337 34805 33340
rect 34839 33337 34851 33371
rect 34793 33331 34851 33337
rect 39485 33371 39543 33377
rect 39485 33337 39497 33371
rect 39531 33368 39543 33371
rect 44082 33368 44088 33380
rect 39531 33340 44088 33368
rect 39531 33337 39543 33340
rect 39485 33331 39543 33337
rect 44082 33328 44088 33340
rect 44140 33328 44146 33380
rect 17920 33272 21312 33300
rect 17920 33260 17926 33272
rect 21450 33260 21456 33312
rect 21508 33300 21514 33312
rect 21634 33300 21640 33312
rect 21508 33272 21640 33300
rect 21508 33260 21514 33272
rect 21634 33260 21640 33272
rect 21692 33300 21698 33312
rect 23753 33303 23811 33309
rect 23753 33300 23765 33303
rect 21692 33272 23765 33300
rect 21692 33260 21698 33272
rect 23753 33269 23765 33272
rect 23799 33269 23811 33303
rect 23753 33263 23811 33269
rect 27246 33260 27252 33312
rect 27304 33300 27310 33312
rect 28905 33303 28963 33309
rect 28905 33300 28917 33303
rect 27304 33272 28917 33300
rect 27304 33260 27310 33272
rect 28905 33269 28917 33272
rect 28951 33269 28963 33303
rect 28905 33263 28963 33269
rect 30466 33260 30472 33312
rect 30524 33300 30530 33312
rect 30742 33300 30748 33312
rect 30524 33272 30748 33300
rect 30524 33260 30530 33272
rect 30742 33260 30748 33272
rect 30800 33260 30806 33312
rect 30834 33260 30840 33312
rect 30892 33300 30898 33312
rect 31757 33303 31815 33309
rect 31757 33300 31769 33303
rect 30892 33272 31769 33300
rect 30892 33260 30898 33272
rect 31757 33269 31769 33272
rect 31803 33269 31815 33303
rect 31757 33263 31815 33269
rect 33042 33260 33048 33312
rect 33100 33300 33106 33312
rect 36170 33300 36176 33312
rect 33100 33272 36176 33300
rect 33100 33260 33106 33272
rect 36170 33260 36176 33272
rect 36228 33260 36234 33312
rect 40865 33303 40923 33309
rect 40865 33269 40877 33303
rect 40911 33300 40923 33303
rect 45830 33300 45836 33312
rect 40911 33272 45836 33300
rect 40911 33269 40923 33272
rect 40865 33263 40923 33269
rect 45830 33260 45836 33272
rect 45888 33260 45894 33312
rect 1104 33210 49864 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 32950 33210
rect 33002 33158 33014 33210
rect 33066 33158 33078 33210
rect 33130 33158 33142 33210
rect 33194 33158 33206 33210
rect 33258 33158 42950 33210
rect 43002 33158 43014 33210
rect 43066 33158 43078 33210
rect 43130 33158 43142 33210
rect 43194 33158 43206 33210
rect 43258 33158 49864 33210
rect 1104 33136 49864 33158
rect 16666 33096 16672 33108
rect 2746 33068 16672 33096
rect 1302 32920 1308 32972
rect 1360 32960 1366 32972
rect 2041 32963 2099 32969
rect 2041 32960 2053 32963
rect 1360 32932 2053 32960
rect 1360 32920 1366 32932
rect 2041 32929 2053 32932
rect 2087 32929 2099 32963
rect 2041 32923 2099 32929
rect 1765 32895 1823 32901
rect 1765 32861 1777 32895
rect 1811 32892 1823 32895
rect 2746 32892 2774 33068
rect 16666 33056 16672 33068
rect 16724 33056 16730 33108
rect 18414 33056 18420 33108
rect 18472 33096 18478 33108
rect 18690 33096 18696 33108
rect 18472 33068 18696 33096
rect 18472 33056 18478 33068
rect 18690 33056 18696 33068
rect 18748 33056 18754 33108
rect 18966 33056 18972 33108
rect 19024 33096 19030 33108
rect 19613 33099 19671 33105
rect 19613 33096 19625 33099
rect 19024 33068 19625 33096
rect 19024 33056 19030 33068
rect 19613 33065 19625 33068
rect 19659 33065 19671 33099
rect 19613 33059 19671 33065
rect 19720 33068 22692 33096
rect 15286 32920 15292 32972
rect 15344 32960 15350 32972
rect 15933 32963 15991 32969
rect 15933 32960 15945 32963
rect 15344 32932 15945 32960
rect 15344 32920 15350 32932
rect 15933 32929 15945 32932
rect 15979 32929 15991 32963
rect 15933 32923 15991 32929
rect 16206 32920 16212 32972
rect 16264 32960 16270 32972
rect 19720 32960 19748 33068
rect 20070 32988 20076 33040
rect 20128 33028 20134 33040
rect 20165 33031 20223 33037
rect 20165 33028 20177 33031
rect 20128 33000 20177 33028
rect 20128 32988 20134 33000
rect 20165 32997 20177 33000
rect 20211 32997 20223 33031
rect 22664 33028 22692 33068
rect 22922 33056 22928 33108
rect 22980 33096 22986 33108
rect 23109 33099 23167 33105
rect 23109 33096 23121 33099
rect 22980 33068 23121 33096
rect 22980 33056 22986 33068
rect 23109 33065 23121 33068
rect 23155 33065 23167 33099
rect 23109 33059 23167 33065
rect 24581 33099 24639 33105
rect 24581 33065 24593 33099
rect 24627 33096 24639 33099
rect 24854 33096 24860 33108
rect 24627 33068 24860 33096
rect 24627 33065 24639 33068
rect 24581 33059 24639 33065
rect 24854 33056 24860 33068
rect 24912 33056 24918 33108
rect 27617 33099 27675 33105
rect 27617 33065 27629 33099
rect 27663 33096 27675 33099
rect 31570 33096 31576 33108
rect 27663 33068 31576 33096
rect 27663 33065 27675 33068
rect 27617 33059 27675 33065
rect 31570 33056 31576 33068
rect 31628 33056 31634 33108
rect 49237 33099 49295 33105
rect 49237 33096 49249 33099
rect 31726 33068 49249 33096
rect 23566 33028 23572 33040
rect 22664 33000 23572 33028
rect 20165 32991 20223 32997
rect 23566 32988 23572 33000
rect 23624 32988 23630 33040
rect 31294 32988 31300 33040
rect 31352 33028 31358 33040
rect 31726 33028 31754 33068
rect 49237 33065 49249 33068
rect 49283 33065 49295 33099
rect 49237 33059 49295 33065
rect 31352 33000 31754 33028
rect 32125 33031 32183 33037
rect 31352 32988 31358 33000
rect 32125 32997 32137 33031
rect 32171 33028 32183 33031
rect 32171 33000 32720 33028
rect 32171 32997 32183 33000
rect 32125 32991 32183 32997
rect 16264 32932 19748 32960
rect 16264 32920 16270 32932
rect 20622 32920 20628 32972
rect 20680 32960 20686 32972
rect 20717 32963 20775 32969
rect 20717 32960 20729 32963
rect 20680 32932 20729 32960
rect 20680 32920 20686 32932
rect 20717 32929 20729 32932
rect 20763 32929 20775 32963
rect 20717 32923 20775 32929
rect 21637 32963 21695 32969
rect 21637 32929 21649 32963
rect 21683 32960 21695 32963
rect 23658 32960 23664 32972
rect 21683 32932 23664 32960
rect 21683 32929 21695 32932
rect 21637 32923 21695 32929
rect 23658 32920 23664 32932
rect 23716 32920 23722 32972
rect 25225 32963 25283 32969
rect 25225 32929 25237 32963
rect 25271 32960 25283 32963
rect 27246 32960 27252 32972
rect 25271 32932 27252 32960
rect 25271 32929 25283 32932
rect 25225 32923 25283 32929
rect 27246 32920 27252 32932
rect 27304 32920 27310 32972
rect 28261 32963 28319 32969
rect 27356 32932 28212 32960
rect 1811 32864 2774 32892
rect 1811 32861 1823 32864
rect 1765 32855 1823 32861
rect 13538 32852 13544 32904
rect 13596 32892 13602 32904
rect 14829 32895 14887 32901
rect 14829 32892 14841 32895
rect 13596 32864 14841 32892
rect 13596 32852 13602 32864
rect 14829 32861 14841 32864
rect 14875 32861 14887 32895
rect 14829 32855 14887 32861
rect 20530 32852 20536 32904
rect 20588 32852 20594 32904
rect 21358 32852 21364 32904
rect 21416 32852 21422 32904
rect 24029 32895 24087 32901
rect 24029 32861 24041 32895
rect 24075 32892 24087 32895
rect 24949 32895 25007 32901
rect 24949 32892 24961 32895
rect 24075 32864 24961 32892
rect 24075 32861 24087 32864
rect 24029 32855 24087 32861
rect 24949 32861 24961 32864
rect 24995 32861 25007 32895
rect 25406 32892 25412 32904
rect 24949 32855 25007 32861
rect 25056 32864 25412 32892
rect 15930 32784 15936 32836
rect 15988 32824 15994 32836
rect 16209 32827 16267 32833
rect 16209 32824 16221 32827
rect 15988 32796 16221 32824
rect 15988 32784 15994 32796
rect 16209 32793 16221 32796
rect 16255 32793 16267 32827
rect 16209 32787 16267 32793
rect 16408 32796 16698 32824
rect 16408 32768 16436 32796
rect 20070 32784 20076 32836
rect 20128 32824 20134 32836
rect 20714 32824 20720 32836
rect 20128 32796 20720 32824
rect 20128 32784 20134 32796
rect 20714 32784 20720 32796
rect 20772 32824 20778 32836
rect 22094 32824 22100 32836
rect 20772 32796 22100 32824
rect 20772 32784 20778 32796
rect 22094 32784 22100 32796
rect 22152 32784 22158 32836
rect 23566 32784 23572 32836
rect 23624 32824 23630 32836
rect 25056 32824 25084 32864
rect 25406 32852 25412 32864
rect 25464 32892 25470 32904
rect 27356 32892 27384 32932
rect 25464 32864 27384 32892
rect 25464 32852 25470 32864
rect 27614 32852 27620 32904
rect 27672 32892 27678 32904
rect 27985 32895 28043 32901
rect 27985 32892 27997 32895
rect 27672 32864 27997 32892
rect 27672 32852 27678 32864
rect 27985 32861 27997 32864
rect 28031 32861 28043 32895
rect 27985 32855 28043 32861
rect 23624 32796 25084 32824
rect 23624 32784 23630 32796
rect 25314 32784 25320 32836
rect 25372 32824 25378 32836
rect 28077 32827 28135 32833
rect 28077 32824 28089 32827
rect 25372 32796 28089 32824
rect 25372 32784 25378 32796
rect 28077 32793 28089 32796
rect 28123 32793 28135 32827
rect 28184 32824 28212 32932
rect 28261 32929 28273 32963
rect 28307 32960 28319 32963
rect 28350 32960 28356 32972
rect 28307 32932 28356 32960
rect 28307 32929 28319 32932
rect 28261 32923 28319 32929
rect 28350 32920 28356 32932
rect 28408 32920 28414 32972
rect 28626 32920 28632 32972
rect 28684 32960 28690 32972
rect 30009 32963 30067 32969
rect 30009 32960 30021 32963
rect 28684 32932 30021 32960
rect 28684 32920 28690 32932
rect 30009 32929 30021 32932
rect 30055 32960 30067 32963
rect 30098 32960 30104 32972
rect 30055 32932 30104 32960
rect 30055 32929 30067 32932
rect 30009 32923 30067 32929
rect 30098 32920 30104 32932
rect 30156 32920 30162 32972
rect 30466 32920 30472 32972
rect 30524 32960 30530 32972
rect 31202 32960 31208 32972
rect 30524 32932 31208 32960
rect 30524 32920 30530 32932
rect 31202 32920 31208 32932
rect 31260 32920 31266 32972
rect 32582 32920 32588 32972
rect 32640 32920 32646 32972
rect 32692 32960 32720 33000
rect 33502 32960 33508 32972
rect 32692 32932 33508 32960
rect 33502 32920 33508 32932
rect 33560 32920 33566 32972
rect 29178 32852 29184 32904
rect 29236 32852 29242 32904
rect 29730 32852 29736 32904
rect 29788 32852 29794 32904
rect 49050 32852 49056 32904
rect 49108 32852 49114 32904
rect 30282 32824 30288 32836
rect 28184 32796 30288 32824
rect 28077 32787 28135 32793
rect 30282 32784 30288 32796
rect 30340 32784 30346 32836
rect 30466 32784 30472 32836
rect 30524 32784 30530 32836
rect 31846 32784 31852 32836
rect 31904 32824 31910 32836
rect 32861 32827 32919 32833
rect 31904 32796 32812 32824
rect 31904 32784 31910 32796
rect 16390 32716 16396 32768
rect 16448 32716 16454 32768
rect 17126 32716 17132 32768
rect 17184 32756 17190 32768
rect 17494 32756 17500 32768
rect 17184 32728 17500 32756
rect 17184 32716 17190 32728
rect 17494 32716 17500 32728
rect 17552 32756 17558 32768
rect 17681 32759 17739 32765
rect 17681 32756 17693 32759
rect 17552 32728 17693 32756
rect 17552 32716 17558 32728
rect 17681 32725 17693 32728
rect 17727 32725 17739 32759
rect 17681 32719 17739 32725
rect 19334 32716 19340 32768
rect 19392 32756 19398 32768
rect 20438 32756 20444 32768
rect 19392 32728 20444 32756
rect 19392 32716 19398 32728
rect 20438 32716 20444 32728
rect 20496 32756 20502 32768
rect 20622 32756 20628 32768
rect 20496 32728 20628 32756
rect 20496 32716 20502 32728
rect 20622 32716 20628 32728
rect 20680 32716 20686 32768
rect 23842 32716 23848 32768
rect 23900 32756 23906 32768
rect 25041 32759 25099 32765
rect 25041 32756 25053 32759
rect 23900 32728 25053 32756
rect 23900 32716 23906 32728
rect 25041 32725 25053 32728
rect 25087 32756 25099 32759
rect 27614 32756 27620 32768
rect 25087 32728 27620 32756
rect 25087 32725 25099 32728
rect 25041 32719 25099 32725
rect 27614 32716 27620 32728
rect 27672 32716 27678 32768
rect 28534 32716 28540 32768
rect 28592 32756 28598 32768
rect 31481 32759 31539 32765
rect 31481 32756 31493 32759
rect 28592 32728 31493 32756
rect 28592 32716 28598 32728
rect 31481 32725 31493 32728
rect 31527 32756 31539 32759
rect 32122 32756 32128 32768
rect 31527 32728 32128 32756
rect 31527 32725 31539 32728
rect 31481 32719 31539 32725
rect 32122 32716 32128 32728
rect 32180 32716 32186 32768
rect 32784 32756 32812 32796
rect 32861 32793 32873 32827
rect 32907 32824 32919 32827
rect 33134 32824 33140 32836
rect 32907 32796 33140 32824
rect 32907 32793 32919 32796
rect 32861 32787 32919 32793
rect 33134 32784 33140 32796
rect 33192 32784 33198 32836
rect 33870 32784 33876 32836
rect 33928 32784 33934 32836
rect 34333 32759 34391 32765
rect 34333 32756 34345 32759
rect 32784 32728 34345 32756
rect 34333 32725 34345 32728
rect 34379 32756 34391 32759
rect 36722 32756 36728 32768
rect 34379 32728 36728 32756
rect 34379 32725 34391 32728
rect 34333 32719 34391 32725
rect 36722 32716 36728 32728
rect 36780 32716 36786 32768
rect 1104 32666 49864 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 27950 32666
rect 28002 32614 28014 32666
rect 28066 32614 28078 32666
rect 28130 32614 28142 32666
rect 28194 32614 28206 32666
rect 28258 32614 37950 32666
rect 38002 32614 38014 32666
rect 38066 32614 38078 32666
rect 38130 32614 38142 32666
rect 38194 32614 38206 32666
rect 38258 32614 47950 32666
rect 48002 32614 48014 32666
rect 48066 32614 48078 32666
rect 48130 32614 48142 32666
rect 48194 32614 48206 32666
rect 48258 32614 49864 32666
rect 1104 32592 49864 32614
rect 12802 32512 12808 32564
rect 12860 32552 12866 32564
rect 12897 32555 12955 32561
rect 12897 32552 12909 32555
rect 12860 32524 12909 32552
rect 12860 32512 12866 32524
rect 12897 32521 12909 32524
rect 12943 32521 12955 32555
rect 16206 32552 16212 32564
rect 12897 32515 12955 32521
rect 14200 32524 16212 32552
rect 12437 32487 12495 32493
rect 12437 32484 12449 32487
rect 2746 32456 12449 32484
rect 1854 32172 1860 32224
rect 1912 32212 1918 32224
rect 2746 32212 2774 32456
rect 12437 32453 12449 32456
rect 12483 32484 12495 32487
rect 13265 32487 13323 32493
rect 13265 32484 13277 32487
rect 12483 32456 13277 32484
rect 12483 32453 12495 32456
rect 12437 32447 12495 32453
rect 13265 32453 13277 32456
rect 13311 32453 13323 32487
rect 13265 32447 13323 32453
rect 12621 32419 12679 32425
rect 12621 32385 12633 32419
rect 12667 32416 12679 32419
rect 14200 32416 14228 32524
rect 16206 32512 16212 32524
rect 16264 32512 16270 32564
rect 20254 32552 20260 32564
rect 16776 32524 20260 32552
rect 14550 32444 14556 32496
rect 14608 32444 14614 32496
rect 16022 32484 16028 32496
rect 15778 32456 16028 32484
rect 16022 32444 16028 32456
rect 16080 32484 16086 32496
rect 16390 32484 16396 32496
rect 16080 32456 16396 32484
rect 16080 32444 16086 32456
rect 16390 32444 16396 32456
rect 16448 32444 16454 32496
rect 12667 32388 14228 32416
rect 14277 32419 14335 32425
rect 12667 32385 12679 32388
rect 12621 32379 12679 32385
rect 14277 32385 14289 32419
rect 14323 32385 14335 32419
rect 14277 32379 14335 32385
rect 13357 32351 13415 32357
rect 13357 32317 13369 32351
rect 13403 32317 13415 32351
rect 13357 32311 13415 32317
rect 13541 32351 13599 32357
rect 13541 32317 13553 32351
rect 13587 32348 13599 32351
rect 13722 32348 13728 32360
rect 13587 32320 13728 32348
rect 13587 32317 13599 32320
rect 13541 32311 13599 32317
rect 13372 32280 13400 32311
rect 13722 32308 13728 32320
rect 13780 32308 13786 32360
rect 14292 32348 14320 32379
rect 15286 32348 15292 32360
rect 14292 32320 15292 32348
rect 15286 32308 15292 32320
rect 15344 32308 15350 32360
rect 16776 32280 16804 32524
rect 20254 32512 20260 32524
rect 20312 32512 20318 32564
rect 20990 32512 20996 32564
rect 21048 32512 21054 32564
rect 21726 32512 21732 32564
rect 21784 32552 21790 32564
rect 22005 32555 22063 32561
rect 22005 32552 22017 32555
rect 21784 32524 22017 32552
rect 21784 32512 21790 32524
rect 22005 32521 22017 32524
rect 22051 32521 22063 32555
rect 22005 32515 22063 32521
rect 22465 32555 22523 32561
rect 22465 32521 22477 32555
rect 22511 32552 22523 32555
rect 22830 32552 22836 32564
rect 22511 32524 22836 32552
rect 22511 32521 22523 32524
rect 22465 32515 22523 32521
rect 22830 32512 22836 32524
rect 22888 32512 22894 32564
rect 26252 32524 29868 32552
rect 17678 32444 17684 32496
rect 17736 32484 17742 32496
rect 19521 32487 19579 32493
rect 19521 32484 19533 32487
rect 17736 32456 19533 32484
rect 17736 32444 17742 32456
rect 19521 32453 19533 32456
rect 19567 32484 19579 32487
rect 19794 32484 19800 32496
rect 19567 32456 19800 32484
rect 19567 32453 19579 32456
rect 19521 32447 19579 32453
rect 19794 32444 19800 32456
rect 19852 32444 19858 32496
rect 20070 32444 20076 32496
rect 20128 32444 20134 32496
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 23842 32484 23848 32496
rect 22336 32456 22876 32484
rect 22336 32444 22342 32456
rect 22848 32428 22876 32456
rect 23584 32456 23848 32484
rect 17310 32376 17316 32428
rect 17368 32416 17374 32428
rect 17405 32419 17463 32425
rect 17405 32416 17417 32419
rect 17368 32388 17417 32416
rect 17368 32376 17374 32388
rect 17405 32385 17417 32388
rect 17451 32385 17463 32419
rect 17405 32379 17463 32385
rect 19058 32376 19064 32428
rect 19116 32416 19122 32428
rect 19245 32419 19303 32425
rect 19245 32416 19257 32419
rect 19116 32388 19257 32416
rect 19116 32376 19122 32388
rect 19245 32385 19257 32388
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 22186 32376 22192 32428
rect 22244 32416 22250 32428
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 22244 32388 22385 32416
rect 22244 32376 22250 32388
rect 22373 32385 22385 32388
rect 22419 32385 22431 32419
rect 22373 32379 22431 32385
rect 22480 32388 22692 32416
rect 17494 32308 17500 32360
rect 17552 32308 17558 32360
rect 17678 32308 17684 32360
rect 17736 32308 17742 32360
rect 18046 32308 18052 32360
rect 18104 32348 18110 32360
rect 22480 32348 22508 32388
rect 18104 32320 22508 32348
rect 18104 32308 18110 32320
rect 22554 32308 22560 32360
rect 22612 32308 22618 32360
rect 22664 32348 22692 32388
rect 22830 32376 22836 32428
rect 22888 32376 22894 32428
rect 23584 32348 23612 32456
rect 23842 32444 23848 32456
rect 23900 32444 23906 32496
rect 23934 32444 23940 32496
rect 23992 32444 23998 32496
rect 24394 32444 24400 32496
rect 24452 32444 24458 32496
rect 22664 32320 23612 32348
rect 23661 32351 23719 32357
rect 23661 32317 23673 32351
rect 23707 32317 23719 32351
rect 26252 32348 26280 32524
rect 28534 32444 28540 32496
rect 28592 32444 28598 32496
rect 29840 32484 29868 32524
rect 30558 32512 30564 32564
rect 30616 32552 30622 32564
rect 30929 32555 30987 32561
rect 30929 32552 30941 32555
rect 30616 32524 30941 32552
rect 30616 32512 30622 32524
rect 30929 32521 30941 32524
rect 30975 32521 30987 32555
rect 30929 32515 30987 32521
rect 32309 32555 32367 32561
rect 32309 32521 32321 32555
rect 32355 32552 32367 32555
rect 33594 32552 33600 32564
rect 32355 32524 33600 32552
rect 32355 32521 32367 32524
rect 32309 32515 32367 32521
rect 33594 32512 33600 32524
rect 33652 32512 33658 32564
rect 35434 32512 35440 32564
rect 35492 32552 35498 32564
rect 36633 32555 36691 32561
rect 36633 32552 36645 32555
rect 35492 32524 36645 32552
rect 35492 32512 35498 32524
rect 36633 32521 36645 32524
rect 36679 32521 36691 32555
rect 36633 32515 36691 32521
rect 31294 32484 31300 32496
rect 29840 32456 31300 32484
rect 31294 32444 31300 32456
rect 31352 32444 31358 32496
rect 31662 32444 31668 32496
rect 31720 32484 31726 32496
rect 31720 32456 34100 32484
rect 31720 32444 31726 32456
rect 30466 32416 30472 32428
rect 29670 32388 30472 32416
rect 30466 32376 30472 32388
rect 30524 32376 30530 32428
rect 30834 32376 30840 32428
rect 30892 32376 30898 32428
rect 32674 32376 32680 32428
rect 32732 32376 32738 32428
rect 32858 32376 32864 32428
rect 32916 32416 32922 32428
rect 32916 32388 33088 32416
rect 32916 32376 32922 32388
rect 23661 32311 23719 32317
rect 23768 32320 26280 32348
rect 28261 32351 28319 32357
rect 13372 32252 14228 32280
rect 1912 32184 2774 32212
rect 1912 32172 1918 32184
rect 12710 32172 12716 32224
rect 12768 32172 12774 32224
rect 14200 32221 14228 32252
rect 15948 32252 16804 32280
rect 14185 32215 14243 32221
rect 14185 32181 14197 32215
rect 14231 32212 14243 32215
rect 15948 32212 15976 32252
rect 17310 32240 17316 32292
rect 17368 32280 17374 32292
rect 19058 32280 19064 32292
rect 17368 32252 19064 32280
rect 17368 32240 17374 32252
rect 19058 32240 19064 32252
rect 19116 32240 19122 32292
rect 22278 32240 22284 32292
rect 22336 32280 22342 32292
rect 23676 32280 23704 32311
rect 22336 32252 23704 32280
rect 22336 32240 22342 32252
rect 14231 32184 15976 32212
rect 14231 32181 14243 32184
rect 14185 32175 14243 32181
rect 16022 32172 16028 32224
rect 16080 32172 16086 32224
rect 17037 32215 17095 32221
rect 17037 32181 17049 32215
rect 17083 32212 17095 32215
rect 19702 32212 19708 32224
rect 17083 32184 19708 32212
rect 17083 32181 17095 32184
rect 17037 32175 17095 32181
rect 19702 32172 19708 32184
rect 19760 32172 19766 32224
rect 20714 32172 20720 32224
rect 20772 32212 20778 32224
rect 21542 32212 21548 32224
rect 20772 32184 21548 32212
rect 20772 32172 20778 32184
rect 21542 32172 21548 32184
rect 21600 32212 21606 32224
rect 23768 32212 23796 32320
rect 28261 32317 28273 32351
rect 28307 32348 28319 32351
rect 29086 32348 29092 32360
rect 28307 32320 29092 32348
rect 28307 32317 28319 32320
rect 28261 32311 28319 32317
rect 29086 32308 29092 32320
rect 29144 32308 29150 32360
rect 29270 32308 29276 32360
rect 29328 32348 29334 32360
rect 30009 32351 30067 32357
rect 30009 32348 30021 32351
rect 29328 32320 30021 32348
rect 29328 32308 29334 32320
rect 30009 32317 30021 32320
rect 30055 32317 30067 32351
rect 30009 32311 30067 32317
rect 30374 32308 30380 32360
rect 30432 32348 30438 32360
rect 31021 32351 31079 32357
rect 31021 32348 31033 32351
rect 30432 32320 31033 32348
rect 30432 32308 30438 32320
rect 31021 32317 31033 32320
rect 31067 32317 31079 32351
rect 31021 32311 31079 32317
rect 32766 32308 32772 32360
rect 32824 32308 32830 32360
rect 32953 32351 33011 32357
rect 32953 32317 32965 32351
rect 32999 32317 33011 32351
rect 33060 32348 33088 32388
rect 33318 32376 33324 32428
rect 33376 32416 33382 32428
rect 33778 32416 33784 32428
rect 33376 32388 33784 32416
rect 33376 32376 33382 32388
rect 33778 32376 33784 32388
rect 33836 32376 33842 32428
rect 33870 32376 33876 32428
rect 33928 32376 33934 32428
rect 34072 32357 34100 32456
rect 36538 32376 36544 32428
rect 36596 32376 36602 32428
rect 33965 32351 34023 32357
rect 33965 32348 33977 32351
rect 33060 32320 33977 32348
rect 32953 32311 33011 32317
rect 33965 32317 33977 32320
rect 34011 32317 34023 32351
rect 33965 32311 34023 32317
rect 34057 32351 34115 32357
rect 34057 32317 34069 32351
rect 34103 32317 34115 32351
rect 34057 32311 34115 32317
rect 30469 32283 30527 32289
rect 30469 32249 30481 32283
rect 30515 32280 30527 32283
rect 32030 32280 32036 32292
rect 30515 32252 32036 32280
rect 30515 32249 30527 32252
rect 30469 32243 30527 32249
rect 32030 32240 32036 32252
rect 32088 32240 32094 32292
rect 21600 32184 23796 32212
rect 21600 32172 21606 32184
rect 23934 32172 23940 32224
rect 23992 32212 23998 32224
rect 25409 32215 25467 32221
rect 25409 32212 25421 32215
rect 23992 32184 25421 32212
rect 23992 32172 23998 32184
rect 25409 32181 25421 32184
rect 25455 32181 25467 32215
rect 25409 32175 25467 32181
rect 28534 32172 28540 32224
rect 28592 32212 28598 32224
rect 28718 32212 28724 32224
rect 28592 32184 28724 32212
rect 28592 32172 28598 32184
rect 28718 32172 28724 32184
rect 28776 32172 28782 32224
rect 30098 32172 30104 32224
rect 30156 32212 30162 32224
rect 31938 32212 31944 32224
rect 30156 32184 31944 32212
rect 30156 32172 30162 32184
rect 31938 32172 31944 32184
rect 31996 32172 32002 32224
rect 32968 32212 32996 32311
rect 36722 32308 36728 32360
rect 36780 32308 36786 32360
rect 33505 32283 33563 32289
rect 33505 32249 33517 32283
rect 33551 32280 33563 32283
rect 37826 32280 37832 32292
rect 33551 32252 37832 32280
rect 33551 32249 33563 32252
rect 33505 32243 33563 32249
rect 37826 32240 37832 32252
rect 37884 32240 37890 32292
rect 34238 32212 34244 32224
rect 32968 32184 34244 32212
rect 34238 32172 34244 32184
rect 34296 32172 34302 32224
rect 34606 32172 34612 32224
rect 34664 32212 34670 32224
rect 36173 32215 36231 32221
rect 36173 32212 36185 32215
rect 34664 32184 36185 32212
rect 34664 32172 34670 32184
rect 36173 32181 36185 32184
rect 36219 32181 36231 32215
rect 36173 32175 36231 32181
rect 1104 32122 49864 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 32950 32122
rect 33002 32070 33014 32122
rect 33066 32070 33078 32122
rect 33130 32070 33142 32122
rect 33194 32070 33206 32122
rect 33258 32070 42950 32122
rect 43002 32070 43014 32122
rect 43066 32070 43078 32122
rect 43130 32070 43142 32122
rect 43194 32070 43206 32122
rect 43258 32070 49864 32122
rect 1104 32048 49864 32070
rect 14752 31980 16528 32008
rect 12710 31940 12716 31952
rect 2746 31912 12716 31940
rect 1302 31832 1308 31884
rect 1360 31872 1366 31884
rect 2041 31875 2099 31881
rect 2041 31872 2053 31875
rect 1360 31844 2053 31872
rect 1360 31832 1366 31844
rect 2041 31841 2053 31844
rect 2087 31841 2099 31875
rect 2041 31835 2099 31841
rect 1765 31807 1823 31813
rect 1765 31773 1777 31807
rect 1811 31804 1823 31807
rect 2746 31804 2774 31912
rect 12710 31900 12716 31912
rect 12768 31900 12774 31952
rect 13630 31872 13636 31884
rect 8128 31844 13636 31872
rect 1811 31776 2774 31804
rect 1811 31773 1823 31776
rect 1765 31767 1823 31773
rect 7374 31764 7380 31816
rect 7432 31804 7438 31816
rect 8021 31807 8079 31813
rect 8021 31804 8033 31807
rect 7432 31776 8033 31804
rect 7432 31764 7438 31776
rect 8021 31773 8033 31776
rect 8067 31773 8079 31807
rect 8021 31767 8079 31773
rect 7837 31739 7895 31745
rect 7837 31705 7849 31739
rect 7883 31736 7895 31739
rect 8128 31736 8156 31844
rect 13630 31832 13636 31844
rect 13688 31832 13694 31884
rect 10965 31807 11023 31813
rect 10965 31773 10977 31807
rect 11011 31804 11023 31807
rect 14752 31804 14780 31980
rect 16500 31940 16528 31980
rect 16574 31968 16580 32020
rect 16632 31968 16638 32020
rect 17310 32008 17316 32020
rect 17144 31980 17316 32008
rect 17144 31940 17172 31980
rect 17310 31968 17316 31980
rect 17368 31968 17374 32020
rect 17494 31968 17500 32020
rect 17552 32008 17558 32020
rect 18046 32008 18052 32020
rect 17552 31980 18052 32008
rect 17552 31968 17558 31980
rect 18046 31968 18052 31980
rect 18104 31968 18110 32020
rect 18782 31968 18788 32020
rect 18840 31968 18846 32020
rect 19426 31968 19432 32020
rect 19484 32008 19490 32020
rect 21085 32011 21143 32017
rect 21085 32008 21097 32011
rect 19484 31980 21097 32008
rect 19484 31968 19490 31980
rect 21085 31977 21097 31980
rect 21131 31977 21143 32011
rect 21085 31971 21143 31977
rect 22646 31968 22652 32020
rect 22704 32008 22710 32020
rect 23658 32008 23664 32020
rect 22704 31980 23664 32008
rect 22704 31968 22710 31980
rect 23658 31968 23664 31980
rect 23716 31968 23722 32020
rect 24026 31968 24032 32020
rect 24084 31968 24090 32020
rect 28261 32011 28319 32017
rect 28261 31977 28273 32011
rect 28307 32008 28319 32011
rect 30098 32008 30104 32020
rect 28307 31980 30104 32008
rect 28307 31977 28319 31980
rect 28261 31971 28319 31977
rect 30098 31968 30104 31980
rect 30156 31968 30162 32020
rect 31846 32008 31852 32020
rect 31036 31980 31852 32008
rect 16500 31912 17172 31940
rect 19058 31900 19064 31952
rect 19116 31940 19122 31952
rect 20714 31940 20720 31952
rect 19116 31912 20720 31940
rect 19116 31900 19122 31912
rect 20714 31900 20720 31912
rect 20772 31900 20778 31952
rect 21450 31940 21456 31952
rect 21192 31912 21456 31940
rect 14829 31875 14887 31881
rect 14829 31841 14841 31875
rect 14875 31872 14887 31875
rect 15194 31872 15200 31884
rect 14875 31844 15200 31872
rect 14875 31841 14887 31844
rect 14829 31835 14887 31841
rect 15194 31832 15200 31844
rect 15252 31872 15258 31884
rect 17313 31875 17371 31881
rect 15252 31844 16344 31872
rect 15252 31832 15258 31844
rect 11011 31776 14780 31804
rect 16316 31804 16344 31844
rect 17313 31841 17325 31875
rect 17359 31872 17371 31875
rect 17359 31844 19196 31872
rect 17359 31841 17371 31844
rect 17313 31835 17371 31841
rect 17037 31807 17095 31813
rect 17037 31804 17049 31807
rect 16316 31776 17049 31804
rect 11011 31773 11023 31776
rect 10965 31767 11023 31773
rect 17037 31773 17049 31776
rect 17083 31773 17095 31807
rect 19168 31804 19196 31844
rect 19242 31832 19248 31884
rect 19300 31872 19306 31884
rect 20257 31875 20315 31881
rect 20257 31872 20269 31875
rect 19300 31844 20269 31872
rect 19300 31832 19306 31844
rect 20257 31841 20269 31844
rect 20303 31841 20315 31875
rect 20257 31835 20315 31841
rect 20441 31875 20499 31881
rect 20441 31841 20453 31875
rect 20487 31872 20499 31875
rect 21192 31872 21220 31912
rect 21450 31900 21456 31912
rect 21508 31900 21514 31952
rect 25869 31943 25927 31949
rect 25869 31909 25881 31943
rect 25915 31940 25927 31943
rect 29454 31940 29460 31952
rect 25915 31912 28672 31940
rect 25915 31909 25927 31912
rect 25869 31903 25927 31909
rect 20487 31844 21220 31872
rect 20487 31841 20499 31844
rect 20441 31835 20499 31841
rect 21358 31832 21364 31884
rect 21416 31832 21422 31884
rect 21634 31832 21640 31884
rect 21692 31832 21698 31884
rect 22278 31872 22284 31884
rect 22066 31844 22284 31872
rect 19610 31804 19616 31816
rect 19168 31776 19616 31804
rect 17037 31767 17095 31773
rect 19610 31764 19616 31776
rect 19668 31804 19674 31816
rect 19668 31776 20300 31804
rect 19668 31764 19674 31776
rect 7883 31708 8156 31736
rect 15105 31739 15163 31745
rect 7883 31705 7895 31708
rect 7837 31699 7895 31705
rect 15105 31705 15117 31739
rect 15151 31736 15163 31739
rect 16390 31736 16396 31748
rect 15151 31708 15516 31736
rect 16330 31708 16396 31736
rect 15151 31705 15163 31708
rect 15105 31699 15163 31705
rect 11054 31628 11060 31680
rect 11112 31628 11118 31680
rect 15488 31668 15516 31708
rect 16390 31696 16396 31708
rect 16448 31736 16454 31748
rect 16850 31736 16856 31748
rect 16448 31708 16856 31736
rect 16448 31696 16454 31708
rect 16850 31696 16856 31708
rect 16908 31696 16914 31748
rect 19058 31736 19064 31748
rect 18538 31708 19064 31736
rect 19058 31696 19064 31708
rect 19116 31736 19122 31748
rect 20070 31736 20076 31748
rect 19116 31708 20076 31736
rect 19116 31696 19122 31708
rect 20070 31696 20076 31708
rect 20128 31696 20134 31748
rect 20162 31696 20168 31748
rect 20220 31696 20226 31748
rect 20272 31736 20300 31776
rect 20806 31764 20812 31816
rect 20864 31804 20870 31816
rect 21376 31804 21404 31832
rect 22066 31804 22094 31844
rect 22278 31832 22284 31844
rect 22336 31832 22342 31884
rect 22557 31875 22615 31881
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23934 31872 23940 31884
rect 22603 31844 23940 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23934 31832 23940 31844
rect 23992 31832 23998 31884
rect 26326 31832 26332 31884
rect 26384 31832 26390 31884
rect 26513 31875 26571 31881
rect 26513 31841 26525 31875
rect 26559 31872 26571 31875
rect 26970 31872 26976 31884
rect 26559 31844 26976 31872
rect 26559 31841 26571 31844
rect 26513 31835 26571 31841
rect 26970 31832 26976 31844
rect 27028 31832 27034 31884
rect 20864 31776 22094 31804
rect 20864 31764 20870 31776
rect 27798 31764 27804 31816
rect 27856 31764 27862 31816
rect 21082 31736 21088 31748
rect 20272 31708 21088 31736
rect 21082 31696 21088 31708
rect 21140 31696 21146 31748
rect 21545 31739 21603 31745
rect 21545 31736 21557 31739
rect 21376 31708 21557 31736
rect 21376 31680 21404 31708
rect 21545 31705 21557 31708
rect 21591 31705 21603 31739
rect 21545 31699 21603 31705
rect 22002 31696 22008 31748
rect 22060 31736 22066 31748
rect 28644 31736 28672 31912
rect 28828 31912 29460 31940
rect 28718 31832 28724 31884
rect 28776 31832 28782 31884
rect 28828 31804 28856 31912
rect 29454 31900 29460 31912
rect 29512 31900 29518 31952
rect 28902 31832 28908 31884
rect 28960 31832 28966 31884
rect 29086 31832 29092 31884
rect 29144 31872 29150 31884
rect 29730 31872 29736 31884
rect 29144 31844 29736 31872
rect 29144 31832 29150 31844
rect 29730 31832 29736 31844
rect 29788 31832 29794 31884
rect 30006 31832 30012 31884
rect 30064 31872 30070 31884
rect 31036 31872 31064 31980
rect 31846 31968 31852 31980
rect 31904 31968 31910 32020
rect 31941 32011 31999 32017
rect 31941 31977 31953 32011
rect 31987 32008 31999 32011
rect 33137 32011 33195 32017
rect 31987 31980 33088 32008
rect 31987 31977 31999 31980
rect 31941 31971 31999 31977
rect 31110 31900 31116 31952
rect 31168 31940 31174 31952
rect 31481 31943 31539 31949
rect 31481 31940 31493 31943
rect 31168 31912 31493 31940
rect 31168 31900 31174 31912
rect 31481 31909 31493 31912
rect 31527 31909 31539 31943
rect 31481 31903 31539 31909
rect 32122 31900 32128 31952
rect 32180 31940 32186 31952
rect 33060 31940 33088 31980
rect 33137 31977 33149 32011
rect 33183 32008 33195 32011
rect 33410 32008 33416 32020
rect 33183 31980 33416 32008
rect 33183 31977 33195 31980
rect 33137 31971 33195 31977
rect 33410 31968 33416 31980
rect 33468 31968 33474 32020
rect 33778 32008 33784 32020
rect 33520 31980 33784 32008
rect 33520 31940 33548 31980
rect 33778 31968 33784 31980
rect 33836 31968 33842 32020
rect 49237 31943 49295 31949
rect 49237 31940 49249 31943
rect 32180 31912 32536 31940
rect 33060 31912 33548 31940
rect 33612 31912 41414 31940
rect 32180 31900 32186 31912
rect 31202 31872 31208 31884
rect 30064 31844 31064 31872
rect 31128 31844 31208 31872
rect 30064 31832 30070 31844
rect 28828 31776 28948 31804
rect 28920 31736 28948 31776
rect 28994 31764 29000 31816
rect 29052 31804 29058 31816
rect 29052 31776 29776 31804
rect 31128 31790 31156 31844
rect 31202 31832 31208 31844
rect 31260 31832 31266 31884
rect 31386 31832 31392 31884
rect 31444 31872 31450 31884
rect 32508 31881 32536 31912
rect 32401 31875 32459 31881
rect 32401 31872 32413 31875
rect 31444 31844 32413 31872
rect 31444 31832 31450 31844
rect 32401 31841 32413 31844
rect 32447 31841 32459 31875
rect 32401 31835 32459 31841
rect 32493 31875 32551 31881
rect 32493 31841 32505 31875
rect 32539 31841 32551 31875
rect 33612 31872 33640 31912
rect 32493 31835 32551 31841
rect 33520 31844 33640 31872
rect 29052 31764 29058 31776
rect 22060 31708 23046 31736
rect 28644 31708 28948 31736
rect 29748 31736 29776 31776
rect 31294 31764 31300 31816
rect 31352 31804 31358 31816
rect 33520 31804 33548 31844
rect 33686 31832 33692 31884
rect 33744 31832 33750 31884
rect 41386 31872 41414 31912
rect 45526 31912 49249 31940
rect 45526 31872 45554 31912
rect 49237 31909 49249 31912
rect 49283 31909 49295 31943
rect 49237 31903 49295 31909
rect 41386 31844 45554 31872
rect 31352 31776 33548 31804
rect 31352 31764 31358 31776
rect 33594 31764 33600 31816
rect 33652 31764 33658 31816
rect 49050 31764 49056 31816
rect 49108 31764 49114 31816
rect 30006 31736 30012 31748
rect 29748 31708 30012 31736
rect 22060 31696 22066 31708
rect 30006 31696 30012 31708
rect 30064 31696 30070 31748
rect 33502 31696 33508 31748
rect 33560 31696 33566 31748
rect 16482 31668 16488 31680
rect 15488 31640 16488 31668
rect 16482 31628 16488 31640
rect 16540 31668 16546 31680
rect 19518 31668 19524 31680
rect 16540 31640 19524 31668
rect 16540 31628 16546 31640
rect 19518 31628 19524 31640
rect 19576 31628 19582 31680
rect 19794 31628 19800 31680
rect 19852 31628 19858 31680
rect 21358 31628 21364 31680
rect 21416 31628 21422 31680
rect 21453 31671 21511 31677
rect 21453 31637 21465 31671
rect 21499 31668 21511 31671
rect 21634 31668 21640 31680
rect 21499 31640 21640 31668
rect 21499 31637 21511 31640
rect 21453 31631 21511 31637
rect 21634 31628 21640 31640
rect 21692 31628 21698 31680
rect 22186 31628 22192 31680
rect 22244 31668 22250 31680
rect 26237 31671 26295 31677
rect 26237 31668 26249 31671
rect 22244 31640 26249 31668
rect 22244 31628 22250 31640
rect 26237 31637 26249 31640
rect 26283 31637 26295 31671
rect 26237 31631 26295 31637
rect 28629 31671 28687 31677
rect 28629 31637 28641 31671
rect 28675 31668 28687 31671
rect 28718 31668 28724 31680
rect 28675 31640 28724 31668
rect 28675 31637 28687 31640
rect 28629 31631 28687 31637
rect 28718 31628 28724 31640
rect 28776 31628 28782 31680
rect 32306 31628 32312 31680
rect 32364 31628 32370 31680
rect 1104 31578 49864 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 27950 31578
rect 28002 31526 28014 31578
rect 28066 31526 28078 31578
rect 28130 31526 28142 31578
rect 28194 31526 28206 31578
rect 28258 31526 37950 31578
rect 38002 31526 38014 31578
rect 38066 31526 38078 31578
rect 38130 31526 38142 31578
rect 38194 31526 38206 31578
rect 38258 31526 47950 31578
rect 48002 31526 48014 31578
rect 48066 31526 48078 31578
rect 48130 31526 48142 31578
rect 48194 31526 48206 31578
rect 48258 31526 49864 31578
rect 1104 31504 49864 31526
rect 13173 31467 13231 31473
rect 13173 31433 13185 31467
rect 13219 31433 13231 31467
rect 13173 31427 13231 31433
rect 11054 31396 11060 31408
rect 6886 31368 11060 31396
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31328 1823 31331
rect 6886 31328 6914 31368
rect 11054 31356 11060 31368
rect 11112 31356 11118 31408
rect 13188 31396 13216 31427
rect 13538 31424 13544 31476
rect 13596 31424 13602 31476
rect 13630 31424 13636 31476
rect 13688 31424 13694 31476
rect 14734 31424 14740 31476
rect 14792 31424 14798 31476
rect 15654 31424 15660 31476
rect 15712 31464 15718 31476
rect 15933 31467 15991 31473
rect 15933 31464 15945 31467
rect 15712 31436 15945 31464
rect 15712 31424 15718 31436
rect 15933 31433 15945 31436
rect 15979 31433 15991 31467
rect 15933 31427 15991 31433
rect 16025 31467 16083 31473
rect 16025 31433 16037 31467
rect 16071 31464 16083 31467
rect 17218 31464 17224 31476
rect 16071 31436 17224 31464
rect 16071 31433 16083 31436
rect 16025 31427 16083 31433
rect 17218 31424 17224 31436
rect 17276 31424 17282 31476
rect 17402 31424 17408 31476
rect 17460 31424 17466 31476
rect 20806 31464 20812 31476
rect 18248 31436 20812 31464
rect 15746 31396 15752 31408
rect 13188 31368 15752 31396
rect 15746 31356 15752 31368
rect 15804 31356 15810 31408
rect 16114 31356 16120 31408
rect 16172 31396 16178 31408
rect 17497 31399 17555 31405
rect 17497 31396 17509 31399
rect 16172 31368 17509 31396
rect 16172 31356 16178 31368
rect 17497 31365 17509 31368
rect 17543 31365 17555 31399
rect 17497 31359 17555 31365
rect 1811 31300 6914 31328
rect 1811 31297 1823 31300
rect 1765 31291 1823 31297
rect 10686 31288 10692 31340
rect 10744 31288 10750 31340
rect 15470 31328 15476 31340
rect 14844 31300 15476 31328
rect 1302 31220 1308 31272
rect 1360 31260 1366 31272
rect 2041 31263 2099 31269
rect 2041 31260 2053 31263
rect 1360 31232 2053 31260
rect 1360 31220 1366 31232
rect 2041 31229 2053 31232
rect 2087 31229 2099 31263
rect 2041 31223 2099 31229
rect 12526 31220 12532 31272
rect 12584 31260 12590 31272
rect 13722 31260 13728 31272
rect 12584 31232 13728 31260
rect 12584 31220 12590 31232
rect 13722 31220 13728 31232
rect 13780 31220 13786 31272
rect 14734 31220 14740 31272
rect 14792 31260 14798 31272
rect 14844 31269 14872 31300
rect 15470 31288 15476 31300
rect 15528 31288 15534 31340
rect 18248 31337 18276 31436
rect 20806 31424 20812 31436
rect 20864 31424 20870 31476
rect 27617 31467 27675 31473
rect 27617 31433 27629 31467
rect 27663 31464 27675 31467
rect 27798 31464 27804 31476
rect 27663 31436 27804 31464
rect 27663 31433 27675 31436
rect 27617 31427 27675 31433
rect 27798 31424 27804 31436
rect 27856 31424 27862 31476
rect 29178 31424 29184 31476
rect 29236 31464 29242 31476
rect 29549 31467 29607 31473
rect 29549 31464 29561 31467
rect 29236 31436 29561 31464
rect 29236 31424 29242 31436
rect 29549 31433 29561 31436
rect 29595 31433 29607 31467
rect 29549 31427 29607 31433
rect 19058 31356 19064 31408
rect 19116 31356 19122 31408
rect 20898 31396 20904 31408
rect 20824 31368 20904 31396
rect 20824 31337 20852 31368
rect 20898 31356 20904 31368
rect 20956 31356 20962 31408
rect 21634 31356 21640 31408
rect 21692 31396 21698 31408
rect 31478 31396 31484 31408
rect 21692 31368 31484 31396
rect 21692 31356 21698 31368
rect 31478 31356 31484 31368
rect 31536 31356 31542 31408
rect 33594 31396 33600 31408
rect 31726 31368 33600 31396
rect 18233 31331 18291 31337
rect 18233 31297 18245 31331
rect 18279 31297 18291 31331
rect 18233 31291 18291 31297
rect 20809 31331 20867 31337
rect 20809 31297 20821 31331
rect 20855 31297 20867 31331
rect 20809 31291 20867 31297
rect 21266 31288 21272 31340
rect 21324 31328 21330 31340
rect 28629 31331 28687 31337
rect 28629 31328 28641 31331
rect 21324 31300 28641 31328
rect 21324 31288 21330 31300
rect 28629 31297 28641 31300
rect 28675 31328 28687 31331
rect 29641 31331 29699 31337
rect 29641 31328 29653 31331
rect 28675 31300 29653 31328
rect 28675 31297 28687 31300
rect 28629 31291 28687 31297
rect 29641 31297 29653 31300
rect 29687 31328 29699 31331
rect 31726 31328 31754 31368
rect 33594 31356 33600 31368
rect 33652 31356 33658 31408
rect 39942 31356 39948 31408
rect 40000 31396 40006 31408
rect 44453 31399 44511 31405
rect 44453 31396 44465 31399
rect 40000 31368 44465 31396
rect 40000 31356 40006 31368
rect 44453 31365 44465 31368
rect 44499 31365 44511 31399
rect 44453 31359 44511 31365
rect 29687 31300 31754 31328
rect 32493 31331 32551 31337
rect 29687 31297 29699 31300
rect 29641 31291 29699 31297
rect 32493 31297 32505 31331
rect 32539 31328 32551 31331
rect 32674 31328 32680 31340
rect 32539 31300 32680 31328
rect 32539 31297 32551 31300
rect 32493 31291 32551 31297
rect 32674 31288 32680 31300
rect 32732 31288 32738 31340
rect 37182 31288 37188 31340
rect 37240 31328 37246 31340
rect 38381 31331 38439 31337
rect 38381 31328 38393 31331
rect 37240 31300 38393 31328
rect 37240 31288 37246 31300
rect 38381 31297 38393 31300
rect 38427 31297 38439 31331
rect 38381 31291 38439 31297
rect 49326 31288 49332 31340
rect 49384 31288 49390 31340
rect 14829 31263 14887 31269
rect 14829 31260 14841 31263
rect 14792 31232 14841 31260
rect 14792 31220 14798 31232
rect 14829 31229 14841 31232
rect 14875 31229 14887 31263
rect 14829 31223 14887 31229
rect 15013 31263 15071 31269
rect 15013 31229 15025 31263
rect 15059 31260 15071 31263
rect 15838 31260 15844 31272
rect 15059 31232 15844 31260
rect 15059 31229 15071 31232
rect 15013 31223 15071 31229
rect 15838 31220 15844 31232
rect 15896 31260 15902 31272
rect 15896 31232 16160 31260
rect 15896 31220 15902 31232
rect 14369 31195 14427 31201
rect 14369 31161 14381 31195
rect 14415 31192 14427 31195
rect 16022 31192 16028 31204
rect 14415 31164 16028 31192
rect 14415 31161 14427 31164
rect 14369 31155 14427 31161
rect 16022 31152 16028 31164
rect 16080 31152 16086 31204
rect 16132 31192 16160 31232
rect 16206 31220 16212 31272
rect 16264 31220 16270 31272
rect 17402 31220 17408 31272
rect 17460 31260 17466 31272
rect 17589 31263 17647 31269
rect 17589 31260 17601 31263
rect 17460 31232 17601 31260
rect 17460 31220 17466 31232
rect 17589 31229 17601 31232
rect 17635 31229 17647 31263
rect 17589 31223 17647 31229
rect 18509 31263 18567 31269
rect 18509 31229 18521 31263
rect 18555 31260 18567 31263
rect 18555 31232 20300 31260
rect 18555 31229 18567 31232
rect 18509 31223 18567 31229
rect 17862 31192 17868 31204
rect 16132 31164 17868 31192
rect 17862 31152 17868 31164
rect 17920 31152 17926 31204
rect 19518 31152 19524 31204
rect 19576 31192 19582 31204
rect 19981 31195 20039 31201
rect 19981 31192 19993 31195
rect 19576 31164 19993 31192
rect 19576 31152 19582 31164
rect 19981 31161 19993 31164
rect 20027 31161 20039 31195
rect 20272 31192 20300 31232
rect 20898 31220 20904 31272
rect 20956 31220 20962 31272
rect 21082 31220 21088 31272
rect 21140 31260 21146 31272
rect 21910 31260 21916 31272
rect 21140 31232 21916 31260
rect 21140 31220 21146 31232
rect 21910 31220 21916 31232
rect 21968 31220 21974 31272
rect 22554 31220 22560 31272
rect 22612 31260 22618 31272
rect 26510 31260 26516 31272
rect 22612 31232 26516 31260
rect 22612 31220 22618 31232
rect 26510 31220 26516 31232
rect 26568 31220 26574 31272
rect 27614 31220 27620 31272
rect 27672 31260 27678 31272
rect 27709 31263 27767 31269
rect 27709 31260 27721 31263
rect 27672 31232 27721 31260
rect 27672 31220 27678 31232
rect 27709 31229 27721 31232
rect 27755 31229 27767 31263
rect 27709 31223 27767 31229
rect 27893 31263 27951 31269
rect 27893 31229 27905 31263
rect 27939 31260 27951 31263
rect 29270 31260 29276 31272
rect 27939 31232 29276 31260
rect 27939 31229 27951 31232
rect 27893 31223 27951 31229
rect 29270 31220 29276 31232
rect 29328 31220 29334 31272
rect 29822 31220 29828 31272
rect 29880 31220 29886 31272
rect 38562 31220 38568 31272
rect 38620 31260 38626 31272
rect 38620 31232 49188 31260
rect 38620 31220 38626 31232
rect 22370 31192 22376 31204
rect 20272 31164 22376 31192
rect 19981 31155 20039 31161
rect 22370 31152 22376 31164
rect 22428 31152 22434 31204
rect 25130 31192 25136 31204
rect 23308 31164 25136 31192
rect 8662 31084 8668 31136
rect 8720 31124 8726 31136
rect 10781 31127 10839 31133
rect 10781 31124 10793 31127
rect 8720 31096 10793 31124
rect 8720 31084 8726 31096
rect 10781 31093 10793 31096
rect 10827 31093 10839 31127
rect 10781 31087 10839 31093
rect 14826 31084 14832 31136
rect 14884 31124 14890 31136
rect 15565 31127 15623 31133
rect 15565 31124 15577 31127
rect 14884 31096 15577 31124
rect 14884 31084 14890 31096
rect 15565 31093 15577 31096
rect 15611 31093 15623 31127
rect 15565 31087 15623 31093
rect 15930 31084 15936 31136
rect 15988 31124 15994 31136
rect 16206 31124 16212 31136
rect 15988 31096 16212 31124
rect 15988 31084 15994 31096
rect 16206 31084 16212 31096
rect 16264 31084 16270 31136
rect 17037 31127 17095 31133
rect 17037 31093 17049 31127
rect 17083 31124 17095 31127
rect 18506 31124 18512 31136
rect 17083 31096 18512 31124
rect 17083 31093 17095 31096
rect 17037 31087 17095 31093
rect 18506 31084 18512 31096
rect 18564 31084 18570 31136
rect 20438 31084 20444 31136
rect 20496 31084 20502 31136
rect 20898 31084 20904 31136
rect 20956 31124 20962 31136
rect 21726 31124 21732 31136
rect 20956 31096 21732 31124
rect 20956 31084 20962 31096
rect 21726 31084 21732 31096
rect 21784 31124 21790 31136
rect 23308 31124 23336 31164
rect 25130 31152 25136 31164
rect 25188 31152 25194 31204
rect 27249 31195 27307 31201
rect 27249 31161 27261 31195
rect 27295 31192 27307 31195
rect 30834 31192 30840 31204
rect 27295 31164 30840 31192
rect 27295 31161 27307 31164
rect 27249 31155 27307 31161
rect 30834 31152 30840 31164
rect 30892 31152 30898 31204
rect 44637 31195 44695 31201
rect 44637 31161 44649 31195
rect 44683 31192 44695 31195
rect 46750 31192 46756 31204
rect 44683 31164 46756 31192
rect 44683 31161 44695 31164
rect 44637 31155 44695 31161
rect 46750 31152 46756 31164
rect 46808 31152 46814 31204
rect 49160 31201 49188 31232
rect 49145 31195 49203 31201
rect 49145 31161 49157 31195
rect 49191 31161 49203 31195
rect 49145 31155 49203 31161
rect 21784 31096 23336 31124
rect 21784 31084 21790 31096
rect 23382 31084 23388 31136
rect 23440 31084 23446 31136
rect 24397 31127 24455 31133
rect 24397 31093 24409 31127
rect 24443 31124 24455 31127
rect 24946 31124 24952 31136
rect 24443 31096 24952 31124
rect 24443 31093 24455 31096
rect 24397 31087 24455 31093
rect 24946 31084 24952 31096
rect 25004 31084 25010 31136
rect 29181 31127 29239 31133
rect 29181 31093 29193 31127
rect 29227 31124 29239 31127
rect 33870 31124 33876 31136
rect 29227 31096 33876 31124
rect 29227 31093 29239 31096
rect 29181 31087 29239 31093
rect 33870 31084 33876 31096
rect 33928 31084 33934 31136
rect 38197 31127 38255 31133
rect 38197 31093 38209 31127
rect 38243 31124 38255 31127
rect 44542 31124 44548 31136
rect 38243 31096 44548 31124
rect 38243 31093 38255 31096
rect 38197 31087 38255 31093
rect 44542 31084 44548 31096
rect 44600 31084 44606 31136
rect 1104 31034 49864 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 32950 31034
rect 33002 30982 33014 31034
rect 33066 30982 33078 31034
rect 33130 30982 33142 31034
rect 33194 30982 33206 31034
rect 33258 30982 42950 31034
rect 43002 30982 43014 31034
rect 43066 30982 43078 31034
rect 43130 30982 43142 31034
rect 43194 30982 43206 31034
rect 43258 30982 49864 31034
rect 1104 30960 49864 30982
rect 10686 30880 10692 30932
rect 10744 30920 10750 30932
rect 22554 30920 22560 30932
rect 10744 30892 19334 30920
rect 10744 30880 10750 30892
rect 19306 30864 19334 30892
rect 19444 30892 22560 30920
rect 19058 30852 19064 30864
rect 17236 30824 19064 30852
rect 14458 30744 14464 30796
rect 14516 30784 14522 30796
rect 14921 30787 14979 30793
rect 14921 30784 14933 30787
rect 14516 30756 14933 30784
rect 14516 30744 14522 30756
rect 14921 30753 14933 30756
rect 14967 30753 14979 30787
rect 14921 30747 14979 30753
rect 15010 30744 15016 30796
rect 15068 30744 15074 30796
rect 16666 30744 16672 30796
rect 16724 30784 16730 30796
rect 16850 30784 16856 30796
rect 16724 30756 16856 30784
rect 16724 30744 16730 30756
rect 16850 30744 16856 30756
rect 16908 30784 16914 30796
rect 17236 30784 17264 30824
rect 19058 30812 19064 30824
rect 19116 30812 19122 30864
rect 19306 30824 19340 30864
rect 19334 30812 19340 30824
rect 19392 30812 19398 30864
rect 16908 30756 17264 30784
rect 16908 30744 16914 30756
rect 11146 30676 11152 30728
rect 11204 30716 11210 30728
rect 13725 30719 13783 30725
rect 13725 30716 13737 30719
rect 11204 30688 13737 30716
rect 11204 30676 11210 30688
rect 13725 30685 13737 30688
rect 13771 30685 13783 30719
rect 13725 30679 13783 30685
rect 14826 30676 14832 30728
rect 14884 30676 14890 30728
rect 15194 30676 15200 30728
rect 15252 30716 15258 30728
rect 15841 30719 15899 30725
rect 15841 30716 15853 30719
rect 15252 30688 15853 30716
rect 15252 30676 15258 30688
rect 15841 30685 15853 30688
rect 15887 30685 15899 30719
rect 17236 30702 17264 30756
rect 17862 30744 17868 30796
rect 17920 30744 17926 30796
rect 19444 30784 19472 30892
rect 22554 30880 22560 30892
rect 22612 30880 22618 30932
rect 23290 30880 23296 30932
rect 23348 30920 23354 30932
rect 24581 30923 24639 30929
rect 24581 30920 24593 30923
rect 23348 30892 24593 30920
rect 23348 30880 23354 30892
rect 24581 30889 24593 30892
rect 24627 30889 24639 30923
rect 24581 30883 24639 30889
rect 26145 30923 26203 30929
rect 26145 30889 26157 30923
rect 26191 30920 26203 30923
rect 30190 30920 30196 30932
rect 26191 30892 30196 30920
rect 26191 30889 26203 30892
rect 26145 30883 26203 30889
rect 30190 30880 30196 30892
rect 30248 30880 30254 30932
rect 20162 30812 20168 30864
rect 20220 30852 20226 30864
rect 20220 30824 22094 30852
rect 20220 30812 20226 30824
rect 18708 30756 19472 30784
rect 15841 30679 15899 30685
rect 12802 30608 12808 30660
rect 12860 30608 12866 30660
rect 13541 30651 13599 30657
rect 13541 30617 13553 30651
rect 13587 30648 13599 30651
rect 16117 30651 16175 30657
rect 13587 30620 16068 30648
rect 13587 30617 13599 30620
rect 13541 30611 13599 30617
rect 11054 30540 11060 30592
rect 11112 30580 11118 30592
rect 12897 30583 12955 30589
rect 12897 30580 12909 30583
rect 11112 30552 12909 30580
rect 11112 30540 11118 30552
rect 12897 30549 12909 30552
rect 12943 30549 12955 30583
rect 12897 30543 12955 30549
rect 14461 30583 14519 30589
rect 14461 30549 14473 30583
rect 14507 30580 14519 30583
rect 15838 30580 15844 30592
rect 14507 30552 15844 30580
rect 14507 30549 14519 30552
rect 14461 30543 14519 30549
rect 15838 30540 15844 30552
rect 15896 30540 15902 30592
rect 16040 30580 16068 30620
rect 16117 30617 16129 30651
rect 16163 30648 16175 30651
rect 16390 30648 16396 30660
rect 16163 30620 16396 30648
rect 16163 30617 16175 30620
rect 16117 30611 16175 30617
rect 16390 30608 16396 30620
rect 16448 30608 16454 30660
rect 18708 30580 18736 30756
rect 20714 30744 20720 30796
rect 20772 30784 20778 30796
rect 20901 30787 20959 30793
rect 20901 30784 20913 30787
rect 20772 30756 20913 30784
rect 20772 30744 20778 30756
rect 20901 30753 20913 30756
rect 20947 30753 20959 30787
rect 20901 30747 20959 30753
rect 20993 30787 21051 30793
rect 20993 30753 21005 30787
rect 21039 30753 21051 30787
rect 22066 30784 22094 30824
rect 23492 30824 25176 30852
rect 23492 30784 23520 30824
rect 22066 30756 23520 30784
rect 20993 30747 21051 30753
rect 18782 30676 18788 30728
rect 18840 30716 18846 30728
rect 21008 30716 21036 30747
rect 23566 30744 23572 30796
rect 23624 30784 23630 30796
rect 23753 30787 23811 30793
rect 23753 30784 23765 30787
rect 23624 30756 23765 30784
rect 23624 30744 23630 30756
rect 23753 30753 23765 30756
rect 23799 30753 23811 30787
rect 23753 30747 23811 30753
rect 23934 30744 23940 30796
rect 23992 30744 23998 30796
rect 18840 30688 21036 30716
rect 18840 30676 18846 30688
rect 24946 30676 24952 30728
rect 25004 30676 25010 30728
rect 25148 30716 25176 30824
rect 25222 30744 25228 30796
rect 25280 30744 25286 30796
rect 26789 30787 26847 30793
rect 26789 30753 26801 30787
rect 26835 30784 26847 30787
rect 26878 30784 26884 30796
rect 26835 30756 26884 30784
rect 26835 30753 26847 30756
rect 26789 30747 26847 30753
rect 26878 30744 26884 30756
rect 26936 30744 26942 30796
rect 26513 30719 26571 30725
rect 26513 30716 26525 30719
rect 25148 30688 26525 30716
rect 26513 30685 26525 30688
rect 26559 30685 26571 30719
rect 26513 30679 26571 30685
rect 42610 30676 42616 30728
rect 42668 30716 42674 30728
rect 45281 30719 45339 30725
rect 45281 30716 45293 30719
rect 42668 30688 45293 30716
rect 42668 30676 42674 30688
rect 45281 30685 45293 30688
rect 45327 30685 45339 30719
rect 45281 30679 45339 30685
rect 20809 30651 20867 30657
rect 20809 30617 20821 30651
rect 20855 30648 20867 30651
rect 22186 30648 22192 30660
rect 20855 30620 22192 30648
rect 20855 30617 20867 30620
rect 20809 30611 20867 30617
rect 22186 30608 22192 30620
rect 22244 30608 22250 30660
rect 25041 30651 25099 30657
rect 25041 30617 25053 30651
rect 25087 30648 25099 30651
rect 28718 30648 28724 30660
rect 25087 30620 28724 30648
rect 25087 30617 25099 30620
rect 25041 30611 25099 30617
rect 28718 30608 28724 30620
rect 28776 30608 28782 30660
rect 45465 30651 45523 30657
rect 45465 30617 45477 30651
rect 45511 30648 45523 30651
rect 46474 30648 46480 30660
rect 45511 30620 46480 30648
rect 45511 30617 45523 30620
rect 45465 30611 45523 30617
rect 46474 30608 46480 30620
rect 46532 30608 46538 30660
rect 16040 30552 18736 30580
rect 18966 30540 18972 30592
rect 19024 30580 19030 30592
rect 20441 30583 20499 30589
rect 20441 30580 20453 30583
rect 19024 30552 20453 30580
rect 19024 30540 19030 30552
rect 20441 30549 20453 30552
rect 20487 30549 20499 30583
rect 20441 30543 20499 30549
rect 21174 30540 21180 30592
rect 21232 30580 21238 30592
rect 23293 30583 23351 30589
rect 23293 30580 23305 30583
rect 21232 30552 23305 30580
rect 21232 30540 21238 30552
rect 23293 30549 23305 30552
rect 23339 30549 23351 30583
rect 23293 30543 23351 30549
rect 23658 30540 23664 30592
rect 23716 30540 23722 30592
rect 26605 30583 26663 30589
rect 26605 30549 26617 30583
rect 26651 30580 26663 30583
rect 26694 30580 26700 30592
rect 26651 30552 26700 30580
rect 26651 30549 26663 30552
rect 26605 30543 26663 30549
rect 26694 30540 26700 30552
rect 26752 30580 26758 30592
rect 27706 30580 27712 30592
rect 26752 30552 27712 30580
rect 26752 30540 26758 30552
rect 27706 30540 27712 30552
rect 27764 30540 27770 30592
rect 1104 30490 49864 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 27950 30490
rect 28002 30438 28014 30490
rect 28066 30438 28078 30490
rect 28130 30438 28142 30490
rect 28194 30438 28206 30490
rect 28258 30438 37950 30490
rect 38002 30438 38014 30490
rect 38066 30438 38078 30490
rect 38130 30438 38142 30490
rect 38194 30438 38206 30490
rect 38258 30438 47950 30490
rect 48002 30438 48014 30490
rect 48066 30438 48078 30490
rect 48130 30438 48142 30490
rect 48194 30438 48206 30490
rect 48258 30438 49864 30490
rect 1104 30416 49864 30438
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 22738 30376 22744 30388
rect 12860 30348 22744 30376
rect 12860 30336 12866 30348
rect 16666 30308 16672 30320
rect 15594 30280 16672 30308
rect 16666 30268 16672 30280
rect 16724 30268 16730 30320
rect 19886 30308 19892 30320
rect 19720 30280 19892 30308
rect 1765 30243 1823 30249
rect 1765 30209 1777 30243
rect 1811 30240 1823 30243
rect 7374 30240 7380 30252
rect 1811 30212 7380 30240
rect 1811 30209 1823 30212
rect 1765 30203 1823 30209
rect 7374 30200 7380 30212
rect 7432 30200 7438 30252
rect 17405 30243 17463 30249
rect 17405 30209 17417 30243
rect 17451 30240 17463 30243
rect 18598 30240 18604 30252
rect 17451 30212 18604 30240
rect 17451 30209 17463 30212
rect 17405 30203 17463 30209
rect 18598 30200 18604 30212
rect 18656 30240 18662 30252
rect 19518 30240 19524 30252
rect 18656 30212 19524 30240
rect 18656 30200 18662 30212
rect 19518 30200 19524 30212
rect 19576 30200 19582 30252
rect 19720 30249 19748 30280
rect 19886 30268 19892 30280
rect 19944 30268 19950 30320
rect 20622 30268 20628 30320
rect 20680 30268 20686 30320
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30209 19763 30243
rect 19705 30203 19763 30209
rect 22186 30200 22192 30252
rect 22244 30200 22250 30252
rect 22664 30240 22692 30348
rect 22738 30336 22744 30348
rect 22796 30336 22802 30388
rect 23201 30379 23259 30385
rect 23201 30345 23213 30379
rect 23247 30376 23259 30379
rect 23382 30376 23388 30388
rect 23247 30348 23388 30376
rect 23247 30345 23259 30348
rect 23201 30339 23259 30345
rect 23382 30336 23388 30348
rect 23440 30336 23446 30388
rect 23658 30336 23664 30388
rect 23716 30376 23722 30388
rect 31018 30376 31024 30388
rect 23716 30348 31024 30376
rect 23716 30336 23722 30348
rect 31018 30336 31024 30348
rect 31076 30336 31082 30388
rect 33594 30336 33600 30388
rect 33652 30376 33658 30388
rect 40126 30376 40132 30388
rect 33652 30348 40132 30376
rect 33652 30336 33658 30348
rect 40126 30336 40132 30348
rect 40184 30336 40190 30388
rect 23293 30311 23351 30317
rect 23293 30277 23305 30311
rect 23339 30308 23351 30311
rect 23566 30308 23572 30320
rect 23339 30280 23572 30308
rect 23339 30277 23351 30280
rect 23293 30271 23351 30277
rect 23566 30268 23572 30280
rect 23624 30268 23630 30320
rect 30006 30240 30012 30252
rect 22664 30212 30012 30240
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 37366 30200 37372 30252
rect 37424 30240 37430 30252
rect 37645 30243 37703 30249
rect 37645 30240 37657 30243
rect 37424 30212 37657 30240
rect 37424 30200 37430 30212
rect 37645 30209 37657 30212
rect 37691 30209 37703 30243
rect 37645 30203 37703 30209
rect 49050 30200 49056 30252
rect 49108 30200 49114 30252
rect 1302 30132 1308 30184
rect 1360 30172 1366 30184
rect 2041 30175 2099 30181
rect 2041 30172 2053 30175
rect 1360 30144 2053 30172
rect 1360 30132 1366 30144
rect 2041 30141 2053 30144
rect 2087 30141 2099 30175
rect 2041 30135 2099 30141
rect 14090 30132 14096 30184
rect 14148 30132 14154 30184
rect 14369 30175 14427 30181
rect 14369 30172 14381 30175
rect 14200 30144 14381 30172
rect 13722 30064 13728 30116
rect 13780 30104 13786 30116
rect 14200 30104 14228 30144
rect 14369 30141 14381 30144
rect 14415 30172 14427 30175
rect 16206 30172 16212 30184
rect 14415 30144 16212 30172
rect 14415 30141 14427 30144
rect 14369 30135 14427 30141
rect 16206 30132 16212 30144
rect 16264 30132 16270 30184
rect 17126 30132 17132 30184
rect 17184 30172 17190 30184
rect 18141 30175 18199 30181
rect 18141 30172 18153 30175
rect 17184 30144 18153 30172
rect 17184 30132 17190 30144
rect 18141 30141 18153 30144
rect 18187 30141 18199 30175
rect 18141 30135 18199 30141
rect 19981 30175 20039 30181
rect 19981 30141 19993 30175
rect 20027 30172 20039 30175
rect 20346 30172 20352 30184
rect 20027 30144 20352 30172
rect 20027 30141 20039 30144
rect 19981 30135 20039 30141
rect 20346 30132 20352 30144
rect 20404 30172 20410 30184
rect 20990 30172 20996 30184
rect 20404 30144 20996 30172
rect 20404 30132 20410 30144
rect 20990 30132 20996 30144
rect 21048 30132 21054 30184
rect 21450 30132 21456 30184
rect 21508 30132 21514 30184
rect 23385 30175 23443 30181
rect 23385 30141 23397 30175
rect 23431 30141 23443 30175
rect 23385 30135 23443 30141
rect 13780 30076 14228 30104
rect 21008 30104 21036 30132
rect 23400 30104 23428 30135
rect 21008 30076 23428 30104
rect 13780 30064 13786 30076
rect 15841 30039 15899 30045
rect 15841 30005 15853 30039
rect 15887 30036 15899 30039
rect 15930 30036 15936 30048
rect 15887 30008 15936 30036
rect 15887 30005 15899 30008
rect 15841 29999 15899 30005
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 16298 29996 16304 30048
rect 16356 30036 16362 30048
rect 22002 30036 22008 30048
rect 16356 30008 22008 30036
rect 16356 29996 16362 30008
rect 22002 29996 22008 30008
rect 22060 29996 22066 30048
rect 22278 29996 22284 30048
rect 22336 30036 22342 30048
rect 22833 30039 22891 30045
rect 22833 30036 22845 30039
rect 22336 30008 22845 30036
rect 22336 29996 22342 30008
rect 22833 30005 22845 30008
rect 22879 30005 22891 30039
rect 22833 29999 22891 30005
rect 29086 29996 29092 30048
rect 29144 30036 29150 30048
rect 29273 30039 29331 30045
rect 29273 30036 29285 30039
rect 29144 30008 29285 30036
rect 29144 29996 29150 30008
rect 29273 30005 29285 30008
rect 29319 30005 29331 30039
rect 29273 29999 29331 30005
rect 37461 30039 37519 30045
rect 37461 30005 37473 30039
rect 37507 30036 37519 30039
rect 39390 30036 39396 30048
rect 37507 30008 39396 30036
rect 37507 30005 37519 30008
rect 37461 29999 37519 30005
rect 39390 29996 39396 30008
rect 39448 29996 39454 30048
rect 49234 29996 49240 30048
rect 49292 29996 49298 30048
rect 1104 29946 49864 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 32950 29946
rect 33002 29894 33014 29946
rect 33066 29894 33078 29946
rect 33130 29894 33142 29946
rect 33194 29894 33206 29946
rect 33258 29894 42950 29946
rect 43002 29894 43014 29946
rect 43066 29894 43078 29946
rect 43130 29894 43142 29946
rect 43194 29894 43206 29946
rect 43258 29894 49864 29946
rect 1104 29872 49864 29894
rect 19518 29792 19524 29844
rect 19576 29832 19582 29844
rect 27157 29835 27215 29841
rect 27157 29832 27169 29835
rect 19576 29804 27169 29832
rect 19576 29792 19582 29804
rect 27157 29801 27169 29804
rect 27203 29832 27215 29835
rect 27522 29832 27528 29844
rect 27203 29804 27528 29832
rect 27203 29801 27215 29804
rect 27157 29795 27215 29801
rect 27522 29792 27528 29804
rect 27580 29792 27586 29844
rect 49234 29832 49240 29844
rect 31726 29804 49240 29832
rect 31726 29764 31754 29804
rect 49234 29792 49240 29804
rect 49292 29792 49298 29844
rect 22066 29736 31754 29764
rect 1302 29656 1308 29708
rect 1360 29696 1366 29708
rect 2041 29699 2099 29705
rect 2041 29696 2053 29699
rect 1360 29668 2053 29696
rect 1360 29656 1366 29668
rect 2041 29665 2053 29668
rect 2087 29665 2099 29699
rect 15010 29696 15016 29708
rect 2041 29659 2099 29665
rect 14660 29668 15016 29696
rect 1765 29631 1823 29637
rect 1765 29597 1777 29631
rect 1811 29628 1823 29631
rect 8662 29628 8668 29640
rect 1811 29600 8668 29628
rect 1811 29597 1823 29600
rect 1765 29591 1823 29597
rect 8662 29588 8668 29600
rect 8720 29588 8726 29640
rect 14090 29588 14096 29640
rect 14148 29628 14154 29640
rect 14660 29637 14688 29668
rect 15010 29656 15016 29668
rect 15068 29696 15074 29708
rect 17126 29696 17132 29708
rect 15068 29668 17132 29696
rect 15068 29656 15074 29668
rect 17126 29656 17132 29668
rect 17184 29656 17190 29708
rect 18874 29656 18880 29708
rect 18932 29656 18938 29708
rect 20165 29699 20223 29705
rect 20165 29665 20177 29699
rect 20211 29696 20223 29699
rect 21450 29696 21456 29708
rect 20211 29668 21456 29696
rect 20211 29665 20223 29668
rect 20165 29659 20223 29665
rect 21450 29656 21456 29668
rect 21508 29656 21514 29708
rect 21910 29656 21916 29708
rect 21968 29656 21974 29708
rect 14645 29631 14703 29637
rect 14645 29628 14657 29631
rect 14148 29600 14657 29628
rect 14148 29588 14154 29600
rect 14645 29597 14657 29600
rect 14691 29597 14703 29631
rect 14645 29591 14703 29597
rect 16850 29588 16856 29640
rect 16908 29588 16914 29640
rect 19886 29588 19892 29640
rect 19944 29588 19950 29640
rect 14918 29520 14924 29572
rect 14976 29520 14982 29572
rect 16666 29560 16672 29572
rect 16146 29532 16672 29560
rect 16666 29520 16672 29532
rect 16724 29520 16730 29572
rect 17129 29563 17187 29569
rect 17129 29529 17141 29563
rect 17175 29529 17187 29563
rect 19058 29560 19064 29572
rect 18354 29532 19064 29560
rect 17129 29523 17187 29529
rect 14936 29492 14964 29520
rect 15930 29492 15936 29504
rect 14936 29464 15936 29492
rect 15930 29452 15936 29464
rect 15988 29452 15994 29504
rect 16390 29452 16396 29504
rect 16448 29452 16454 29504
rect 17144 29492 17172 29523
rect 19058 29520 19064 29532
rect 19116 29560 19122 29572
rect 20622 29560 20628 29572
rect 19116 29532 20628 29560
rect 19116 29520 19122 29532
rect 20622 29520 20628 29532
rect 20680 29520 20686 29572
rect 22066 29560 22094 29736
rect 28626 29656 28632 29708
rect 28684 29696 28690 29708
rect 28997 29699 29055 29705
rect 28997 29696 29009 29699
rect 28684 29668 29009 29696
rect 28684 29656 28690 29668
rect 28997 29665 29009 29668
rect 29043 29665 29055 29699
rect 49329 29699 49387 29705
rect 49329 29696 49341 29699
rect 28997 29659 29055 29665
rect 45526 29668 49341 29696
rect 22370 29588 22376 29640
rect 22428 29628 22434 29640
rect 22557 29631 22615 29637
rect 22557 29628 22569 29631
rect 22428 29600 22569 29628
rect 22428 29588 22434 29600
rect 22557 29597 22569 29600
rect 22603 29597 22615 29631
rect 22557 29591 22615 29597
rect 28813 29631 28871 29637
rect 28813 29597 28825 29631
rect 28859 29628 28871 29631
rect 29917 29631 29975 29637
rect 29917 29628 29929 29631
rect 28859 29600 29929 29628
rect 28859 29597 28871 29600
rect 28813 29591 28871 29597
rect 29917 29597 29929 29600
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 30006 29588 30012 29640
rect 30064 29628 30070 29640
rect 45526 29628 45554 29668
rect 49329 29665 49341 29668
rect 49375 29665 49387 29699
rect 49329 29659 49387 29665
rect 46569 29631 46627 29637
rect 46569 29628 46581 29631
rect 30064 29600 45554 29628
rect 45756 29600 46581 29628
rect 30064 29588 30070 29600
rect 21468 29532 22094 29560
rect 18782 29492 18788 29504
rect 17144 29464 18788 29492
rect 18782 29452 18788 29464
rect 18840 29452 18846 29504
rect 20530 29452 20536 29504
rect 20588 29492 20594 29504
rect 21468 29492 21496 29532
rect 25866 29520 25872 29572
rect 25924 29520 25930 29572
rect 32306 29560 32312 29572
rect 28460 29532 32312 29560
rect 20588 29464 21496 29492
rect 20588 29452 20594 29464
rect 22002 29452 22008 29504
rect 22060 29492 22066 29504
rect 24486 29492 24492 29504
rect 22060 29464 24492 29492
rect 22060 29452 22066 29464
rect 24486 29452 24492 29464
rect 24544 29452 24550 29504
rect 28460 29501 28488 29532
rect 32306 29520 32312 29532
rect 32364 29520 32370 29572
rect 28445 29495 28503 29501
rect 28445 29461 28457 29495
rect 28491 29461 28503 29495
rect 28445 29455 28503 29461
rect 28905 29495 28963 29501
rect 28905 29461 28917 29495
rect 28951 29492 28963 29495
rect 29178 29492 29184 29504
rect 28951 29464 29184 29492
rect 28951 29461 28963 29464
rect 28905 29455 28963 29461
rect 29178 29452 29184 29464
rect 29236 29452 29242 29504
rect 44174 29452 44180 29504
rect 44232 29492 44238 29504
rect 45756 29492 45784 29600
rect 46569 29597 46581 29600
rect 46615 29597 46627 29631
rect 46569 29591 46627 29597
rect 45830 29520 45836 29572
rect 45888 29520 45894 29572
rect 46753 29563 46811 29569
rect 46753 29529 46765 29563
rect 46799 29560 46811 29563
rect 47762 29560 47768 29572
rect 46799 29532 47768 29560
rect 46799 29529 46811 29532
rect 46753 29523 46811 29529
rect 47762 29520 47768 29532
rect 47820 29520 47826 29572
rect 49142 29520 49148 29572
rect 49200 29520 49206 29572
rect 44232 29464 45784 29492
rect 44232 29452 44238 29464
rect 45922 29452 45928 29504
rect 45980 29452 45986 29504
rect 1104 29402 49864 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 27950 29402
rect 28002 29350 28014 29402
rect 28066 29350 28078 29402
rect 28130 29350 28142 29402
rect 28194 29350 28206 29402
rect 28258 29350 37950 29402
rect 38002 29350 38014 29402
rect 38066 29350 38078 29402
rect 38130 29350 38142 29402
rect 38194 29350 38206 29402
rect 38258 29350 47950 29402
rect 48002 29350 48014 29402
rect 48066 29350 48078 29402
rect 48130 29350 48142 29402
rect 48194 29350 48206 29402
rect 48258 29350 49864 29402
rect 1104 29328 49864 29350
rect 14642 29248 14648 29300
rect 14700 29288 14706 29300
rect 15565 29291 15623 29297
rect 15565 29288 15577 29291
rect 14700 29260 15577 29288
rect 14700 29248 14706 29260
rect 15565 29257 15577 29260
rect 15611 29257 15623 29291
rect 15565 29251 15623 29257
rect 16022 29248 16028 29300
rect 16080 29248 16086 29300
rect 16114 29248 16120 29300
rect 16172 29288 16178 29300
rect 16298 29288 16304 29300
rect 16172 29260 16304 29288
rect 16172 29248 16178 29260
rect 16298 29248 16304 29260
rect 16356 29248 16362 29300
rect 16850 29248 16856 29300
rect 16908 29288 16914 29300
rect 16908 29260 19748 29288
rect 16908 29248 16914 29260
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29152 15991 29155
rect 16022 29152 16028 29164
rect 15979 29124 16028 29152
rect 15979 29121 15991 29124
rect 15933 29115 15991 29121
rect 16022 29112 16028 29124
rect 16080 29112 16086 29164
rect 17328 29161 17356 29260
rect 19058 29220 19064 29232
rect 18814 29192 19064 29220
rect 19058 29180 19064 29192
rect 19116 29180 19122 29232
rect 19720 29220 19748 29260
rect 21450 29248 21456 29300
rect 21508 29248 21514 29300
rect 21818 29248 21824 29300
rect 21876 29288 21882 29300
rect 22005 29291 22063 29297
rect 22005 29288 22017 29291
rect 21876 29260 22017 29288
rect 21876 29248 21882 29260
rect 22005 29257 22017 29260
rect 22051 29257 22063 29291
rect 22005 29251 22063 29257
rect 22370 29248 22376 29300
rect 22428 29248 22434 29300
rect 24949 29291 25007 29297
rect 24949 29257 24961 29291
rect 24995 29288 25007 29291
rect 25314 29288 25320 29300
rect 24995 29260 25320 29288
rect 24995 29257 25007 29260
rect 24949 29251 25007 29257
rect 25314 29248 25320 29260
rect 25372 29248 25378 29300
rect 28721 29291 28779 29297
rect 28721 29257 28733 29291
rect 28767 29288 28779 29291
rect 28810 29288 28816 29300
rect 28767 29260 28816 29288
rect 28767 29257 28779 29260
rect 28721 29251 28779 29257
rect 28810 29248 28816 29260
rect 28868 29248 28874 29300
rect 29086 29248 29092 29300
rect 29144 29248 29150 29300
rect 19886 29220 19892 29232
rect 19720 29192 19892 29220
rect 19720 29161 19748 29192
rect 19886 29180 19892 29192
rect 19944 29220 19950 29232
rect 20254 29220 20260 29232
rect 19944 29192 20260 29220
rect 19944 29180 19950 29192
rect 20254 29180 20260 29192
rect 20312 29180 20318 29232
rect 20622 29180 20628 29232
rect 20680 29180 20686 29232
rect 24486 29180 24492 29232
rect 24544 29220 24550 29232
rect 25409 29223 25467 29229
rect 25409 29220 25421 29223
rect 24544 29192 25421 29220
rect 24544 29180 24550 29192
rect 25409 29189 25421 29192
rect 25455 29220 25467 29223
rect 32398 29220 32404 29232
rect 25455 29192 32404 29220
rect 25455 29189 25467 29192
rect 25409 29183 25467 29189
rect 32398 29180 32404 29192
rect 32456 29220 32462 29232
rect 32766 29220 32772 29232
rect 32456 29192 32772 29220
rect 32456 29180 32462 29192
rect 32766 29180 32772 29192
rect 32824 29180 32830 29232
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29121 17371 29155
rect 17313 29115 17371 29121
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 22465 29155 22523 29161
rect 22465 29121 22477 29155
rect 22511 29152 22523 29155
rect 25314 29152 25320 29164
rect 22511 29124 25320 29152
rect 22511 29121 22523 29124
rect 22465 29115 22523 29121
rect 25314 29112 25320 29124
rect 25372 29112 25378 29164
rect 28902 29112 28908 29164
rect 28960 29152 28966 29164
rect 28960 29124 29316 29152
rect 28960 29112 28966 29124
rect 16209 29087 16267 29093
rect 16209 29053 16221 29087
rect 16255 29084 16267 29087
rect 17218 29084 17224 29096
rect 16255 29056 17224 29084
rect 16255 29053 16267 29056
rect 16209 29047 16267 29053
rect 17218 29044 17224 29056
rect 17276 29044 17282 29096
rect 17586 29044 17592 29096
rect 17644 29044 17650 29096
rect 17678 29044 17684 29096
rect 17736 29084 17742 29096
rect 18598 29084 18604 29096
rect 17736 29056 18604 29084
rect 17736 29044 17742 29056
rect 18598 29044 18604 29056
rect 18656 29084 18662 29096
rect 19061 29087 19119 29093
rect 19061 29084 19073 29087
rect 18656 29056 19073 29084
rect 18656 29044 18662 29056
rect 19061 29053 19073 29056
rect 19107 29053 19119 29087
rect 19061 29047 19119 29053
rect 22646 29044 22652 29096
rect 22704 29044 22710 29096
rect 25593 29087 25651 29093
rect 25593 29053 25605 29087
rect 25639 29084 25651 29087
rect 27062 29084 27068 29096
rect 25639 29056 27068 29084
rect 25639 29053 25651 29056
rect 25593 29047 25651 29053
rect 27062 29044 27068 29056
rect 27120 29044 27126 29096
rect 29178 29044 29184 29096
rect 29236 29044 29242 29096
rect 29288 29093 29316 29124
rect 29273 29087 29331 29093
rect 29273 29053 29285 29087
rect 29319 29053 29331 29087
rect 29273 29047 29331 29053
rect 17402 28908 17408 28960
rect 17460 28948 17466 28960
rect 17678 28948 17684 28960
rect 17460 28920 17684 28948
rect 17460 28908 17466 28920
rect 17678 28908 17684 28920
rect 17736 28908 17742 28960
rect 19968 28951 20026 28957
rect 19968 28917 19980 28951
rect 20014 28948 20026 28951
rect 21542 28948 21548 28960
rect 20014 28920 21548 28948
rect 20014 28917 20026 28920
rect 19968 28911 20026 28917
rect 21542 28908 21548 28920
rect 21600 28908 21606 28960
rect 1104 28858 49864 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 32950 28858
rect 33002 28806 33014 28858
rect 33066 28806 33078 28858
rect 33130 28806 33142 28858
rect 33194 28806 33206 28858
rect 33258 28806 42950 28858
rect 43002 28806 43014 28858
rect 43066 28806 43078 28858
rect 43130 28806 43142 28858
rect 43194 28806 43206 28858
rect 43258 28806 49864 28858
rect 1104 28784 49864 28806
rect 17586 28704 17592 28756
rect 17644 28744 17650 28756
rect 18690 28744 18696 28756
rect 17644 28716 18696 28744
rect 17644 28704 17650 28716
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 18782 28704 18788 28756
rect 18840 28744 18846 28756
rect 18877 28747 18935 28753
rect 18877 28744 18889 28747
rect 18840 28716 18889 28744
rect 18840 28704 18846 28716
rect 18877 28713 18889 28716
rect 18923 28713 18935 28747
rect 18877 28707 18935 28713
rect 19886 28704 19892 28756
rect 19944 28744 19950 28756
rect 28442 28744 28448 28756
rect 19944 28716 28448 28744
rect 19944 28704 19950 28716
rect 28442 28704 28448 28716
rect 28500 28704 28506 28756
rect 19242 28636 19248 28688
rect 19300 28676 19306 28688
rect 23750 28676 23756 28688
rect 19300 28648 23756 28676
rect 19300 28636 19306 28648
rect 23750 28636 23756 28648
rect 23808 28636 23814 28688
rect 1302 28568 1308 28620
rect 1360 28608 1366 28620
rect 2041 28611 2099 28617
rect 2041 28608 2053 28611
rect 1360 28580 2053 28608
rect 1360 28568 1366 28580
rect 2041 28577 2053 28580
rect 2087 28577 2099 28611
rect 2041 28571 2099 28577
rect 15930 28568 15936 28620
rect 15988 28568 15994 28620
rect 17126 28568 17132 28620
rect 17184 28568 17190 28620
rect 17402 28568 17408 28620
rect 17460 28568 17466 28620
rect 21542 28568 21548 28620
rect 21600 28568 21606 28620
rect 1765 28543 1823 28549
rect 1765 28509 1777 28543
rect 1811 28540 1823 28543
rect 11054 28540 11060 28552
rect 1811 28512 11060 28540
rect 1811 28509 1823 28512
rect 1765 28503 1823 28509
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 15746 28500 15752 28552
rect 15804 28500 15810 28552
rect 19518 28500 19524 28552
rect 19576 28500 19582 28552
rect 21269 28543 21327 28549
rect 21269 28509 21281 28543
rect 21315 28540 21327 28543
rect 22278 28540 22284 28552
rect 21315 28512 22284 28540
rect 21315 28509 21327 28512
rect 21269 28503 21327 28509
rect 22278 28500 22284 28512
rect 22336 28500 22342 28552
rect 34790 28500 34796 28552
rect 34848 28540 34854 28552
rect 37277 28543 37335 28549
rect 37277 28540 37289 28543
rect 34848 28512 37289 28540
rect 34848 28500 34854 28512
rect 37277 28509 37289 28512
rect 37323 28509 37335 28543
rect 37277 28503 37335 28509
rect 49050 28500 49056 28552
rect 49108 28500 49114 28552
rect 19058 28472 19064 28484
rect 18630 28444 19064 28472
rect 19058 28432 19064 28444
rect 19116 28432 19122 28484
rect 20254 28432 20260 28484
rect 20312 28432 20318 28484
rect 26510 28432 26516 28484
rect 26568 28472 26574 28484
rect 26568 28444 45554 28472
rect 26568 28432 26574 28444
rect 15378 28364 15384 28416
rect 15436 28364 15442 28416
rect 15841 28407 15899 28413
rect 15841 28373 15853 28407
rect 15887 28404 15899 28407
rect 16942 28404 16948 28416
rect 15887 28376 16948 28404
rect 15887 28373 15899 28376
rect 15841 28367 15899 28373
rect 16942 28364 16948 28376
rect 17000 28364 17006 28416
rect 17310 28364 17316 28416
rect 17368 28404 17374 28416
rect 20162 28404 20168 28416
rect 17368 28376 20168 28404
rect 17368 28364 17374 28376
rect 20162 28364 20168 28376
rect 20220 28364 20226 28416
rect 20898 28364 20904 28416
rect 20956 28364 20962 28416
rect 21358 28364 21364 28416
rect 21416 28364 21422 28416
rect 37093 28407 37151 28413
rect 37093 28373 37105 28407
rect 37139 28404 37151 28407
rect 43898 28404 43904 28416
rect 37139 28376 43904 28404
rect 37139 28373 37151 28376
rect 37093 28367 37151 28373
rect 43898 28364 43904 28376
rect 43956 28364 43962 28416
rect 45526 28404 45554 28444
rect 49237 28407 49295 28413
rect 49237 28404 49249 28407
rect 45526 28376 49249 28404
rect 49237 28373 49249 28376
rect 49283 28373 49295 28407
rect 49237 28367 49295 28373
rect 1104 28314 49864 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 27950 28314
rect 28002 28262 28014 28314
rect 28066 28262 28078 28314
rect 28130 28262 28142 28314
rect 28194 28262 28206 28314
rect 28258 28262 37950 28314
rect 38002 28262 38014 28314
rect 38066 28262 38078 28314
rect 38130 28262 38142 28314
rect 38194 28262 38206 28314
rect 38258 28262 47950 28314
rect 48002 28262 48014 28314
rect 48066 28262 48078 28314
rect 48130 28262 48142 28314
rect 48194 28262 48206 28314
rect 48258 28262 49864 28314
rect 1104 28240 49864 28262
rect 15286 28160 15292 28212
rect 15344 28160 15350 28212
rect 16942 28160 16948 28212
rect 17000 28160 17006 28212
rect 17405 28203 17463 28209
rect 17405 28169 17417 28203
rect 17451 28200 17463 28203
rect 18509 28203 18567 28209
rect 18509 28200 18521 28203
rect 17451 28172 18521 28200
rect 17451 28169 17463 28172
rect 17405 28163 17463 28169
rect 18509 28169 18521 28172
rect 18555 28169 18567 28203
rect 18509 28163 18567 28169
rect 18877 28203 18935 28209
rect 18877 28169 18889 28203
rect 18923 28200 18935 28203
rect 19150 28200 19156 28212
rect 18923 28172 19156 28200
rect 18923 28169 18935 28172
rect 18877 28163 18935 28169
rect 19150 28160 19156 28172
rect 19208 28160 19214 28212
rect 19705 28203 19763 28209
rect 19705 28169 19717 28203
rect 19751 28200 19763 28203
rect 21358 28200 21364 28212
rect 19751 28172 21364 28200
rect 19751 28169 19763 28172
rect 19705 28163 19763 28169
rect 21358 28160 21364 28172
rect 21416 28160 21422 28212
rect 14277 28135 14335 28141
rect 14277 28101 14289 28135
rect 14323 28132 14335 28135
rect 15749 28135 15807 28141
rect 15749 28132 15761 28135
rect 14323 28104 15761 28132
rect 14323 28101 14335 28104
rect 14277 28095 14335 28101
rect 15749 28101 15761 28104
rect 15795 28132 15807 28135
rect 31754 28132 31760 28144
rect 15795 28104 31760 28132
rect 15795 28101 15807 28104
rect 15749 28095 15807 28101
rect 31754 28092 31760 28104
rect 31812 28092 31818 28144
rect 44082 28092 44088 28144
rect 44140 28132 44146 28144
rect 45189 28135 45247 28141
rect 45189 28132 45201 28135
rect 44140 28104 45201 28132
rect 44140 28092 44146 28104
rect 45189 28101 45201 28104
rect 45235 28101 45247 28135
rect 45189 28095 45247 28101
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28064 1823 28067
rect 11146 28064 11152 28076
rect 1811 28036 11152 28064
rect 1811 28033 1823 28036
rect 1765 28027 1823 28033
rect 11146 28024 11152 28036
rect 11204 28024 11210 28076
rect 14734 28024 14740 28076
rect 14792 28064 14798 28076
rect 15657 28067 15715 28073
rect 15657 28064 15669 28067
rect 14792 28036 15669 28064
rect 14792 28024 14798 28036
rect 15657 28033 15669 28036
rect 15703 28033 15715 28067
rect 15657 28027 15715 28033
rect 16206 28024 16212 28076
rect 16264 28064 16270 28076
rect 16264 28036 16620 28064
rect 16264 28024 16270 28036
rect 1302 27956 1308 28008
rect 1360 27996 1366 28008
rect 2041 27999 2099 28005
rect 2041 27996 2053 27999
rect 1360 27968 2053 27996
rect 1360 27956 1366 27968
rect 2041 27965 2053 27968
rect 2087 27965 2099 27999
rect 2041 27959 2099 27965
rect 15933 27999 15991 28005
rect 15933 27965 15945 27999
rect 15979 27996 15991 27999
rect 16482 27996 16488 28008
rect 15979 27968 16488 27996
rect 15979 27965 15991 27968
rect 15933 27959 15991 27965
rect 16482 27956 16488 27968
rect 16540 27956 16546 28008
rect 16592 27996 16620 28036
rect 17310 28024 17316 28076
rect 17368 28024 17374 28076
rect 18874 28024 18880 28076
rect 18932 28064 18938 28076
rect 18932 28036 19104 28064
rect 18932 28024 18938 28036
rect 19076 28005 19104 28036
rect 20070 28024 20076 28076
rect 20128 28064 20134 28076
rect 21634 28064 21640 28076
rect 20128 28036 21640 28064
rect 20128 28024 20134 28036
rect 21634 28024 21640 28036
rect 21692 28024 21698 28076
rect 49326 28024 49332 28076
rect 49384 28024 49390 28076
rect 17497 27999 17555 28005
rect 17497 27996 17509 27999
rect 16592 27968 17509 27996
rect 17497 27965 17509 27968
rect 17543 27965 17555 27999
rect 17497 27959 17555 27965
rect 18969 27999 19027 28005
rect 18969 27965 18981 27999
rect 19015 27965 19027 27999
rect 18969 27959 19027 27965
rect 19061 27999 19119 28005
rect 19061 27965 19073 27999
rect 19107 27965 19119 27999
rect 19061 27959 19119 27965
rect 18874 27888 18880 27940
rect 18932 27928 18938 27940
rect 18984 27928 19012 27959
rect 19702 27956 19708 28008
rect 19760 27996 19766 28008
rect 20165 27999 20223 28005
rect 20165 27996 20177 27999
rect 19760 27968 20177 27996
rect 19760 27956 19766 27968
rect 20165 27965 20177 27968
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 20346 27956 20352 28008
rect 20404 27956 20410 28008
rect 19242 27928 19248 27940
rect 18932 27900 19248 27928
rect 18932 27888 18938 27900
rect 19242 27888 19248 27900
rect 19300 27888 19306 27940
rect 36538 27888 36544 27940
rect 36596 27928 36602 27940
rect 49145 27931 49203 27937
rect 49145 27928 49157 27931
rect 36596 27900 49157 27928
rect 36596 27888 36602 27900
rect 49145 27897 49157 27900
rect 49191 27897 49203 27931
rect 49145 27891 49203 27897
rect 14734 27820 14740 27872
rect 14792 27820 14798 27872
rect 45278 27820 45284 27872
rect 45336 27820 45342 27872
rect 1104 27770 49864 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 32950 27770
rect 33002 27718 33014 27770
rect 33066 27718 33078 27770
rect 33130 27718 33142 27770
rect 33194 27718 33206 27770
rect 33258 27718 42950 27770
rect 43002 27718 43014 27770
rect 43066 27718 43078 27770
rect 43130 27718 43142 27770
rect 43194 27718 43206 27770
rect 43258 27718 49864 27770
rect 1104 27696 49864 27718
rect 18340 27628 19288 27656
rect 15381 27591 15439 27597
rect 15381 27557 15393 27591
rect 15427 27588 15439 27591
rect 16850 27588 16856 27600
rect 15427 27560 16856 27588
rect 15427 27557 15439 27560
rect 15381 27551 15439 27557
rect 16850 27548 16856 27560
rect 16908 27548 16914 27600
rect 18340 27588 18368 27628
rect 17052 27560 18368 27588
rect 15838 27480 15844 27532
rect 15896 27480 15902 27532
rect 16025 27523 16083 27529
rect 16025 27489 16037 27523
rect 16071 27520 16083 27523
rect 16390 27520 16396 27532
rect 16071 27492 16396 27520
rect 16071 27489 16083 27492
rect 16025 27483 16083 27489
rect 16390 27480 16396 27492
rect 16448 27480 16454 27532
rect 17052 27529 17080 27560
rect 18414 27548 18420 27600
rect 18472 27588 18478 27600
rect 19150 27588 19156 27600
rect 18472 27560 19156 27588
rect 18472 27548 18478 27560
rect 19150 27548 19156 27560
rect 19208 27548 19214 27600
rect 19260 27588 19288 27628
rect 20438 27588 20444 27600
rect 19260 27560 20444 27588
rect 20438 27548 20444 27560
rect 20496 27548 20502 27600
rect 17037 27523 17095 27529
rect 17037 27489 17049 27523
rect 17083 27489 17095 27523
rect 17037 27483 17095 27489
rect 17221 27523 17279 27529
rect 17221 27489 17233 27523
rect 17267 27520 17279 27523
rect 17586 27520 17592 27532
rect 17267 27492 17592 27520
rect 17267 27489 17279 27492
rect 17221 27483 17279 27489
rect 17586 27480 17592 27492
rect 17644 27480 17650 27532
rect 18598 27480 18604 27532
rect 18656 27520 18662 27532
rect 18693 27523 18751 27529
rect 18693 27520 18705 27523
rect 18656 27492 18705 27520
rect 18656 27480 18662 27492
rect 18693 27489 18705 27492
rect 18739 27489 18751 27523
rect 18693 27483 18751 27489
rect 15378 27412 15384 27464
rect 15436 27452 15442 27464
rect 15749 27455 15807 27461
rect 15749 27452 15761 27455
rect 15436 27424 15761 27452
rect 15436 27412 15442 27424
rect 15749 27421 15761 27424
rect 15795 27421 15807 27455
rect 15749 27415 15807 27421
rect 16942 27412 16948 27464
rect 17000 27412 17006 27464
rect 18509 27455 18567 27461
rect 18509 27421 18521 27455
rect 18555 27452 18567 27455
rect 18966 27452 18972 27464
rect 18555 27424 18972 27452
rect 18555 27421 18567 27424
rect 18509 27415 18567 27421
rect 18966 27412 18972 27424
rect 19024 27412 19030 27464
rect 18601 27387 18659 27393
rect 18601 27384 18613 27387
rect 16592 27356 18613 27384
rect 16592 27325 16620 27356
rect 18601 27353 18613 27356
rect 18647 27353 18659 27387
rect 18601 27347 18659 27353
rect 28350 27344 28356 27396
rect 28408 27384 28414 27396
rect 38933 27387 38991 27393
rect 38933 27384 38945 27387
rect 28408 27356 38945 27384
rect 28408 27344 28414 27356
rect 38933 27353 38945 27356
rect 38979 27353 38991 27387
rect 38933 27347 38991 27353
rect 39117 27387 39175 27393
rect 39117 27353 39129 27387
rect 39163 27384 39175 27387
rect 46842 27384 46848 27396
rect 39163 27356 46848 27384
rect 39163 27353 39175 27356
rect 39117 27347 39175 27353
rect 46842 27344 46848 27356
rect 46900 27344 46906 27396
rect 16577 27319 16635 27325
rect 16577 27285 16589 27319
rect 16623 27285 16635 27319
rect 16577 27279 16635 27285
rect 18141 27319 18199 27325
rect 18141 27285 18153 27319
rect 18187 27316 18199 27319
rect 18414 27316 18420 27328
rect 18187 27288 18420 27316
rect 18187 27285 18199 27288
rect 18141 27279 18199 27285
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 1104 27226 49864 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 27950 27226
rect 28002 27174 28014 27226
rect 28066 27174 28078 27226
rect 28130 27174 28142 27226
rect 28194 27174 28206 27226
rect 28258 27174 37950 27226
rect 38002 27174 38014 27226
rect 38066 27174 38078 27226
rect 38130 27174 38142 27226
rect 38194 27174 38206 27226
rect 38258 27174 47950 27226
rect 48002 27174 48014 27226
rect 48066 27174 48078 27226
rect 48130 27174 48142 27226
rect 48194 27174 48206 27226
rect 48258 27174 49864 27226
rect 1104 27152 49864 27174
rect 20898 27072 20904 27124
rect 20956 27112 20962 27124
rect 21085 27115 21143 27121
rect 21085 27112 21097 27115
rect 20956 27084 21097 27112
rect 20956 27072 20962 27084
rect 21085 27081 21097 27084
rect 21131 27081 21143 27115
rect 21085 27075 21143 27081
rect 19794 27004 19800 27056
rect 19852 27044 19858 27056
rect 21177 27047 21235 27053
rect 21177 27044 21189 27047
rect 19852 27016 21189 27044
rect 19852 27004 19858 27016
rect 21177 27013 21189 27016
rect 21223 27013 21235 27047
rect 21177 27007 21235 27013
rect 44542 27004 44548 27056
rect 44600 27004 44606 27056
rect 934 26936 940 26988
rect 992 26976 998 26988
rect 1673 26979 1731 26985
rect 1673 26976 1685 26979
rect 992 26948 1685 26976
rect 992 26936 998 26948
rect 1673 26945 1685 26948
rect 1719 26945 1731 26979
rect 1673 26939 1731 26945
rect 46750 26936 46756 26988
rect 46808 26976 46814 26988
rect 47949 26979 48007 26985
rect 47949 26976 47961 26979
rect 46808 26948 47961 26976
rect 46808 26936 46814 26948
rect 47949 26945 47961 26948
rect 47995 26945 48007 26979
rect 47949 26939 48007 26945
rect 21361 26911 21419 26917
rect 21361 26877 21373 26911
rect 21407 26908 21419 26911
rect 21450 26908 21456 26920
rect 21407 26880 21456 26908
rect 21407 26877 21419 26880
rect 21361 26871 21419 26877
rect 21450 26868 21456 26880
rect 21508 26868 21514 26920
rect 49142 26868 49148 26920
rect 49200 26868 49206 26920
rect 44726 26800 44732 26852
rect 44784 26800 44790 26852
rect 1765 26775 1823 26781
rect 1765 26741 1777 26775
rect 1811 26772 1823 26775
rect 12434 26772 12440 26784
rect 1811 26744 12440 26772
rect 1811 26741 1823 26744
rect 1765 26735 1823 26741
rect 12434 26732 12440 26744
rect 12492 26732 12498 26784
rect 20717 26775 20775 26781
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 22278 26772 22284 26784
rect 20763 26744 22284 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 22278 26732 22284 26744
rect 22336 26732 22342 26784
rect 1104 26682 49864 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 32950 26682
rect 33002 26630 33014 26682
rect 33066 26630 33078 26682
rect 33130 26630 33142 26682
rect 33194 26630 33206 26682
rect 33258 26630 42950 26682
rect 43002 26630 43014 26682
rect 43066 26630 43078 26682
rect 43130 26630 43142 26682
rect 43194 26630 43206 26682
rect 43258 26630 49864 26682
rect 1104 26608 49864 26630
rect 18141 26503 18199 26509
rect 18141 26469 18153 26503
rect 18187 26500 18199 26503
rect 20162 26500 20168 26512
rect 18187 26472 20168 26500
rect 18187 26469 18199 26472
rect 18141 26463 18199 26469
rect 20162 26460 20168 26472
rect 20220 26460 20226 26512
rect 18598 26392 18604 26444
rect 18656 26392 18662 26444
rect 18782 26392 18788 26444
rect 18840 26392 18846 26444
rect 48222 26392 48228 26444
rect 48280 26432 48286 26444
rect 48409 26435 48467 26441
rect 48409 26432 48421 26435
rect 48280 26404 48421 26432
rect 48280 26392 48286 26404
rect 48409 26401 48421 26404
rect 48455 26401 48467 26435
rect 48409 26395 48467 26401
rect 1857 26367 1915 26373
rect 1857 26333 1869 26367
rect 1903 26364 1915 26367
rect 12618 26364 12624 26376
rect 1903 26336 12624 26364
rect 1903 26333 1915 26336
rect 1857 26327 1915 26333
rect 12618 26324 12624 26336
rect 12676 26324 12682 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18509 26367 18567 26373
rect 18509 26364 18521 26367
rect 18472 26336 18521 26364
rect 18472 26324 18478 26336
rect 18509 26333 18521 26336
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 46474 26324 46480 26376
rect 46532 26364 46538 26376
rect 47949 26367 48007 26373
rect 47949 26364 47961 26367
rect 46532 26336 47961 26364
rect 46532 26324 46538 26336
rect 47949 26333 47961 26336
rect 47995 26333 48007 26367
rect 47949 26327 48007 26333
rect 1670 26256 1676 26308
rect 1728 26256 1734 26308
rect 1104 26138 49864 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 27950 26138
rect 28002 26086 28014 26138
rect 28066 26086 28078 26138
rect 28130 26086 28142 26138
rect 28194 26086 28206 26138
rect 28258 26086 37950 26138
rect 38002 26086 38014 26138
rect 38066 26086 38078 26138
rect 38130 26086 38142 26138
rect 38194 26086 38206 26138
rect 38258 26086 47950 26138
rect 48002 26086 48014 26138
rect 48066 26086 48078 26138
rect 48130 26086 48142 26138
rect 48194 26086 48206 26138
rect 48258 26086 49864 26138
rect 1104 26064 49864 26086
rect 29638 25916 29644 25968
rect 29696 25956 29702 25968
rect 38841 25959 38899 25965
rect 38841 25956 38853 25959
rect 29696 25928 38853 25956
rect 29696 25916 29702 25928
rect 38841 25925 38853 25928
rect 38887 25925 38899 25959
rect 38841 25919 38899 25925
rect 37826 25848 37832 25900
rect 37884 25888 37890 25900
rect 38197 25891 38255 25897
rect 38197 25888 38209 25891
rect 37884 25860 38209 25888
rect 37884 25848 37890 25860
rect 38197 25857 38209 25860
rect 38243 25857 38255 25891
rect 38197 25851 38255 25857
rect 39025 25755 39083 25761
rect 39025 25721 39037 25755
rect 39071 25752 39083 25755
rect 44266 25752 44272 25764
rect 39071 25724 44272 25752
rect 39071 25721 39083 25724
rect 39025 25715 39083 25721
rect 44266 25712 44272 25724
rect 44324 25712 44330 25764
rect 38013 25687 38071 25693
rect 38013 25653 38025 25687
rect 38059 25684 38071 25687
rect 39942 25684 39948 25696
rect 38059 25656 39948 25684
rect 38059 25653 38071 25656
rect 38013 25647 38071 25653
rect 39942 25644 39948 25656
rect 40000 25644 40006 25696
rect 1104 25594 49864 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 32950 25594
rect 33002 25542 33014 25594
rect 33066 25542 33078 25594
rect 33130 25542 33142 25594
rect 33194 25542 33206 25594
rect 33258 25542 42950 25594
rect 43002 25542 43014 25594
rect 43066 25542 43078 25594
rect 43130 25542 43142 25594
rect 43194 25542 43206 25594
rect 43258 25542 49864 25594
rect 1104 25520 49864 25542
rect 1857 25347 1915 25353
rect 1857 25313 1869 25347
rect 1903 25344 1915 25347
rect 3418 25344 3424 25356
rect 1903 25316 3424 25344
rect 1903 25313 1915 25316
rect 1857 25307 1915 25313
rect 3418 25304 3424 25316
rect 3476 25304 3482 25356
rect 934 25236 940 25288
rect 992 25276 998 25288
rect 1581 25279 1639 25285
rect 1581 25276 1593 25279
rect 992 25248 1593 25276
rect 992 25236 998 25248
rect 1581 25245 1593 25248
rect 1627 25245 1639 25279
rect 1581 25239 1639 25245
rect 45922 25236 45928 25288
rect 45980 25276 45986 25288
rect 47949 25279 48007 25285
rect 47949 25276 47961 25279
rect 45980 25248 47961 25276
rect 45980 25236 45986 25248
rect 47949 25245 47961 25248
rect 47995 25245 48007 25279
rect 47949 25239 48007 25245
rect 49142 25236 49148 25288
rect 49200 25236 49206 25288
rect 1104 25050 49864 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 27950 25050
rect 28002 24998 28014 25050
rect 28066 24998 28078 25050
rect 28130 24998 28142 25050
rect 28194 24998 28206 25050
rect 28258 24998 37950 25050
rect 38002 24998 38014 25050
rect 38066 24998 38078 25050
rect 38130 24998 38142 25050
rect 38194 24998 38206 25050
rect 38258 24998 47950 25050
rect 48002 24998 48014 25050
rect 48066 24998 48078 25050
rect 48130 24998 48142 25050
rect 48194 24998 48206 25050
rect 48258 24998 49864 25050
rect 1104 24976 49864 24998
rect 934 24760 940 24812
rect 992 24800 998 24812
rect 1673 24803 1731 24809
rect 1673 24800 1685 24803
rect 992 24772 1685 24800
rect 992 24760 998 24772
rect 1673 24769 1685 24772
rect 1719 24769 1731 24803
rect 1673 24763 1731 24769
rect 28442 24760 28448 24812
rect 28500 24800 28506 24812
rect 39577 24803 39635 24809
rect 39577 24800 39589 24803
rect 28500 24772 39589 24800
rect 28500 24760 28506 24772
rect 39577 24769 39589 24772
rect 39623 24769 39635 24803
rect 39577 24763 39635 24769
rect 39945 24803 40003 24809
rect 39945 24769 39957 24803
rect 39991 24769 40003 24803
rect 39945 24763 40003 24769
rect 39298 24692 39304 24744
rect 39356 24732 39362 24744
rect 39960 24732 39988 24763
rect 47762 24760 47768 24812
rect 47820 24800 47826 24812
rect 47949 24803 48007 24809
rect 47949 24800 47961 24803
rect 47820 24772 47961 24800
rect 47820 24760 47826 24772
rect 47949 24769 47961 24772
rect 47995 24769 48007 24803
rect 47949 24763 48007 24769
rect 39356 24704 39988 24732
rect 39356 24692 39362 24704
rect 49142 24692 49148 24744
rect 49200 24692 49206 24744
rect 39761 24667 39819 24673
rect 39761 24633 39773 24667
rect 39807 24664 39819 24667
rect 44174 24664 44180 24676
rect 39807 24636 44180 24664
rect 39807 24633 39819 24636
rect 39761 24627 39819 24633
rect 44174 24624 44180 24636
rect 44232 24624 44238 24676
rect 1949 24599 2007 24605
rect 1949 24565 1961 24599
rect 1995 24596 2007 24599
rect 14826 24596 14832 24608
rect 1995 24568 14832 24596
rect 1995 24565 2007 24568
rect 1949 24559 2007 24565
rect 14826 24556 14832 24568
rect 14884 24556 14890 24608
rect 40037 24599 40095 24605
rect 40037 24565 40049 24599
rect 40083 24596 40095 24599
rect 46934 24596 46940 24608
rect 40083 24568 46940 24596
rect 40083 24565 40095 24568
rect 40037 24559 40095 24565
rect 46934 24556 46940 24568
rect 46992 24556 46998 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 13354 24148 13360 24200
rect 13412 24188 13418 24200
rect 15841 24191 15899 24197
rect 15841 24188 15853 24191
rect 13412 24160 15853 24188
rect 13412 24148 13418 24160
rect 15841 24157 15853 24160
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 37645 24191 37703 24197
rect 37645 24188 37657 24191
rect 33836 24160 37657 24188
rect 33836 24148 33842 24160
rect 37645 24157 37657 24160
rect 37691 24157 37703 24191
rect 37645 24151 37703 24157
rect 39390 24148 39396 24200
rect 39448 24188 39454 24200
rect 44085 24191 44143 24197
rect 44085 24188 44097 24191
rect 39448 24160 44097 24188
rect 39448 24148 39454 24160
rect 44085 24157 44097 24160
rect 44131 24157 44143 24191
rect 44085 24151 44143 24157
rect 44269 24123 44327 24129
rect 44269 24089 44281 24123
rect 44315 24120 44327 24123
rect 45094 24120 45100 24132
rect 44315 24092 45100 24120
rect 44315 24089 44327 24092
rect 44269 24083 44327 24089
rect 45094 24080 45100 24092
rect 45152 24080 45158 24132
rect 15654 24012 15660 24064
rect 15712 24012 15718 24064
rect 37461 24055 37519 24061
rect 37461 24021 37473 24055
rect 37507 24052 37519 24055
rect 43438 24052 43444 24064
rect 37507 24024 43444 24052
rect 37507 24021 37519 24024
rect 37461 24015 37519 24021
rect 43438 24012 43444 24024
rect 43496 24012 43502 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 1857 23783 1915 23789
rect 1857 23749 1869 23783
rect 1903 23780 1915 23783
rect 4890 23780 4896 23792
rect 1903 23752 4896 23780
rect 1903 23749 1915 23752
rect 1857 23743 1915 23749
rect 4890 23740 4896 23752
rect 4948 23740 4954 23792
rect 33410 23740 33416 23792
rect 33468 23780 33474 23792
rect 39117 23783 39175 23789
rect 39117 23780 39129 23783
rect 33468 23752 39129 23780
rect 33468 23740 33474 23752
rect 39117 23749 39129 23752
rect 39163 23749 39175 23783
rect 39117 23743 39175 23749
rect 934 23672 940 23724
rect 992 23712 998 23724
rect 1673 23715 1731 23721
rect 1673 23712 1685 23715
rect 992 23684 1685 23712
rect 992 23672 998 23684
rect 1673 23681 1685 23684
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 32030 23672 32036 23724
rect 32088 23712 32094 23724
rect 36909 23715 36967 23721
rect 36909 23712 36921 23715
rect 32088 23684 36921 23712
rect 32088 23672 32094 23684
rect 36909 23681 36921 23684
rect 36955 23681 36967 23715
rect 36909 23675 36967 23681
rect 46842 23672 46848 23724
rect 46900 23712 46906 23724
rect 47949 23715 48007 23721
rect 47949 23712 47961 23715
rect 46900 23684 47961 23712
rect 46900 23672 46906 23684
rect 47949 23681 47961 23684
rect 47995 23681 48007 23715
rect 47949 23675 48007 23681
rect 49142 23604 49148 23656
rect 49200 23604 49206 23656
rect 39301 23579 39359 23585
rect 39301 23545 39313 23579
rect 39347 23576 39359 23579
rect 47026 23576 47032 23588
rect 39347 23548 47032 23576
rect 39347 23545 39359 23548
rect 39301 23539 39359 23545
rect 47026 23536 47032 23548
rect 47084 23536 47090 23588
rect 36722 23468 36728 23520
rect 36780 23468 36786 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 1857 23171 1915 23177
rect 1857 23137 1869 23171
rect 1903 23168 1915 23171
rect 4798 23168 4804 23180
rect 1903 23140 4804 23168
rect 1903 23137 1915 23140
rect 1857 23131 1915 23137
rect 4798 23128 4804 23140
rect 4856 23128 4862 23180
rect 934 23060 940 23112
rect 992 23100 998 23112
rect 1581 23103 1639 23109
rect 1581 23100 1593 23103
rect 992 23072 1593 23100
rect 992 23060 998 23072
rect 1581 23069 1593 23072
rect 1627 23069 1639 23103
rect 1581 23063 1639 23069
rect 45278 23060 45284 23112
rect 45336 23100 45342 23112
rect 47949 23103 48007 23109
rect 47949 23100 47961 23103
rect 45336 23072 47961 23100
rect 45336 23060 45342 23072
rect 47949 23069 47961 23072
rect 47995 23069 48007 23103
rect 47949 23063 48007 23069
rect 49142 22992 49148 23044
rect 49200 22992 49206 23044
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 43898 21972 43904 22024
rect 43956 21972 43962 22024
rect 44726 21972 44732 22024
rect 44784 22012 44790 22024
rect 47949 22015 48007 22021
rect 47949 22012 47961 22015
rect 44784 21984 47961 22012
rect 44784 21972 44790 21984
rect 47949 21981 47961 21984
rect 47995 21981 48007 22015
rect 47949 21975 48007 21981
rect 49142 21972 49148 22024
rect 49200 21972 49206 22024
rect 934 21904 940 21956
rect 992 21944 998 21956
rect 1673 21947 1731 21953
rect 1673 21944 1685 21947
rect 992 21916 1685 21944
rect 992 21904 998 21916
rect 1673 21913 1685 21916
rect 1719 21913 1731 21947
rect 1673 21907 1731 21913
rect 44085 21947 44143 21953
rect 44085 21913 44097 21947
rect 44131 21944 44143 21947
rect 44818 21944 44824 21956
rect 44131 21916 44824 21944
rect 44131 21913 44143 21916
rect 44085 21907 44143 21913
rect 44818 21904 44824 21916
rect 44876 21904 44882 21956
rect 1949 21879 2007 21885
rect 1949 21845 1961 21879
rect 1995 21876 2007 21879
rect 19150 21876 19156 21888
rect 1995 21848 19156 21876
rect 1995 21845 2007 21848
rect 1949 21839 2007 21845
rect 19150 21836 19156 21848
rect 19208 21836 19214 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 934 21496 940 21548
rect 992 21536 998 21548
rect 1673 21539 1731 21545
rect 1673 21536 1685 21539
rect 992 21508 1685 21536
rect 992 21496 998 21508
rect 1673 21505 1685 21508
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 26694 21496 26700 21548
rect 26752 21536 26758 21548
rect 37553 21539 37611 21545
rect 37553 21536 37565 21539
rect 26752 21508 37565 21536
rect 26752 21496 26758 21508
rect 37553 21505 37565 21508
rect 37599 21505 37611 21539
rect 37553 21499 37611 21505
rect 44266 21496 44272 21548
rect 44324 21536 44330 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 44324 21508 47961 21536
rect 44324 21496 44330 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 37737 21403 37795 21409
rect 37737 21369 37749 21403
rect 37783 21400 37795 21403
rect 42794 21400 42800 21412
rect 37783 21372 42800 21400
rect 37783 21369 37795 21372
rect 37737 21363 37795 21369
rect 42794 21360 42800 21372
rect 42852 21360 42858 21412
rect 1949 21335 2007 21341
rect 1949 21301 1961 21335
rect 1995 21332 2007 21335
rect 19886 21332 19892 21344
rect 1995 21304 19892 21332
rect 1995 21301 2007 21304
rect 1949 21295 2007 21301
rect 19886 21292 19892 21304
rect 19944 21292 19950 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 32214 20816 32220 20868
rect 32272 20856 32278 20868
rect 40129 20859 40187 20865
rect 40129 20856 40141 20859
rect 32272 20828 40141 20856
rect 32272 20816 32278 20828
rect 40129 20825 40141 20828
rect 40175 20825 40187 20859
rect 40129 20819 40187 20825
rect 40313 20859 40371 20865
rect 40313 20825 40325 20859
rect 40359 20856 40371 20859
rect 47762 20856 47768 20868
rect 40359 20828 47768 20856
rect 40359 20825 40371 20828
rect 40313 20819 40371 20825
rect 47762 20816 47768 20828
rect 47820 20816 47826 20868
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 934 20408 940 20460
rect 992 20448 998 20460
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 992 20420 1685 20448
rect 992 20408 998 20420
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 44174 20408 44180 20460
rect 44232 20448 44238 20460
rect 47949 20451 48007 20457
rect 47949 20448 47961 20451
rect 44232 20420 47961 20448
rect 44232 20408 44238 20420
rect 47949 20417 47961 20420
rect 47995 20417 48007 20451
rect 47949 20411 48007 20417
rect 49142 20340 49148 20392
rect 49200 20340 49206 20392
rect 1949 20247 2007 20253
rect 1949 20213 1961 20247
rect 1995 20244 2007 20247
rect 16758 20244 16764 20256
rect 1995 20216 16764 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 46934 19796 46940 19848
rect 46992 19836 46998 19848
rect 47949 19839 48007 19845
rect 47949 19836 47961 19839
rect 46992 19808 47961 19836
rect 46992 19796 46998 19808
rect 47949 19805 47961 19808
rect 47995 19805 48007 19839
rect 47949 19799 48007 19805
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 1673 19771 1731 19777
rect 1673 19768 1685 19771
rect 992 19740 1685 19768
rect 992 19728 998 19740
rect 1673 19737 1685 19740
rect 1719 19737 1731 19771
rect 1673 19731 1731 19737
rect 49142 19728 49148 19780
rect 49200 19728 49206 19780
rect 1765 19703 1823 19709
rect 1765 19669 1777 19703
rect 1811 19700 1823 19703
rect 17034 19700 17040 19712
rect 1811 19672 17040 19700
rect 1811 19669 1823 19672
rect 1765 19663 1823 19669
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 17773 19499 17831 19505
rect 17773 19465 17785 19499
rect 17819 19496 17831 19499
rect 19978 19496 19984 19508
rect 17819 19468 19984 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 22186 19496 22192 19508
rect 22143 19468 22192 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 22186 19456 22192 19468
rect 22244 19456 22250 19508
rect 39942 19388 39948 19440
rect 40000 19428 40006 19440
rect 44453 19431 44511 19437
rect 44453 19428 44465 19431
rect 40000 19400 44465 19428
rect 40000 19388 40006 19400
rect 44453 19397 44465 19400
rect 44499 19397 44511 19431
rect 44453 19391 44511 19397
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17957 19363 18015 19369
rect 17957 19360 17969 19363
rect 16908 19332 17969 19360
rect 16908 19320 16914 19332
rect 17957 19329 17969 19332
rect 18003 19329 18015 19363
rect 17957 19323 18015 19329
rect 22278 19320 22284 19372
rect 22336 19320 22342 19372
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 38657 19363 38715 19369
rect 38657 19360 38669 19363
rect 32456 19332 38669 19360
rect 32456 19320 32462 19332
rect 38657 19329 38669 19332
rect 38703 19329 38715 19363
rect 38657 19323 38715 19329
rect 38841 19227 38899 19233
rect 38841 19193 38853 19227
rect 38887 19224 38899 19227
rect 44266 19224 44272 19236
rect 38887 19196 44272 19224
rect 38887 19193 38899 19196
rect 38841 19187 38899 19193
rect 44266 19184 44272 19196
rect 44324 19184 44330 19236
rect 44637 19227 44695 19233
rect 44637 19193 44649 19227
rect 44683 19224 44695 19227
rect 46934 19224 46940 19236
rect 44683 19196 46940 19224
rect 44683 19193 44695 19196
rect 44637 19187 44695 19193
rect 46934 19184 46940 19196
rect 46992 19184 46998 19236
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1581 18751 1639 18757
rect 1581 18748 1593 18751
rect 992 18720 1593 18748
rect 992 18708 998 18720
rect 1581 18717 1593 18720
rect 1627 18717 1639 18751
rect 1581 18711 1639 18717
rect 20162 18708 20168 18760
rect 20220 18708 20226 18760
rect 40126 18708 40132 18760
rect 40184 18708 40190 18760
rect 45094 18708 45100 18760
rect 45152 18748 45158 18760
rect 47949 18751 48007 18757
rect 47949 18748 47961 18751
rect 45152 18720 47961 18748
rect 45152 18708 45158 18720
rect 47949 18717 47961 18720
rect 47995 18717 48007 18751
rect 47949 18711 48007 18717
rect 49142 18708 49148 18760
rect 49200 18708 49206 18760
rect 33410 18680 33416 18692
rect 6886 18652 33416 18680
rect 1765 18615 1823 18621
rect 1765 18581 1777 18615
rect 1811 18612 1823 18615
rect 6886 18612 6914 18652
rect 33410 18640 33416 18652
rect 33468 18640 33474 18692
rect 40313 18683 40371 18689
rect 40313 18649 40325 18683
rect 40359 18680 40371 18683
rect 47854 18680 47860 18692
rect 40359 18652 47860 18680
rect 40359 18649 40371 18652
rect 40313 18643 40371 18649
rect 47854 18640 47860 18652
rect 47912 18640 47918 18692
rect 1811 18584 6914 18612
rect 19981 18615 20039 18621
rect 1811 18581 1823 18584
rect 1765 18575 1823 18581
rect 19981 18581 19993 18615
rect 20027 18612 20039 18615
rect 21910 18612 21916 18624
rect 20027 18584 21916 18612
rect 20027 18581 20039 18584
rect 19981 18575 20039 18581
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 1578 18232 1584 18284
rect 1636 18232 1642 18284
rect 47026 18232 47032 18284
rect 47084 18272 47090 18284
rect 47949 18275 48007 18281
rect 47949 18272 47961 18275
rect 47084 18244 47961 18272
rect 47084 18232 47090 18244
rect 47949 18241 47961 18244
rect 47995 18241 48007 18275
rect 47949 18235 48007 18241
rect 49142 18164 49148 18216
rect 49200 18164 49206 18216
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 26694 18068 26700 18080
rect 1811 18040 26700 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 26694 18028 26700 18040
rect 26752 18028 26758 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 29178 17620 29184 17672
rect 29236 17660 29242 17672
rect 38013 17663 38071 17669
rect 38013 17660 38025 17663
rect 29236 17632 38025 17660
rect 29236 17620 29242 17632
rect 38013 17629 38025 17632
rect 38059 17629 38071 17663
rect 38013 17623 38071 17629
rect 38197 17595 38255 17601
rect 38197 17561 38209 17595
rect 38243 17592 38255 17595
rect 43346 17592 43352 17604
rect 38243 17564 43352 17592
rect 38243 17561 38255 17564
rect 38197 17555 38255 17561
rect 43346 17552 43352 17564
rect 43404 17552 43410 17604
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 992 17156 1685 17184
rect 992 17144 998 17156
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 2038 17144 2044 17196
rect 2096 17144 2102 17196
rect 27706 17144 27712 17196
rect 27764 17184 27770 17196
rect 38105 17187 38163 17193
rect 38105 17184 38117 17187
rect 27764 17156 38117 17184
rect 27764 17144 27770 17156
rect 38105 17153 38117 17156
rect 38151 17153 38163 17187
rect 38105 17147 38163 17153
rect 42794 17144 42800 17196
rect 42852 17184 42858 17196
rect 47949 17187 48007 17193
rect 47949 17184 47961 17187
rect 42852 17156 47961 17184
rect 42852 17144 42858 17156
rect 47949 17153 47961 17156
rect 47995 17153 48007 17187
rect 47949 17147 48007 17153
rect 49142 17076 49148 17128
rect 49200 17076 49206 17128
rect 38286 17008 38292 17060
rect 38344 17008 38350 17060
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 18322 16640 18328 16652
rect 1903 16612 18328 16640
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 38105 16643 38163 16649
rect 38105 16609 38117 16643
rect 38151 16640 38163 16643
rect 38562 16640 38568 16652
rect 38151 16612 38568 16640
rect 38151 16609 38163 16612
rect 38105 16603 38163 16609
rect 38562 16600 38568 16612
rect 38620 16600 38626 16652
rect 44361 16643 44419 16649
rect 44361 16609 44373 16643
rect 44407 16640 44419 16643
rect 46198 16640 46204 16652
rect 44407 16612 46204 16640
rect 44407 16609 44419 16612
rect 44361 16603 44419 16609
rect 46198 16600 46204 16612
rect 46256 16600 46262 16652
rect 43438 16532 43444 16584
rect 43496 16572 43502 16584
rect 44177 16575 44235 16581
rect 44177 16572 44189 16575
rect 43496 16544 44189 16572
rect 43496 16532 43502 16544
rect 44177 16541 44189 16544
rect 44223 16541 44235 16575
rect 44177 16535 44235 16541
rect 47762 16532 47768 16584
rect 47820 16572 47826 16584
rect 47949 16575 48007 16581
rect 47949 16572 47961 16575
rect 47820 16544 47961 16572
rect 47820 16532 47826 16544
rect 47949 16541 47961 16544
rect 47995 16541 48007 16575
rect 47949 16535 48007 16541
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1673 16507 1731 16513
rect 1673 16504 1685 16507
rect 992 16476 1685 16504
rect 992 16464 998 16476
rect 1673 16473 1685 16476
rect 1719 16473 1731 16507
rect 1673 16467 1731 16473
rect 21818 16464 21824 16516
rect 21876 16504 21882 16516
rect 37921 16507 37979 16513
rect 37921 16504 37933 16507
rect 21876 16476 37933 16504
rect 21876 16464 21882 16476
rect 37921 16473 37933 16476
rect 37967 16473 37979 16507
rect 37921 16467 37979 16473
rect 49142 16464 49148 16516
rect 49200 16464 49206 16516
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 23566 16124 23572 16176
rect 23624 16164 23630 16176
rect 24949 16167 25007 16173
rect 24949 16164 24961 16167
rect 23624 16136 24961 16164
rect 23624 16124 23630 16136
rect 24949 16133 24961 16136
rect 24995 16133 25007 16167
rect 24949 16127 25007 16133
rect 38197 16099 38255 16105
rect 38197 16096 38209 16099
rect 26206 16068 38209 16096
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 25225 16031 25283 16037
rect 25225 15997 25237 16031
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 22830 15920 22836 15972
rect 22888 15960 22894 15972
rect 25240 15960 25268 15991
rect 22888 15932 25268 15960
rect 22888 15920 22894 15932
rect 18966 15852 18972 15904
rect 19024 15892 19030 15904
rect 26206 15892 26234 16068
rect 38197 16065 38209 16068
rect 38243 16096 38255 16099
rect 38841 16099 38899 16105
rect 38841 16096 38853 16099
rect 38243 16068 38853 16096
rect 38243 16065 38255 16068
rect 38197 16059 38255 16065
rect 38841 16065 38853 16068
rect 38887 16065 38899 16099
rect 38841 16059 38899 16065
rect 38381 15963 38439 15969
rect 38381 15929 38393 15963
rect 38427 15960 38439 15963
rect 38470 15960 38476 15972
rect 38427 15932 38476 15960
rect 38427 15929 38439 15932
rect 38381 15923 38439 15929
rect 38470 15920 38476 15932
rect 38528 15920 38534 15972
rect 19024 15864 26234 15892
rect 19024 15852 19030 15864
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 25590 15512 25596 15564
rect 25648 15552 25654 15564
rect 26697 15555 26755 15561
rect 26697 15552 26709 15555
rect 25648 15524 26709 15552
rect 25648 15512 25654 15524
rect 26697 15521 26709 15524
rect 26743 15521 26755 15555
rect 26697 15515 26755 15521
rect 26234 15444 26240 15496
rect 26292 15444 26298 15496
rect 44818 15444 44824 15496
rect 44876 15484 44882 15496
rect 47949 15487 48007 15493
rect 47949 15484 47961 15487
rect 44876 15456 47961 15484
rect 44876 15444 44882 15456
rect 47949 15453 47961 15456
rect 47995 15453 48007 15487
rect 47949 15447 48007 15453
rect 49142 15444 49148 15496
rect 49200 15444 49206 15496
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 1673 15419 1731 15425
rect 1673 15416 1685 15419
rect 992 15388 1685 15416
rect 992 15376 998 15388
rect 1673 15385 1685 15388
rect 1719 15385 1731 15419
rect 1673 15379 1731 15385
rect 24670 15376 24676 15428
rect 24728 15416 24734 15428
rect 26421 15419 26479 15425
rect 26421 15416 26433 15419
rect 24728 15388 26433 15416
rect 24728 15376 24734 15388
rect 26421 15385 26433 15388
rect 26467 15385 26479 15419
rect 26421 15379 26479 15385
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 15838 15348 15844 15360
rect 1995 15320 15844 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 15838 15308 15844 15320
rect 15896 15308 15902 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 22646 15104 22652 15156
rect 22704 15144 22710 15156
rect 22704 15116 29408 15144
rect 22704 15104 22710 15116
rect 25498 15036 25504 15088
rect 25556 15076 25562 15088
rect 28169 15079 28227 15085
rect 28169 15076 28181 15079
rect 25556 15048 28181 15076
rect 25556 15036 25562 15048
rect 28169 15045 28181 15048
rect 28215 15045 28227 15079
rect 28169 15039 28227 15045
rect 934 14968 940 15020
rect 992 15008 998 15020
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 992 14980 1685 15008
rect 992 14968 998 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 27985 14943 28043 14949
rect 27985 14909 27997 14943
rect 28031 14940 28043 14943
rect 28350 14940 28356 14952
rect 28031 14912 28356 14940
rect 28031 14909 28043 14912
rect 27985 14903 28043 14909
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 29380 14949 29408 15116
rect 36722 15036 36728 15088
rect 36780 15076 36786 15088
rect 43717 15079 43775 15085
rect 43717 15076 43729 15079
rect 36780 15048 43729 15076
rect 36780 15036 36786 15048
rect 43717 15045 43729 15048
rect 43763 15045 43775 15079
rect 43717 15039 43775 15045
rect 44266 14968 44272 15020
rect 44324 15008 44330 15020
rect 47949 15011 48007 15017
rect 47949 15008 47961 15011
rect 44324 14980 47961 15008
rect 44324 14968 44330 14980
rect 47949 14977 47961 14980
rect 47995 14977 48007 15011
rect 47949 14971 48007 14977
rect 29365 14943 29423 14949
rect 29365 14909 29377 14943
rect 29411 14909 29423 14943
rect 29365 14903 29423 14909
rect 49142 14900 49148 14952
rect 49200 14900 49206 14952
rect 1949 14807 2007 14813
rect 1949 14773 1961 14807
rect 1995 14804 2007 14807
rect 21542 14804 21548 14816
rect 1995 14776 21548 14804
rect 1995 14773 2007 14776
rect 1949 14767 2007 14773
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 43806 14764 43812 14816
rect 43864 14764 43870 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 30374 14424 30380 14476
rect 30432 14424 30438 14476
rect 29822 14356 29828 14408
rect 29880 14356 29886 14408
rect 27154 14288 27160 14340
rect 27212 14328 27218 14340
rect 30009 14331 30067 14337
rect 30009 14328 30021 14331
rect 27212 14300 30021 14328
rect 27212 14288 27218 14300
rect 30009 14297 30021 14300
rect 30055 14297 30067 14331
rect 30009 14291 30067 14297
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 934 13880 940 13932
rect 992 13920 998 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 992 13892 1593 13920
rect 992 13880 998 13892
rect 1581 13889 1593 13892
rect 1627 13889 1639 13923
rect 1581 13883 1639 13889
rect 28626 13880 28632 13932
rect 28684 13920 28690 13932
rect 37553 13923 37611 13929
rect 37553 13920 37565 13923
rect 28684 13892 37565 13920
rect 28684 13880 28690 13892
rect 37553 13889 37565 13892
rect 37599 13889 37611 13923
rect 37553 13883 37611 13889
rect 47854 13880 47860 13932
rect 47912 13920 47918 13932
rect 47949 13923 48007 13929
rect 47949 13920 47961 13923
rect 47912 13892 47961 13920
rect 47912 13880 47918 13892
rect 47949 13889 47961 13892
rect 47995 13889 48007 13923
rect 47949 13883 48007 13889
rect 29178 13852 29184 13864
rect 1780 13824 29184 13852
rect 1780 13793 1808 13824
rect 29178 13812 29184 13824
rect 29236 13812 29242 13864
rect 37734 13812 37740 13864
rect 37792 13812 37798 13864
rect 49142 13812 49148 13864
rect 49200 13812 49206 13864
rect 1765 13787 1823 13793
rect 1765 13753 1777 13787
rect 1811 13753 1823 13787
rect 1765 13747 1823 13753
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 1854 13336 1860 13388
rect 1912 13336 1918 13388
rect 15654 13336 15660 13388
rect 15712 13376 15718 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 15712 13348 18245 13376
rect 15712 13336 15718 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 992 13280 1593 13308
rect 992 13268 998 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 18414 13268 18420 13320
rect 18472 13268 18478 13320
rect 31018 13268 31024 13320
rect 31076 13308 31082 13320
rect 37645 13311 37703 13317
rect 37645 13308 37657 13311
rect 31076 13280 37657 13308
rect 31076 13268 31082 13280
rect 37645 13277 37657 13280
rect 37691 13277 37703 13311
rect 37645 13271 37703 13277
rect 43346 13268 43352 13320
rect 43404 13308 43410 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 43404 13280 47961 13308
rect 43404 13268 43410 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 37829 13243 37887 13249
rect 37829 13209 37841 13243
rect 37875 13240 37887 13243
rect 38562 13240 38568 13252
rect 37875 13212 38568 13240
rect 37875 13209 37887 13212
rect 37829 13203 37887 13209
rect 38562 13200 38568 13212
rect 38620 13200 38626 13252
rect 49142 13200 49148 13252
rect 49200 13200 49206 13252
rect 18877 13175 18935 13181
rect 18877 13141 18889 13175
rect 18923 13172 18935 13175
rect 19518 13172 19524 13184
rect 18923 13144 19524 13172
rect 18923 13141 18935 13144
rect 18877 13135 18935 13141
rect 19518 13132 19524 13144
rect 19576 13132 19582 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 23566 12977 23572 12980
rect 23523 12971 23572 12977
rect 23523 12937 23535 12971
rect 23569 12937 23572 12971
rect 23523 12931 23572 12937
rect 23566 12928 23572 12931
rect 23624 12928 23630 12980
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 23452 12835 23510 12841
rect 23452 12832 23464 12835
rect 18472 12804 23464 12832
rect 18472 12792 18478 12804
rect 23452 12801 23464 12804
rect 23498 12832 23510 12835
rect 24854 12832 24860 12844
rect 23498 12804 24860 12832
rect 23498 12801 23510 12804
rect 23452 12795 23510 12801
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 38289 12835 38347 12841
rect 38289 12832 38301 12835
rect 26206 12804 38301 12832
rect 20070 12724 20076 12776
rect 20128 12764 20134 12776
rect 26206 12764 26234 12804
rect 38289 12801 38301 12804
rect 38335 12801 38347 12835
rect 38289 12795 38347 12801
rect 20128 12736 26234 12764
rect 20128 12724 20134 12736
rect 38378 12588 38384 12640
rect 38436 12588 38442 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 24670 12384 24676 12436
rect 24728 12433 24734 12436
rect 25498 12433 25504 12436
rect 24728 12427 24777 12433
rect 24728 12393 24731 12427
rect 24765 12393 24777 12427
rect 24728 12387 24777 12393
rect 25455 12427 25504 12433
rect 25455 12393 25467 12427
rect 25501 12393 25504 12427
rect 25455 12387 25504 12393
rect 24728 12384 24734 12387
rect 25498 12384 25504 12387
rect 25556 12384 25562 12436
rect 26743 12427 26801 12433
rect 26743 12393 26755 12427
rect 26789 12424 26801 12427
rect 27154 12424 27160 12436
rect 26789 12396 27160 12424
rect 26789 12393 26801 12396
rect 26743 12387 26801 12393
rect 27154 12384 27160 12396
rect 27212 12384 27218 12436
rect 27522 12288 27528 12300
rect 24596 12260 27528 12288
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 24596 12229 24624 12260
rect 27522 12248 27528 12260
rect 27580 12248 27586 12300
rect 24596 12223 24674 12229
rect 24596 12220 24628 12223
rect 20220 12192 24628 12220
rect 20220 12180 20226 12192
rect 24616 12189 24628 12192
rect 24662 12189 24674 12223
rect 24616 12183 24674 12189
rect 25314 12180 25320 12232
rect 25372 12229 25378 12232
rect 25372 12223 25410 12229
rect 25398 12189 25410 12223
rect 25372 12183 25410 12189
rect 25372 12180 25378 12183
rect 25498 12180 25504 12232
rect 25556 12220 25562 12232
rect 26640 12223 26698 12229
rect 26640 12220 26652 12223
rect 25556 12192 26652 12220
rect 25556 12180 25562 12192
rect 26640 12189 26652 12192
rect 26686 12189 26698 12223
rect 26640 12183 26698 12189
rect 46934 12180 46940 12232
rect 46992 12220 46998 12232
rect 47949 12223 48007 12229
rect 47949 12220 47961 12223
rect 46992 12192 47961 12220
rect 46992 12180 46998 12192
rect 47949 12189 47961 12192
rect 47995 12189 48007 12223
rect 47949 12183 48007 12189
rect 49142 12180 49148 12232
rect 49200 12180 49206 12232
rect 934 12112 940 12164
rect 992 12152 998 12164
rect 1673 12155 1731 12161
rect 1673 12152 1685 12155
rect 992 12124 1685 12152
rect 992 12112 998 12124
rect 1673 12121 1685 12124
rect 1719 12121 1731 12155
rect 1673 12115 1731 12121
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 17494 12084 17500 12096
rect 1995 12056 17500 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 992 11716 1685 11744
rect 992 11704 998 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 19978 11704 19984 11756
rect 20036 11704 20042 11756
rect 37826 11704 37832 11756
rect 37884 11744 37890 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 37884 11716 47961 11744
rect 37884 11704 37890 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 18598 11636 18604 11688
rect 18656 11676 18662 11688
rect 20162 11676 20168 11688
rect 18656 11648 20168 11676
rect 18656 11636 18662 11648
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 49142 11636 49148 11688
rect 49200 11636 49206 11688
rect 1949 11611 2007 11617
rect 1949 11577 1961 11611
rect 1995 11608 2007 11611
rect 21818 11608 21824 11620
rect 1995 11580 21824 11608
rect 1995 11577 2007 11580
rect 1949 11571 2007 11577
rect 21818 11568 21824 11580
rect 21876 11568 21882 11620
rect 20625 11543 20683 11549
rect 20625 11509 20637 11543
rect 20671 11540 20683 11543
rect 21358 11540 21364 11552
rect 20671 11512 21364 11540
rect 20671 11509 20683 11512
rect 20625 11503 20683 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17368 11308 26234 11336
rect 17368 11296 17374 11308
rect 25314 11268 25320 11280
rect 22112 11240 25320 11268
rect 21910 11160 21916 11212
rect 21968 11160 21974 11212
rect 22112 11209 22140 11240
rect 25314 11228 25320 11240
rect 25372 11228 25378 11280
rect 26206 11268 26234 11308
rect 36725 11271 36783 11277
rect 36725 11268 36737 11271
rect 26206 11240 36737 11268
rect 36725 11237 36737 11240
rect 36771 11237 36783 11271
rect 36725 11231 36783 11237
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11169 22155 11203
rect 22097 11163 22155 11169
rect 22186 11160 22192 11212
rect 22244 11200 22250 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 22244 11172 24593 11200
rect 22244 11160 22250 11172
rect 24581 11169 24593 11172
rect 24627 11169 24639 11203
rect 24581 11163 24639 11169
rect 24765 11203 24823 11209
rect 24765 11169 24777 11203
rect 24811 11200 24823 11203
rect 25498 11200 25504 11212
rect 24811 11172 25504 11200
rect 24811 11169 24823 11172
rect 24765 11163 24823 11169
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 24780 11132 24808 11163
rect 25498 11160 25504 11172
rect 25556 11160 25562 11212
rect 23440 11104 24808 11132
rect 36740 11132 36768 11231
rect 37369 11135 37427 11141
rect 37369 11132 37381 11135
rect 36740 11104 37381 11132
rect 23440 11092 23446 11104
rect 37369 11101 37381 11104
rect 37415 11101 37427 11135
rect 37369 11095 37427 11101
rect 22557 11067 22615 11073
rect 22557 11033 22569 11067
rect 22603 11064 22615 11067
rect 24578 11064 24584 11076
rect 22603 11036 24584 11064
rect 22603 11033 22615 11036
rect 22557 11027 22615 11033
rect 24578 11024 24584 11036
rect 24636 11024 24642 11076
rect 25225 11067 25283 11073
rect 25225 11033 25237 11067
rect 25271 11064 25283 11067
rect 26602 11064 26608 11076
rect 25271 11036 26608 11064
rect 25271 11033 25283 11036
rect 25225 11027 25283 11033
rect 26602 11024 26608 11036
rect 26660 11024 26666 11076
rect 37458 11024 37464 11076
rect 37516 11064 37522 11076
rect 37553 11067 37611 11073
rect 37553 11064 37565 11067
rect 37516 11036 37565 11064
rect 37516 11024 37522 11036
rect 37553 11033 37565 11036
rect 37599 11033 37611 11067
rect 37553 11027 37611 11033
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 992 10628 1685 10656
rect 992 10616 998 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 37553 10659 37611 10665
rect 37553 10656 37565 10659
rect 1673 10619 1731 10625
rect 26206 10628 37565 10656
rect 15838 10480 15844 10532
rect 15896 10520 15902 10532
rect 16390 10520 16396 10532
rect 15896 10492 16396 10520
rect 15896 10480 15902 10492
rect 16390 10480 16396 10492
rect 16448 10520 16454 10532
rect 26206 10520 26234 10628
rect 37553 10625 37565 10628
rect 37599 10656 37611 10659
rect 38197 10659 38255 10665
rect 38197 10656 38209 10659
rect 37599 10628 38209 10656
rect 37599 10625 37611 10628
rect 37553 10619 37611 10625
rect 38197 10625 38209 10628
rect 38243 10625 38255 10659
rect 38197 10619 38255 10625
rect 38286 10616 38292 10668
rect 38344 10656 38350 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 38344 10628 47961 10656
rect 38344 10616 38350 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 49142 10548 49148 10600
rect 49200 10548 49206 10600
rect 16448 10492 26234 10520
rect 37737 10523 37795 10529
rect 16448 10480 16454 10492
rect 37737 10489 37749 10523
rect 37783 10520 37795 10523
rect 37826 10520 37832 10532
rect 37783 10492 37832 10520
rect 37783 10489 37795 10492
rect 37737 10483 37795 10489
rect 37826 10480 37832 10492
rect 37884 10480 37890 10532
rect 1949 10455 2007 10461
rect 1949 10421 1961 10455
rect 1995 10452 2007 10455
rect 18966 10452 18972 10464
rect 1995 10424 18972 10452
rect 1995 10421 2007 10424
rect 1949 10415 2007 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10112 26111 10115
rect 27062 10112 27068 10124
rect 26099 10084 27068 10112
rect 26099 10081 26111 10084
rect 26053 10075 26111 10081
rect 27062 10072 27068 10084
rect 27120 10072 27126 10124
rect 38470 10004 38476 10056
rect 38528 10044 38534 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 38528 10016 47961 10044
rect 38528 10004 38534 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 934 9936 940 9988
rect 992 9976 998 9988
rect 1673 9979 1731 9985
rect 1673 9976 1685 9979
rect 992 9948 1685 9976
rect 992 9936 998 9948
rect 1673 9945 1685 9948
rect 1719 9945 1731 9979
rect 1673 9939 1731 9945
rect 25406 9936 25412 9988
rect 25464 9976 25470 9988
rect 26329 9979 26387 9985
rect 26329 9976 26341 9979
rect 25464 9948 26341 9976
rect 25464 9936 25470 9948
rect 26329 9945 26341 9948
rect 26375 9945 26387 9979
rect 33318 9976 33324 9988
rect 27554 9948 33324 9976
rect 26329 9939 26387 9945
rect 1765 9911 1823 9917
rect 1765 9877 1777 9911
rect 1811 9908 1823 9911
rect 14642 9908 14648 9920
rect 1811 9880 14648 9908
rect 1811 9877 1823 9880
rect 1765 9871 1823 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 27632 9908 27660 9948
rect 33318 9936 33324 9948
rect 33376 9936 33382 9988
rect 49142 9936 49148 9988
rect 49200 9936 49206 9988
rect 22428 9880 27660 9908
rect 22428 9868 22434 9880
rect 27798 9868 27804 9920
rect 27856 9868 27862 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 22428 9608 22770 9636
rect 22428 9596 22434 9608
rect 20254 9528 20260 9580
rect 20312 9568 20318 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 20312 9540 22017 9568
rect 20312 9528 20318 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 25222 9528 25228 9580
rect 25280 9568 25286 9580
rect 36265 9571 36323 9577
rect 36265 9568 36277 9571
rect 25280 9540 36277 9568
rect 25280 9528 25286 9540
rect 36265 9537 36277 9540
rect 36311 9537 36323 9571
rect 36265 9531 36323 9537
rect 22278 9460 22284 9512
rect 22336 9460 22342 9512
rect 36446 9392 36452 9444
rect 36504 9392 36510 9444
rect 23753 9367 23811 9373
rect 23753 9333 23765 9367
rect 23799 9364 23811 9367
rect 25406 9364 25412 9376
rect 23799 9336 25412 9364
rect 23799 9333 23811 9336
rect 23753 9327 23811 9333
rect 25406 9324 25412 9336
rect 25464 9324 25470 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 992 8928 1593 8956
rect 992 8916 998 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 46198 8916 46204 8968
rect 46256 8956 46262 8968
rect 47949 8959 48007 8965
rect 47949 8956 47961 8959
rect 46256 8928 47961 8956
rect 46256 8916 46262 8928
rect 47949 8925 47961 8928
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 49142 8916 49148 8968
rect 49200 8916 49206 8968
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8820 1823 8823
rect 28626 8820 28632 8832
rect 1811 8792 28632 8820
rect 1811 8789 1823 8792
rect 1765 8783 1823 8789
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 25314 8576 25320 8628
rect 25372 8616 25378 8628
rect 25590 8616 25596 8628
rect 25372 8588 25596 8616
rect 25372 8576 25378 8588
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 30742 8616 30748 8628
rect 27632 8588 30748 8616
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 24670 8440 24676 8492
rect 24728 8480 24734 8492
rect 25133 8483 25191 8489
rect 25133 8480 25145 8483
rect 24728 8452 25145 8480
rect 24728 8440 24734 8452
rect 25133 8449 25145 8452
rect 25179 8480 25191 8483
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 25179 8452 27169 8480
rect 25179 8449 25191 8452
rect 25133 8443 25191 8449
rect 27157 8449 27169 8452
rect 27203 8480 27215 8483
rect 27632 8480 27660 8588
rect 30742 8576 30748 8588
rect 30800 8576 30806 8628
rect 33318 8576 33324 8628
rect 33376 8576 33382 8628
rect 33336 8548 33364 8576
rect 33336 8520 33442 8548
rect 31018 8480 31024 8492
rect 27203 8452 27660 8480
rect 27724 8452 31024 8480
rect 27203 8449 27215 8452
rect 27157 8443 27215 8449
rect 27724 8412 27752 8452
rect 31018 8440 31024 8452
rect 31076 8440 31082 8492
rect 32674 8440 32680 8492
rect 32732 8440 32738 8492
rect 37734 8440 37740 8492
rect 37792 8480 37798 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 37792 8452 47961 8480
rect 37792 8440 37798 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 26206 8384 27752 8412
rect 1765 8347 1823 8353
rect 1765 8313 1777 8347
rect 1811 8344 1823 8347
rect 26206 8344 26234 8384
rect 27798 8372 27804 8424
rect 27856 8412 27862 8424
rect 32953 8415 33011 8421
rect 32953 8412 32965 8415
rect 27856 8384 32965 8412
rect 27856 8372 27862 8384
rect 32953 8381 32965 8384
rect 32999 8381 33011 8415
rect 32953 8375 33011 8381
rect 49142 8372 49148 8424
rect 49200 8372 49206 8424
rect 27816 8344 27844 8372
rect 1811 8316 26234 8344
rect 27540 8316 27844 8344
rect 1811 8313 1823 8316
rect 1765 8307 1823 8313
rect 25406 8236 25412 8288
rect 25464 8236 25470 8288
rect 27433 8279 27491 8285
rect 27433 8245 27445 8279
rect 27479 8276 27491 8279
rect 27540 8276 27568 8316
rect 27479 8248 27568 8276
rect 27479 8245 27491 8248
rect 27433 8239 27491 8245
rect 27614 8236 27620 8288
rect 27672 8236 27678 8288
rect 34422 8236 34428 8288
rect 34480 8236 34486 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 22278 8032 22284 8084
rect 22336 8072 22342 8084
rect 23017 8075 23075 8081
rect 23017 8072 23029 8075
rect 22336 8044 23029 8072
rect 22336 8032 22342 8044
rect 23017 8041 23029 8044
rect 23063 8041 23075 8075
rect 23017 8035 23075 8041
rect 23382 8032 23388 8084
rect 23440 8032 23446 8084
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7868 22983 7871
rect 24670 7868 24676 7880
rect 22971 7840 24676 7868
rect 22971 7837 22983 7840
rect 22925 7831 22983 7837
rect 24670 7828 24676 7840
rect 24728 7828 24734 7880
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 992 7364 1685 7392
rect 992 7352 998 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 30742 7352 30748 7404
rect 30800 7352 30806 7404
rect 38562 7352 38568 7404
rect 38620 7392 38626 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 38620 7364 47961 7392
rect 38620 7352 38626 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 49142 7284 49148 7336
rect 49200 7284 49206 7336
rect 18414 7216 18420 7268
rect 18472 7256 18478 7268
rect 24854 7256 24860 7268
rect 18472 7228 24860 7256
rect 18472 7216 18478 7228
rect 24854 7216 24860 7228
rect 24912 7256 24918 7268
rect 31205 7259 31263 7265
rect 31205 7256 31217 7259
rect 24912 7228 31217 7256
rect 24912 7216 24918 7228
rect 31205 7225 31217 7228
rect 31251 7225 31263 7259
rect 31205 7219 31263 7225
rect 1949 7191 2007 7197
rect 1949 7157 1961 7191
rect 1995 7188 2007 7191
rect 20070 7188 20076 7200
rect 1995 7160 20076 7188
rect 1995 7157 2007 7160
rect 1949 7151 2007 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 30285 7191 30343 7197
rect 30285 7157 30297 7191
rect 30331 7188 30343 7191
rect 31021 7191 31079 7197
rect 31021 7188 31033 7191
rect 30331 7160 31033 7188
rect 30331 7157 30343 7160
rect 30285 7151 30343 7157
rect 31021 7157 31033 7160
rect 31067 7188 31079 7191
rect 34422 7188 34428 7200
rect 31067 7160 34428 7188
rect 31067 7157 31079 7160
rect 31021 7151 31079 7157
rect 34422 7148 34428 7160
rect 34480 7148 34486 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 19518 6740 19524 6792
rect 19576 6740 19582 6792
rect 38378 6740 38384 6792
rect 38436 6780 38442 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 38436 6752 47961 6780
rect 38436 6740 38442 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 992 6684 1685 6712
rect 992 6672 998 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 1673 6675 1731 6681
rect 49142 6672 49148 6724
rect 49200 6672 49206 6724
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 16942 6644 16948 6656
rect 1811 6616 16948 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 19610 6604 19616 6656
rect 19668 6604 19674 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 12989 5831 13047 5837
rect 12989 5797 13001 5831
rect 13035 5828 13047 5831
rect 22278 5828 22284 5840
rect 13035 5800 22284 5828
rect 13035 5797 13047 5800
rect 12989 5791 13047 5797
rect 22278 5788 22284 5800
rect 22336 5788 22342 5840
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5760 11299 5763
rect 14090 5760 14096 5772
rect 11287 5732 14096 5760
rect 11287 5729 11299 5732
rect 11241 5723 11299 5729
rect 14090 5720 14096 5732
rect 14148 5720 14154 5772
rect 21358 5652 21364 5704
rect 21416 5652 21422 5704
rect 22370 5692 22376 5704
rect 21468 5664 22376 5692
rect 934 5584 940 5636
rect 992 5624 998 5636
rect 1673 5627 1731 5633
rect 1673 5624 1685 5627
rect 992 5596 1685 5624
rect 992 5584 998 5596
rect 1673 5593 1685 5596
rect 1719 5593 1731 5627
rect 1673 5587 1731 5593
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 11517 5627 11575 5633
rect 11517 5624 11529 5627
rect 9732 5596 11529 5624
rect 9732 5584 9738 5596
rect 11517 5593 11529 5596
rect 11563 5593 11575 5627
rect 21468 5624 21496 5664
rect 22370 5652 22376 5664
rect 22428 5652 22434 5704
rect 24670 5652 24676 5704
rect 24728 5652 24734 5704
rect 26602 5652 26608 5704
rect 26660 5652 26666 5704
rect 43806 5652 43812 5704
rect 43864 5692 43870 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 43864 5664 47961 5692
rect 43864 5652 43870 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 49142 5652 49148 5704
rect 49200 5652 49206 5704
rect 12742 5596 21496 5624
rect 21545 5627 21603 5633
rect 11517 5587 11575 5593
rect 21545 5593 21557 5627
rect 21591 5624 21603 5627
rect 22186 5624 22192 5636
rect 21591 5596 22192 5624
rect 21591 5593 21603 5596
rect 21545 5587 21603 5593
rect 22186 5584 22192 5596
rect 22244 5584 22250 5636
rect 24857 5627 24915 5633
rect 24857 5593 24869 5627
rect 24903 5624 24915 5627
rect 25222 5624 25228 5636
rect 24903 5596 25228 5624
rect 24903 5593 24915 5596
rect 24857 5587 24915 5593
rect 25222 5584 25228 5596
rect 25280 5584 25286 5636
rect 26789 5627 26847 5633
rect 26789 5593 26801 5627
rect 26835 5624 26847 5627
rect 28810 5624 28816 5636
rect 26835 5596 28816 5624
rect 26835 5593 26847 5596
rect 26789 5587 26847 5593
rect 28810 5584 28816 5596
rect 28868 5584 28874 5636
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 17218 5556 17224 5568
rect 1995 5528 17224 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 13541 5287 13599 5293
rect 13541 5253 13553 5287
rect 13587 5284 13599 5287
rect 18414 5284 18420 5296
rect 13587 5256 18420 5284
rect 13587 5253 13599 5256
rect 13541 5247 13599 5253
rect 18414 5244 18420 5256
rect 18472 5244 18478 5296
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 992 5188 1685 5216
rect 992 5176 998 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 37458 5176 37464 5228
rect 37516 5216 37522 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 37516 5188 47961 5216
rect 37516 5176 37522 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 49142 5108 49148 5160
rect 49200 5108 49206 5160
rect 15838 5080 15844 5092
rect 6886 5052 15844 5080
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 6886 5012 6914 5052
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 1995 4984 6914 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 13630 4972 13636 5024
rect 13688 4972 13694 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 17589 4675 17647 4681
rect 17589 4672 17601 4675
rect 14240 4644 17601 4672
rect 14240 4632 14246 4644
rect 17589 4641 17601 4644
rect 17635 4641 17647 4675
rect 17589 4635 17647 4641
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 18598 4604 18604 4616
rect 15335 4576 18604 4604
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4604 19579 4607
rect 23382 4604 23388 4616
rect 19567 4576 23388 4604
rect 19567 4573 19579 4576
rect 19521 4567 19579 4573
rect 23382 4564 23388 4576
rect 23440 4564 23446 4616
rect 17405 4539 17463 4545
rect 17405 4505 17417 4539
rect 17451 4536 17463 4539
rect 25590 4536 25596 4548
rect 17451 4508 25596 4536
rect 17451 4505 17463 4508
rect 17405 4499 17463 4505
rect 25590 4496 25596 4508
rect 25648 4496 25654 4548
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 15381 4471 15439 4477
rect 15381 4468 15393 4471
rect 11112 4440 15393 4468
rect 11112 4428 11118 4440
rect 15381 4437 15393 4440
rect 15427 4437 15439 4471
rect 15381 4431 15439 4437
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 19613 4471 19671 4477
rect 19613 4468 19625 4471
rect 17920 4440 19625 4468
rect 17920 4428 17926 4440
rect 19613 4437 19625 4440
rect 19659 4437 19671 4471
rect 19613 4431 19671 4437
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 992 4100 1593 4128
rect 992 4088 998 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 37826 4088 37832 4140
rect 37884 4128 37890 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 37884 4100 47961 4128
rect 37884 4088 37890 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49142 4020 49148 4072
rect 49200 4020 49206 4072
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 25314 3924 25320 3936
rect 1811 3896 25320 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 36446 3476 36452 3528
rect 36504 3516 36510 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 36504 3488 47961 3516
rect 36504 3476 36510 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1673 3451 1731 3457
rect 1673 3448 1685 3451
rect 992 3420 1685 3448
rect 992 3408 998 3420
rect 1673 3417 1685 3420
rect 1719 3417 1731 3451
rect 1673 3411 1731 3417
rect 25866 3408 25872 3460
rect 25924 3448 25930 3460
rect 48590 3448 48596 3460
rect 25924 3420 48596 3448
rect 25924 3408 25930 3420
rect 48590 3408 48596 3420
rect 48648 3408 48654 3460
rect 49142 3408 49148 3460
rect 49200 3408 49206 3460
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3380 1823 3383
rect 14734 3380 14740 3392
rect 1811 3352 14740 3380
rect 1811 3349 1823 3352
rect 1765 3343 1823 3349
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 28810 3000 28816 3052
rect 28868 3000 28874 3052
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 29273 2975 29331 2981
rect 29273 2972 29285 2975
rect 28776 2944 29285 2972
rect 28776 2932 28782 2944
rect 29273 2941 29285 2944
rect 29319 2941 29331 2975
rect 29273 2935 29331 2941
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 34422 2592 34428 2644
rect 34480 2632 34486 2644
rect 34480 2604 45554 2632
rect 34480 2592 34486 2604
rect 28350 2524 28356 2576
rect 28408 2564 28414 2576
rect 28408 2536 38976 2564
rect 28408 2524 28414 2536
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 5592 2468 7021 2496
rect 5592 2456 5598 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 8904 2468 9689 2496
rect 8904 2456 8910 2468
rect 9677 2465 9689 2468
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12216 2468 12725 2496
rect 12216 2456 12222 2468
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 15470 2456 15476 2508
rect 15528 2456 15534 2508
rect 18782 2456 18788 2508
rect 18840 2496 18846 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 18840 2468 19901 2496
rect 18840 2456 18846 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22649 2499 22707 2505
rect 22649 2496 22661 2499
rect 22152 2468 22661 2496
rect 22152 2456 22158 2468
rect 22649 2465 22661 2468
rect 22695 2465 22707 2499
rect 22649 2459 22707 2465
rect 25406 2456 25412 2508
rect 25464 2496 25470 2508
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25464 2468 25697 2496
rect 25464 2456 25470 2468
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 29822 2456 29828 2508
rect 29880 2496 29886 2508
rect 38948 2505 38976 2536
rect 38933 2499 38991 2505
rect 29880 2468 38884 2496
rect 29880 2456 29886 2468
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2280 2400 2513 2428
rect 2280 2388 2286 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 9309 2431 9367 2437
rect 6779 2400 6914 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 6886 2360 6914 2400
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 11054 2428 11060 2440
rect 9355 2400 11060 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 14182 2428 14188 2440
rect 12391 2400 14188 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2428 15163 2431
rect 17862 2428 17868 2440
rect 15151 2400 17868 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 22186 2388 22192 2440
rect 22244 2388 22250 2440
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 32030 2388 32036 2440
rect 32088 2428 32094 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32088 2400 32505 2428
rect 32088 2388 32094 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32493 2391 32551 2397
rect 35342 2388 35348 2440
rect 35400 2428 35406 2440
rect 35437 2431 35495 2437
rect 35437 2428 35449 2431
rect 35400 2400 35449 2428
rect 35400 2388 35406 2400
rect 35437 2397 35449 2400
rect 35483 2397 35495 2431
rect 35437 2391 35495 2397
rect 35713 2431 35771 2437
rect 35713 2397 35725 2431
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 13630 2360 13636 2372
rect 6886 2332 13636 2360
rect 13630 2320 13636 2332
rect 13688 2320 13694 2372
rect 26234 2320 26240 2372
rect 26292 2360 26298 2372
rect 35728 2360 35756 2391
rect 38654 2388 38660 2440
rect 38712 2388 38718 2440
rect 38856 2428 38884 2468
rect 38933 2465 38945 2499
rect 38979 2465 38991 2499
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 38933 2459 38991 2465
rect 39040 2468 42901 2496
rect 39040 2428 39068 2468
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 38856 2400 39068 2428
rect 41966 2388 41972 2440
rect 42024 2428 42030 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 42024 2400 42625 2428
rect 42024 2388 42030 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 45526 2428 45554 2604
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 45526 2400 47961 2428
rect 42613 2391 42671 2397
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 26292 2332 35756 2360
rect 26292 2320 26298 2332
rect 45278 2320 45284 2372
rect 45336 2360 45342 2372
rect 45465 2363 45523 2369
rect 45465 2360 45477 2363
rect 45336 2332 45477 2360
rect 45336 2320 45342 2332
rect 45465 2329 45477 2332
rect 45511 2329 45523 2363
rect 45465 2323 45523 2329
rect 49142 2320 49148 2372
rect 49200 2320 49206 2372
rect 2317 2295 2375 2301
rect 2317 2261 2329 2295
rect 2363 2292 2375 2295
rect 9674 2292 9680 2304
rect 2363 2264 9680 2292
rect 2363 2261 2375 2264
rect 2317 2255 2375 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 24762 2252 24768 2304
rect 24820 2292 24826 2304
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 24820 2264 32321 2292
rect 24820 2252 24826 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 45554 2252 45560 2304
rect 45612 2252 45618 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 30742 2048 30748 2100
rect 30800 2088 30806 2100
rect 45554 2088 45560 2100
rect 30800 2060 45560 2088
rect 30800 2048 30806 2060
rect 45554 2048 45560 2060
rect 45612 2048 45618 2100
<< via1 >>
rect 30564 54612 30616 54664
rect 37464 54612 37516 54664
rect 32496 54544 32548 54596
rect 45836 54544 45888 54596
rect 34520 54476 34572 54528
rect 40684 54476 40736 54528
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 27950 54374 28002 54426
rect 28014 54374 28066 54426
rect 28078 54374 28130 54426
rect 28142 54374 28194 54426
rect 28206 54374 28258 54426
rect 37950 54374 38002 54426
rect 38014 54374 38066 54426
rect 38078 54374 38130 54426
rect 38142 54374 38194 54426
rect 38206 54374 38258 54426
rect 47950 54374 48002 54426
rect 48014 54374 48066 54426
rect 48078 54374 48130 54426
rect 48142 54374 48194 54426
rect 48206 54374 48258 54426
rect 3516 54204 3568 54256
rect 5540 54204 5592 54256
rect 8668 54204 8720 54256
rect 10600 54204 10652 54256
rect 13820 54204 13872 54256
rect 15752 54204 15804 54256
rect 18972 54204 19024 54256
rect 4896 54136 4948 54188
rect 5448 54111 5500 54120
rect 5448 54077 5457 54111
rect 5457 54077 5491 54111
rect 5491 54077 5500 54111
rect 5448 54068 5500 54077
rect 10508 54136 10560 54188
rect 13728 54136 13780 54188
rect 15016 54179 15068 54188
rect 15016 54145 15025 54179
rect 15025 54145 15059 54179
rect 15059 54145 15068 54179
rect 15016 54136 15068 54145
rect 20720 54204 20772 54256
rect 30104 54272 30156 54324
rect 32220 54272 32272 54324
rect 28264 54204 28316 54256
rect 30196 54204 30248 54256
rect 33692 54204 33744 54256
rect 35256 54204 35308 54256
rect 15384 54068 15436 54120
rect 20260 54068 20312 54120
rect 22836 54136 22888 54188
rect 23480 54136 23532 54188
rect 24124 54136 24176 54188
rect 24768 54136 24820 54188
rect 25412 54136 25464 54188
rect 26240 54136 26292 54188
rect 26700 54136 26752 54188
rect 27436 54136 27488 54188
rect 28356 54136 28408 54188
rect 29276 54136 29328 54188
rect 30288 54136 30340 54188
rect 30656 54136 30708 54188
rect 31852 54136 31904 54188
rect 32588 54136 32640 54188
rect 33232 54136 33284 54188
rect 35072 54136 35124 54188
rect 35900 54136 35952 54188
rect 23572 54068 23624 54120
rect 27712 54068 27764 54120
rect 28816 54068 28868 54120
rect 29736 54068 29788 54120
rect 37188 54204 37240 54256
rect 37004 54136 37056 54188
rect 37740 54136 37792 54188
rect 38384 54136 38436 54188
rect 39120 54204 39172 54256
rect 40776 54204 40828 54256
rect 42156 54204 42208 54256
rect 39580 54136 39632 54188
rect 40316 54136 40368 54188
rect 44732 54136 44784 54188
rect 45836 54272 45888 54324
rect 45652 54204 45704 54256
rect 46112 54136 46164 54188
rect 47308 54136 47360 54188
rect 47860 54136 47912 54188
rect 27896 54000 27948 54052
rect 31944 54000 31996 54052
rect 25412 53932 25464 53984
rect 26056 53932 26108 53984
rect 27436 53932 27488 53984
rect 28356 53932 28408 53984
rect 29092 53932 29144 53984
rect 30380 53975 30432 53984
rect 30380 53941 30389 53975
rect 30389 53941 30423 53975
rect 30423 53941 30432 53975
rect 30380 53932 30432 53941
rect 30748 53932 30800 53984
rect 32312 53975 32364 53984
rect 32312 53941 32321 53975
rect 32321 53941 32355 53975
rect 32355 53941 32364 53975
rect 32312 53932 32364 53941
rect 32588 53932 32640 53984
rect 33600 53975 33652 53984
rect 33600 53941 33609 53975
rect 33609 53941 33643 53975
rect 33643 53941 33652 53975
rect 33600 53932 33652 53941
rect 33692 53932 33744 53984
rect 37464 53975 37516 53984
rect 37464 53941 37473 53975
rect 37473 53941 37507 53975
rect 37507 53941 37516 53975
rect 37464 53932 37516 53941
rect 37556 53932 37608 53984
rect 40684 54043 40736 54052
rect 40684 54009 40693 54043
rect 40693 54009 40727 54043
rect 40727 54009 40736 54043
rect 40684 54000 40736 54009
rect 40776 54000 40828 54052
rect 43904 53975 43956 53984
rect 43904 53941 43913 53975
rect 43913 53941 43947 53975
rect 43947 53941 43956 53975
rect 43904 53932 43956 53941
rect 48688 53975 48740 53984
rect 48688 53941 48697 53975
rect 48697 53941 48731 53975
rect 48731 53941 48740 53975
rect 48688 53932 48740 53941
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 32950 53830 33002 53882
rect 33014 53830 33066 53882
rect 33078 53830 33130 53882
rect 33142 53830 33194 53882
rect 33206 53830 33258 53882
rect 42950 53830 43002 53882
rect 43014 53830 43066 53882
rect 43078 53830 43130 53882
rect 43142 53830 43194 53882
rect 43206 53830 43258 53882
rect 2872 53635 2924 53644
rect 2872 53601 2881 53635
rect 2881 53601 2915 53635
rect 2915 53601 2924 53635
rect 2872 53592 2924 53601
rect 6092 53635 6144 53644
rect 6092 53601 6101 53635
rect 6101 53601 6135 53635
rect 6135 53601 6144 53635
rect 6092 53592 6144 53601
rect 7840 53635 7892 53644
rect 7840 53601 7849 53635
rect 7849 53601 7883 53635
rect 7883 53601 7892 53635
rect 7840 53592 7892 53601
rect 11244 53635 11296 53644
rect 11244 53601 11253 53635
rect 11253 53601 11287 53635
rect 11287 53601 11296 53635
rect 11244 53592 11296 53601
rect 13360 53635 13412 53644
rect 13360 53601 13369 53635
rect 13369 53601 13403 53635
rect 13403 53601 13412 53635
rect 13360 53592 13412 53601
rect 2044 53567 2096 53576
rect 2044 53533 2053 53567
rect 2053 53533 2087 53567
rect 2087 53533 2096 53567
rect 2044 53524 2096 53533
rect 8484 53524 8536 53576
rect 8392 53456 8444 53508
rect 15200 53524 15252 53576
rect 22100 53660 22152 53712
rect 16396 53635 16448 53644
rect 16396 53601 16405 53635
rect 16405 53601 16439 53635
rect 16439 53601 16448 53635
rect 16396 53592 16448 53601
rect 18328 53635 18380 53644
rect 18328 53601 18337 53635
rect 18337 53601 18371 53635
rect 18371 53601 18380 53635
rect 18328 53592 18380 53601
rect 29460 53660 29512 53712
rect 38660 53660 38712 53712
rect 34428 53592 34480 53644
rect 38292 53592 38344 53644
rect 13544 53456 13596 53508
rect 22192 53524 22244 53576
rect 26240 53524 26292 53576
rect 28632 53524 28684 53576
rect 31208 53524 31260 53576
rect 33784 53524 33836 53576
rect 20904 53456 20956 53508
rect 29644 53456 29696 53508
rect 36360 53524 36412 53576
rect 38936 53524 38988 53576
rect 44088 53524 44140 53576
rect 46664 53524 46716 53576
rect 48320 53524 48372 53576
rect 48596 53524 48648 53576
rect 37372 53456 37424 53508
rect 22652 53388 22704 53440
rect 23388 53388 23440 53440
rect 28632 53388 28684 53440
rect 30472 53388 30524 53440
rect 31760 53388 31812 53440
rect 39028 53431 39080 53440
rect 39028 53397 39037 53431
rect 39037 53397 39071 53431
rect 39071 53397 39080 53431
rect 39028 53388 39080 53397
rect 48872 53431 48924 53440
rect 48872 53397 48881 53431
rect 48881 53397 48915 53431
rect 48915 53397 48924 53431
rect 48872 53388 48924 53397
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 27950 53286 28002 53338
rect 28014 53286 28066 53338
rect 28078 53286 28130 53338
rect 28142 53286 28194 53338
rect 28206 53286 28258 53338
rect 37950 53286 38002 53338
rect 38014 53286 38066 53338
rect 38078 53286 38130 53338
rect 38142 53286 38194 53338
rect 38206 53286 38258 53338
rect 47950 53286 48002 53338
rect 48014 53286 48066 53338
rect 48078 53286 48130 53338
rect 48142 53286 48194 53338
rect 48206 53286 48258 53338
rect 20720 53184 20772 53236
rect 23572 53184 23624 53236
rect 2228 53116 2280 53168
rect 5816 53048 5868 53100
rect 4804 52980 4856 53032
rect 9680 53048 9732 53100
rect 12440 53048 12492 53100
rect 16212 53116 16264 53168
rect 24860 53116 24912 53168
rect 47768 53116 47820 53168
rect 15292 53048 15344 53100
rect 19340 53048 19392 53100
rect 19892 53091 19944 53100
rect 19892 53057 19901 53091
rect 19901 53057 19935 53091
rect 19935 53057 19944 53091
rect 19892 53048 19944 53057
rect 21548 53048 21600 53100
rect 27344 53048 27396 53100
rect 7380 52980 7432 53032
rect 9956 52980 10008 53032
rect 12532 52980 12584 53032
rect 15108 52980 15160 53032
rect 17684 52980 17736 53032
rect 19616 52980 19668 53032
rect 33692 52980 33744 53032
rect 48504 53023 48556 53032
rect 48504 52989 48513 53023
rect 48513 52989 48547 53023
rect 48547 52989 48556 53023
rect 48504 52980 48556 52989
rect 12808 52912 12860 52964
rect 25320 52844 25372 52896
rect 46204 52844 46256 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 32950 52742 33002 52794
rect 33014 52742 33066 52794
rect 33078 52742 33130 52794
rect 33142 52742 33194 52794
rect 33206 52742 33258 52794
rect 42950 52742 43002 52794
rect 43014 52742 43066 52794
rect 43078 52742 43130 52794
rect 43142 52742 43194 52794
rect 43206 52742 43258 52794
rect 19892 52640 19944 52692
rect 22652 52640 22704 52692
rect 15384 52572 15436 52624
rect 1584 52504 1636 52556
rect 4160 52504 4212 52556
rect 6736 52504 6788 52556
rect 9312 52504 9364 52556
rect 11888 52504 11940 52556
rect 14464 52504 14516 52556
rect 17040 52504 17092 52556
rect 1676 52479 1728 52488
rect 1676 52445 1685 52479
rect 1685 52445 1719 52479
rect 1719 52445 1728 52479
rect 1676 52436 1728 52445
rect 4712 52436 4764 52488
rect 8300 52436 8352 52488
rect 9772 52436 9824 52488
rect 13820 52436 13872 52488
rect 16856 52436 16908 52488
rect 19432 52436 19484 52488
rect 24768 52504 24820 52556
rect 36360 52504 36412 52556
rect 48504 52479 48556 52488
rect 48504 52445 48513 52479
rect 48513 52445 48547 52479
rect 48547 52445 48556 52479
rect 48504 52436 48556 52445
rect 35532 52368 35584 52420
rect 24952 52300 25004 52352
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 27950 52198 28002 52250
rect 28014 52198 28066 52250
rect 28078 52198 28130 52250
rect 28142 52198 28194 52250
rect 28206 52198 28258 52250
rect 37950 52198 38002 52250
rect 38014 52198 38066 52250
rect 38078 52198 38130 52250
rect 38142 52198 38194 52250
rect 38206 52198 38258 52250
rect 47950 52198 48002 52250
rect 48014 52198 48066 52250
rect 48078 52198 48130 52250
rect 48142 52198 48194 52250
rect 48206 52198 48258 52250
rect 5816 52096 5868 52148
rect 10692 51960 10744 52012
rect 49240 51960 49292 52012
rect 38936 51756 38988 51808
rect 43444 51756 43496 51808
rect 49148 51799 49200 51808
rect 49148 51765 49157 51799
rect 49157 51765 49191 51799
rect 49191 51765 49200 51799
rect 49148 51756 49200 51765
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 32950 51654 33002 51706
rect 33014 51654 33066 51706
rect 33078 51654 33130 51706
rect 33142 51654 33194 51706
rect 33206 51654 33258 51706
rect 42950 51654 43002 51706
rect 43014 51654 43066 51706
rect 43078 51654 43130 51706
rect 43142 51654 43194 51706
rect 43206 51654 43258 51706
rect 4896 51552 4948 51604
rect 42156 51552 42208 51604
rect 43904 51552 43956 51604
rect 1308 51416 1360 51468
rect 49148 51416 49200 51468
rect 7564 51348 7616 51400
rect 37280 51348 37332 51400
rect 43444 51391 43496 51400
rect 43444 51357 43453 51391
rect 43453 51357 43487 51391
rect 43487 51357 43496 51391
rect 43444 51348 43496 51357
rect 48504 51391 48556 51400
rect 48504 51357 48513 51391
rect 48513 51357 48547 51391
rect 48547 51357 48556 51391
rect 48504 51348 48556 51357
rect 10968 51280 11020 51332
rect 39304 51280 39356 51332
rect 42156 51280 42208 51332
rect 23940 51212 23992 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 27950 51110 28002 51162
rect 28014 51110 28066 51162
rect 28078 51110 28130 51162
rect 28142 51110 28194 51162
rect 28206 51110 28258 51162
rect 37950 51110 38002 51162
rect 38014 51110 38066 51162
rect 38078 51110 38130 51162
rect 38142 51110 38194 51162
rect 38206 51110 38258 51162
rect 47950 51110 48002 51162
rect 48014 51110 48066 51162
rect 48078 51110 48130 51162
rect 48142 51110 48194 51162
rect 48206 51110 48258 51162
rect 8300 51008 8352 51060
rect 9680 51008 9732 51060
rect 10508 51008 10560 51060
rect 15200 51008 15252 51060
rect 19340 51008 19392 51060
rect 26240 51051 26292 51060
rect 26240 51017 26249 51051
rect 26249 51017 26283 51051
rect 26283 51017 26292 51051
rect 26240 51008 26292 51017
rect 27344 51051 27396 51060
rect 27344 51017 27353 51051
rect 27353 51017 27387 51051
rect 27387 51017 27396 51051
rect 27344 51008 27396 51017
rect 35164 50940 35216 50992
rect 5632 50872 5684 50924
rect 9956 50872 10008 50924
rect 11612 50872 11664 50924
rect 14924 50872 14976 50924
rect 19248 50872 19300 50924
rect 24492 50872 24544 50924
rect 1308 50804 1360 50856
rect 27528 50915 27580 50924
rect 27528 50881 27537 50915
rect 27537 50881 27571 50915
rect 27571 50881 27580 50915
rect 27528 50872 27580 50881
rect 31300 50872 31352 50924
rect 32312 50872 32364 50924
rect 49332 50915 49384 50924
rect 49332 50881 49341 50915
rect 49341 50881 49375 50915
rect 49375 50881 49384 50915
rect 49332 50872 49384 50881
rect 28908 50804 28960 50856
rect 29092 50804 29144 50856
rect 24860 50736 24912 50788
rect 26700 50668 26752 50720
rect 30380 50668 30432 50720
rect 30564 50668 30616 50720
rect 31024 50711 31076 50720
rect 31024 50677 31033 50711
rect 31033 50677 31067 50711
rect 31067 50677 31076 50711
rect 31024 50668 31076 50677
rect 31576 50668 31628 50720
rect 42800 50668 42852 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 32950 50566 33002 50618
rect 33014 50566 33066 50618
rect 33078 50566 33130 50618
rect 33142 50566 33194 50618
rect 33206 50566 33258 50618
rect 42950 50566 43002 50618
rect 43014 50566 43066 50618
rect 43078 50566 43130 50618
rect 43142 50566 43194 50618
rect 43206 50566 43258 50618
rect 12440 50464 12492 50516
rect 16856 50464 16908 50516
rect 19432 50464 19484 50516
rect 27528 50464 27580 50516
rect 32312 50464 32364 50516
rect 32956 50464 33008 50516
rect 8392 50439 8444 50448
rect 8392 50405 8401 50439
rect 8401 50405 8435 50439
rect 8435 50405 8444 50439
rect 8392 50396 8444 50405
rect 13728 50396 13780 50448
rect 27620 50396 27672 50448
rect 30012 50396 30064 50448
rect 13820 50328 13872 50380
rect 15108 50328 15160 50380
rect 25872 50328 25924 50380
rect 18328 50260 18380 50312
rect 30564 50260 30616 50312
rect 9588 50192 9640 50244
rect 14832 50192 14884 50244
rect 17500 50235 17552 50244
rect 17500 50201 17509 50235
rect 17509 50201 17543 50235
rect 17543 50201 17552 50235
rect 17500 50192 17552 50201
rect 25596 50192 25648 50244
rect 22468 50124 22520 50176
rect 30656 50192 30708 50244
rect 30288 50167 30340 50176
rect 30288 50133 30297 50167
rect 30297 50133 30331 50167
rect 30331 50133 30340 50167
rect 30288 50124 30340 50133
rect 35256 50396 35308 50448
rect 33508 50328 33560 50380
rect 31668 50192 31720 50244
rect 34520 50192 34572 50244
rect 31116 50124 31168 50176
rect 34428 50124 34480 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 27950 50022 28002 50074
rect 28014 50022 28066 50074
rect 28078 50022 28130 50074
rect 28142 50022 28194 50074
rect 28206 50022 28258 50074
rect 37950 50022 38002 50074
rect 38014 50022 38066 50074
rect 38078 50022 38130 50074
rect 38142 50022 38194 50074
rect 38206 50022 38258 50074
rect 47950 50022 48002 50074
rect 48014 50022 48066 50074
rect 48078 50022 48130 50074
rect 48142 50022 48194 50074
rect 48206 50022 48258 50074
rect 12808 49920 12860 49972
rect 13544 49920 13596 49972
rect 5724 49784 5776 49836
rect 16120 49920 16172 49972
rect 16212 49963 16264 49972
rect 16212 49929 16221 49963
rect 16221 49929 16255 49963
rect 16255 49929 16264 49963
rect 16212 49920 16264 49929
rect 22100 49920 22152 49972
rect 26332 49920 26384 49972
rect 15108 49895 15160 49904
rect 15108 49861 15117 49895
rect 15117 49861 15151 49895
rect 15151 49861 15160 49895
rect 15108 49852 15160 49861
rect 1308 49716 1360 49768
rect 15016 49784 15068 49836
rect 18972 49784 19024 49836
rect 21916 49784 21968 49836
rect 26608 49784 26660 49836
rect 29000 49784 29052 49836
rect 27620 49759 27672 49768
rect 27620 49725 27629 49759
rect 27629 49725 27663 49759
rect 27663 49725 27672 49759
rect 27620 49716 27672 49725
rect 31668 49920 31720 49972
rect 32588 49920 32640 49972
rect 32772 49920 32824 49972
rect 32864 49920 32916 49972
rect 34520 49920 34572 49972
rect 30472 49852 30524 49904
rect 30748 49852 30800 49904
rect 33600 49852 33652 49904
rect 35164 49963 35216 49972
rect 35164 49929 35173 49963
rect 35173 49929 35207 49963
rect 35207 49929 35216 49963
rect 35164 49920 35216 49929
rect 39028 49920 39080 49972
rect 37004 49852 37056 49904
rect 31944 49784 31996 49836
rect 32588 49784 32640 49836
rect 32680 49784 32732 49836
rect 16672 49648 16724 49700
rect 27344 49648 27396 49700
rect 30196 49716 30248 49768
rect 31576 49759 31628 49768
rect 31576 49725 31585 49759
rect 31585 49725 31619 49759
rect 31619 49725 31628 49759
rect 31576 49716 31628 49725
rect 31668 49716 31720 49768
rect 32956 49784 33008 49836
rect 34060 49716 34112 49768
rect 15200 49580 15252 49632
rect 27160 49580 27212 49632
rect 29092 49580 29144 49632
rect 29368 49623 29420 49632
rect 29368 49589 29377 49623
rect 29377 49589 29411 49623
rect 29411 49589 29420 49623
rect 29368 49580 29420 49589
rect 32496 49580 32548 49632
rect 34244 49716 34296 49768
rect 37096 49784 37148 49836
rect 49332 49827 49384 49836
rect 49332 49793 49341 49827
rect 49341 49793 49375 49827
rect 49375 49793 49384 49827
rect 49332 49784 49384 49793
rect 36636 49716 36688 49768
rect 43444 49716 43496 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 32950 49478 33002 49530
rect 33014 49478 33066 49530
rect 33078 49478 33130 49530
rect 33142 49478 33194 49530
rect 33206 49478 33258 49530
rect 42950 49478 43002 49530
rect 43014 49478 43066 49530
rect 43078 49478 43130 49530
rect 43142 49478 43194 49530
rect 43206 49478 43258 49530
rect 8484 49376 8536 49428
rect 9772 49308 9824 49360
rect 15292 49376 15344 49428
rect 24952 49376 25004 49428
rect 30104 49376 30156 49428
rect 27160 49351 27212 49360
rect 27160 49317 27169 49351
rect 27169 49317 27203 49351
rect 27203 49317 27212 49351
rect 27160 49308 27212 49317
rect 1308 49240 1360 49292
rect 29460 49308 29512 49360
rect 5816 49172 5868 49224
rect 25412 49215 25464 49224
rect 25412 49181 25421 49215
rect 25421 49181 25455 49215
rect 25455 49181 25464 49215
rect 25412 49172 25464 49181
rect 26792 49172 26844 49224
rect 26976 49172 27028 49224
rect 29368 49240 29420 49292
rect 33324 49308 33376 49360
rect 33508 49419 33560 49428
rect 33508 49385 33517 49419
rect 33517 49385 33551 49419
rect 33551 49385 33560 49419
rect 33508 49376 33560 49385
rect 34428 49376 34480 49428
rect 36544 49308 36596 49360
rect 34152 49240 34204 49292
rect 31760 49215 31812 49224
rect 31760 49181 31769 49215
rect 31769 49181 31803 49215
rect 31803 49181 31812 49215
rect 31760 49172 31812 49181
rect 33324 49172 33376 49224
rect 33600 49172 33652 49224
rect 34704 49172 34756 49224
rect 11980 49104 12032 49156
rect 16396 49104 16448 49156
rect 22744 49104 22796 49156
rect 25688 49147 25740 49156
rect 25688 49113 25697 49147
rect 25697 49113 25731 49147
rect 25731 49113 25740 49147
rect 25688 49104 25740 49113
rect 29184 49104 29236 49156
rect 30104 49147 30156 49156
rect 30104 49113 30113 49147
rect 30113 49113 30147 49147
rect 30147 49113 30156 49147
rect 30104 49104 30156 49113
rect 31024 49104 31076 49156
rect 32036 49147 32088 49156
rect 32036 49113 32045 49147
rect 32045 49113 32079 49147
rect 32079 49113 32088 49147
rect 32036 49104 32088 49113
rect 33784 49104 33836 49156
rect 37188 49104 37240 49156
rect 49056 49215 49108 49224
rect 49056 49181 49065 49215
rect 49065 49181 49099 49215
rect 49099 49181 49108 49215
rect 49056 49172 49108 49181
rect 27252 49036 27304 49088
rect 29000 49036 29052 49088
rect 30380 49036 30432 49088
rect 33416 49036 33468 49088
rect 35348 49079 35400 49088
rect 35348 49045 35357 49079
rect 35357 49045 35391 49079
rect 35391 49045 35400 49079
rect 35348 49036 35400 49045
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 27950 48934 28002 48986
rect 28014 48934 28066 48986
rect 28078 48934 28130 48986
rect 28142 48934 28194 48986
rect 28206 48934 28258 48986
rect 37950 48934 38002 48986
rect 38014 48934 38066 48986
rect 38078 48934 38130 48986
rect 38142 48934 38194 48986
rect 38206 48934 38258 48986
rect 47950 48934 48002 48986
rect 48014 48934 48066 48986
rect 48078 48934 48130 48986
rect 48142 48934 48194 48986
rect 48206 48934 48258 48986
rect 24768 48832 24820 48884
rect 27252 48764 27304 48816
rect 31852 48832 31904 48884
rect 32036 48832 32088 48884
rect 33048 48832 33100 48884
rect 33416 48832 33468 48884
rect 35256 48832 35308 48884
rect 29276 48764 29328 48816
rect 25044 48696 25096 48748
rect 23480 48628 23532 48680
rect 20996 48560 21048 48612
rect 18880 48492 18932 48544
rect 27436 48696 27488 48748
rect 26424 48671 26476 48680
rect 26424 48637 26433 48671
rect 26433 48637 26467 48671
rect 26467 48637 26476 48671
rect 26424 48628 26476 48637
rect 26516 48628 26568 48680
rect 29552 48739 29604 48748
rect 29552 48705 29561 48739
rect 29561 48705 29595 48739
rect 29595 48705 29604 48739
rect 29552 48696 29604 48705
rect 30656 48628 30708 48680
rect 31208 48628 31260 48680
rect 31852 48696 31904 48748
rect 33784 48696 33836 48748
rect 32312 48628 32364 48680
rect 28540 48560 28592 48612
rect 28908 48560 28960 48612
rect 29276 48560 29328 48612
rect 30288 48560 30340 48612
rect 27068 48492 27120 48544
rect 27160 48535 27212 48544
rect 27160 48501 27169 48535
rect 27169 48501 27203 48535
rect 27203 48501 27212 48535
rect 27160 48492 27212 48501
rect 30748 48492 30800 48544
rect 33048 48628 33100 48680
rect 34152 48671 34204 48680
rect 34152 48637 34161 48671
rect 34161 48637 34195 48671
rect 34195 48637 34204 48671
rect 34152 48628 34204 48637
rect 34336 48628 34388 48680
rect 34520 48560 34572 48612
rect 33968 48492 34020 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 32950 48390 33002 48442
rect 33014 48390 33066 48442
rect 33078 48390 33130 48442
rect 33142 48390 33194 48442
rect 33206 48390 33258 48442
rect 42950 48390 43002 48442
rect 43014 48390 43066 48442
rect 43078 48390 43130 48442
rect 43142 48390 43194 48442
rect 43206 48390 43258 48442
rect 25228 48288 25280 48340
rect 27160 48288 27212 48340
rect 27712 48288 27764 48340
rect 32312 48288 32364 48340
rect 34796 48288 34848 48340
rect 35348 48288 35400 48340
rect 28632 48220 28684 48272
rect 1308 48152 1360 48204
rect 21456 48152 21508 48204
rect 25412 48152 25464 48204
rect 26056 48152 26108 48204
rect 27712 48152 27764 48204
rect 28356 48152 28408 48204
rect 28724 48152 28776 48204
rect 30656 48152 30708 48204
rect 31024 48195 31076 48204
rect 31024 48161 31033 48195
rect 31033 48161 31067 48195
rect 31067 48161 31076 48195
rect 31024 48152 31076 48161
rect 31392 48152 31444 48204
rect 37372 48220 37424 48272
rect 35348 48152 35400 48204
rect 11060 48084 11112 48136
rect 18512 48084 18564 48136
rect 22100 48084 22152 48136
rect 24676 48084 24728 48136
rect 30012 48084 30064 48136
rect 32128 48084 32180 48136
rect 36820 48152 36872 48204
rect 22560 48059 22612 48068
rect 22560 48025 22569 48059
rect 22569 48025 22603 48059
rect 22603 48025 22612 48059
rect 22560 48016 22612 48025
rect 24584 48016 24636 48068
rect 25136 48016 25188 48068
rect 25504 48016 25556 48068
rect 27436 48016 27488 48068
rect 29092 48016 29144 48068
rect 31300 48016 31352 48068
rect 16580 47948 16632 48000
rect 19800 47948 19852 48000
rect 22008 47948 22060 48000
rect 22652 47948 22704 48000
rect 24768 47948 24820 48000
rect 27252 47948 27304 48000
rect 27712 47948 27764 48000
rect 32680 48016 32732 48068
rect 36360 48016 36412 48068
rect 36728 48059 36780 48068
rect 36728 48025 36737 48059
rect 36737 48025 36771 48059
rect 36771 48025 36780 48059
rect 36728 48016 36780 48025
rect 32772 47948 32824 48000
rect 33416 47991 33468 48000
rect 33416 47957 33425 47991
rect 33425 47957 33459 47991
rect 33459 47957 33468 47991
rect 33416 47948 33468 47957
rect 34980 47948 35032 48000
rect 35440 47948 35492 48000
rect 35716 47948 35768 48000
rect 36268 47991 36320 48000
rect 36268 47957 36277 47991
rect 36277 47957 36311 47991
rect 36311 47957 36320 47991
rect 36268 47948 36320 47957
rect 49332 48127 49384 48136
rect 49332 48093 49341 48127
rect 49341 48093 49375 48127
rect 49375 48093 49384 48127
rect 49332 48084 49384 48093
rect 39028 47948 39080 48000
rect 43352 47948 43404 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 27950 47846 28002 47898
rect 28014 47846 28066 47898
rect 28078 47846 28130 47898
rect 28142 47846 28194 47898
rect 28206 47846 28258 47898
rect 37950 47846 38002 47898
rect 38014 47846 38066 47898
rect 38078 47846 38130 47898
rect 38142 47846 38194 47898
rect 38206 47846 38258 47898
rect 47950 47846 48002 47898
rect 48014 47846 48066 47898
rect 48078 47846 48130 47898
rect 48142 47846 48194 47898
rect 48206 47846 48258 47898
rect 10692 47744 10744 47796
rect 19524 47676 19576 47728
rect 4068 47608 4120 47660
rect 15108 47608 15160 47660
rect 21088 47608 21140 47660
rect 1308 47540 1360 47592
rect 19708 47583 19760 47592
rect 19708 47549 19717 47583
rect 19717 47549 19751 47583
rect 19751 47549 19760 47583
rect 19708 47540 19760 47549
rect 21456 47787 21508 47796
rect 21456 47753 21465 47787
rect 21465 47753 21499 47787
rect 21499 47753 21508 47787
rect 21456 47744 21508 47753
rect 22008 47787 22060 47796
rect 22008 47753 22017 47787
rect 22017 47753 22051 47787
rect 22051 47753 22060 47787
rect 22008 47744 22060 47753
rect 22192 47744 22244 47796
rect 25688 47744 25740 47796
rect 22468 47719 22520 47728
rect 22468 47685 22477 47719
rect 22477 47685 22511 47719
rect 22511 47685 22520 47719
rect 22468 47676 22520 47685
rect 25136 47676 25188 47728
rect 26792 47744 26844 47796
rect 22836 47608 22888 47660
rect 24584 47608 24636 47660
rect 25504 47608 25556 47660
rect 25688 47608 25740 47660
rect 26240 47608 26292 47660
rect 27620 47719 27672 47728
rect 27620 47685 27629 47719
rect 27629 47685 27663 47719
rect 27663 47685 27672 47719
rect 27620 47676 27672 47685
rect 28264 47744 28316 47796
rect 29368 47744 29420 47796
rect 29000 47676 29052 47728
rect 28356 47608 28408 47660
rect 31760 47744 31812 47796
rect 31944 47744 31996 47796
rect 31300 47676 31352 47728
rect 32128 47676 32180 47728
rect 34796 47744 34848 47796
rect 42800 47744 42852 47796
rect 33508 47676 33560 47728
rect 33784 47676 33836 47728
rect 40132 47676 40184 47728
rect 48872 47676 48924 47728
rect 35256 47608 35308 47660
rect 37556 47608 37608 47660
rect 39764 47608 39816 47660
rect 48688 47608 48740 47660
rect 49332 47651 49384 47660
rect 49332 47617 49341 47651
rect 49341 47617 49375 47651
rect 49375 47617 49384 47651
rect 49332 47608 49384 47617
rect 22652 47583 22704 47592
rect 22652 47549 22661 47583
rect 22661 47549 22695 47583
rect 22695 47549 22704 47583
rect 22652 47540 22704 47549
rect 22100 47472 22152 47524
rect 23572 47540 23624 47592
rect 24768 47540 24820 47592
rect 27436 47540 27488 47592
rect 21272 47404 21324 47456
rect 27252 47472 27304 47524
rect 29368 47540 29420 47592
rect 31024 47540 31076 47592
rect 31760 47472 31812 47524
rect 31852 47472 31904 47524
rect 32128 47472 32180 47524
rect 32772 47472 32824 47524
rect 34888 47540 34940 47592
rect 35808 47540 35860 47592
rect 38936 47583 38988 47592
rect 38936 47549 38945 47583
rect 38945 47549 38979 47583
rect 38979 47549 38988 47583
rect 38936 47540 38988 47549
rect 25136 47404 25188 47456
rect 25504 47404 25556 47456
rect 30196 47404 30248 47456
rect 34612 47404 34664 47456
rect 34980 47404 35032 47456
rect 35716 47404 35768 47456
rect 37464 47404 37516 47456
rect 37832 47404 37884 47456
rect 42800 47404 42852 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 32950 47302 33002 47354
rect 33014 47302 33066 47354
rect 33078 47302 33130 47354
rect 33142 47302 33194 47354
rect 33206 47302 33258 47354
rect 42950 47302 43002 47354
rect 43014 47302 43066 47354
rect 43078 47302 43130 47354
rect 43142 47302 43194 47354
rect 43206 47302 43258 47354
rect 15200 47200 15252 47252
rect 22836 47200 22888 47252
rect 25688 47200 25740 47252
rect 26884 47200 26936 47252
rect 27528 47200 27580 47252
rect 28356 47243 28408 47252
rect 28356 47209 28365 47243
rect 28365 47209 28399 47243
rect 28399 47209 28408 47243
rect 28356 47200 28408 47209
rect 28632 47200 28684 47252
rect 19156 47132 19208 47184
rect 20904 47064 20956 47116
rect 22192 47132 22244 47184
rect 21456 47064 21508 47116
rect 21272 46996 21324 47048
rect 22100 46996 22152 47048
rect 25504 47132 25556 47184
rect 27620 47132 27672 47184
rect 29092 47132 29144 47184
rect 29276 47132 29328 47184
rect 29828 47132 29880 47184
rect 30932 47243 30984 47252
rect 30932 47209 30941 47243
rect 30941 47209 30975 47243
rect 30975 47209 30984 47243
rect 30932 47200 30984 47209
rect 34888 47243 34940 47252
rect 34888 47209 34897 47243
rect 34897 47209 34931 47243
rect 34931 47209 34940 47243
rect 34888 47200 34940 47209
rect 37188 47200 37240 47252
rect 24860 47064 24912 47116
rect 25872 47064 25924 47116
rect 26056 47064 26108 47116
rect 26792 47064 26844 47116
rect 29920 47064 29972 47116
rect 30196 47064 30248 47116
rect 31024 47064 31076 47116
rect 31484 47107 31536 47116
rect 31484 47073 31493 47107
rect 31493 47073 31527 47107
rect 31527 47073 31536 47107
rect 31484 47064 31536 47073
rect 32588 47107 32640 47116
rect 32588 47073 32597 47107
rect 32597 47073 32631 47107
rect 32631 47073 32640 47107
rect 32588 47064 32640 47073
rect 32680 47107 32732 47116
rect 32680 47073 32689 47107
rect 32689 47073 32723 47107
rect 32723 47073 32732 47107
rect 32680 47064 32732 47073
rect 37096 47132 37148 47184
rect 33876 47064 33928 47116
rect 34336 47064 34388 47116
rect 34428 47064 34480 47116
rect 35808 47064 35860 47116
rect 36544 47107 36596 47116
rect 36544 47073 36553 47107
rect 36553 47073 36587 47107
rect 36587 47073 36596 47107
rect 36544 47064 36596 47073
rect 36636 47107 36688 47116
rect 36636 47073 36645 47107
rect 36645 47073 36679 47107
rect 36679 47073 36688 47107
rect 36636 47064 36688 47073
rect 39028 47107 39080 47116
rect 39028 47073 39037 47107
rect 39037 47073 39071 47107
rect 39071 47073 39080 47107
rect 39028 47064 39080 47073
rect 24952 46996 25004 47048
rect 25320 47039 25372 47048
rect 25320 47005 25329 47039
rect 25329 47005 25363 47039
rect 25363 47005 25372 47039
rect 25320 46996 25372 47005
rect 28816 46996 28868 47048
rect 30472 46996 30524 47048
rect 33692 47039 33744 47048
rect 33692 47005 33701 47039
rect 33701 47005 33735 47039
rect 33735 47005 33744 47039
rect 33692 46996 33744 47005
rect 34704 46996 34756 47048
rect 35256 47039 35308 47048
rect 35256 47005 35265 47039
rect 35265 47005 35299 47039
rect 35299 47005 35308 47039
rect 35256 46996 35308 47005
rect 38292 46996 38344 47048
rect 43444 46996 43496 47048
rect 20720 46928 20772 46980
rect 22008 46928 22060 46980
rect 23848 46928 23900 46980
rect 24584 46928 24636 46980
rect 25780 46928 25832 46980
rect 26148 46928 26200 46980
rect 21180 46860 21232 46912
rect 23480 46860 23532 46912
rect 26884 46928 26936 46980
rect 28356 46928 28408 46980
rect 28540 46928 28592 46980
rect 30288 46928 30340 46980
rect 30564 46928 30616 46980
rect 28632 46860 28684 46912
rect 29092 46860 29144 46912
rect 31576 46860 31628 46912
rect 36084 46928 36136 46980
rect 36452 46971 36504 46980
rect 36452 46937 36461 46971
rect 36461 46937 36495 46971
rect 36495 46937 36504 46971
rect 36452 46928 36504 46937
rect 40132 46928 40184 46980
rect 33324 46903 33376 46912
rect 33324 46869 33333 46903
rect 33333 46869 33367 46903
rect 33367 46869 33376 46903
rect 33324 46860 33376 46869
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 27950 46758 28002 46810
rect 28014 46758 28066 46810
rect 28078 46758 28130 46810
rect 28142 46758 28194 46810
rect 28206 46758 28258 46810
rect 37950 46758 38002 46810
rect 38014 46758 38066 46810
rect 38078 46758 38130 46810
rect 38142 46758 38194 46810
rect 38206 46758 38258 46810
rect 47950 46758 48002 46810
rect 48014 46758 48066 46810
rect 48078 46758 48130 46810
rect 48142 46758 48194 46810
rect 48206 46758 48258 46810
rect 10968 46656 11020 46708
rect 22560 46656 22612 46708
rect 24768 46656 24820 46708
rect 21640 46588 21692 46640
rect 23848 46588 23900 46640
rect 24676 46588 24728 46640
rect 26056 46656 26108 46708
rect 26792 46656 26844 46708
rect 28908 46656 28960 46708
rect 29184 46699 29236 46708
rect 29184 46665 29193 46699
rect 29193 46665 29227 46699
rect 29227 46665 29236 46699
rect 29184 46656 29236 46665
rect 29460 46656 29512 46708
rect 25688 46588 25740 46640
rect 27896 46631 27948 46640
rect 27896 46597 27905 46631
rect 27905 46597 27939 46631
rect 27939 46597 27948 46631
rect 27896 46588 27948 46597
rect 28540 46588 28592 46640
rect 28632 46588 28684 46640
rect 32588 46656 32640 46708
rect 31300 46588 31352 46640
rect 31668 46588 31720 46640
rect 33692 46656 33744 46708
rect 36544 46588 36596 46640
rect 39304 46588 39356 46640
rect 8668 46520 8720 46572
rect 13728 46520 13780 46572
rect 21088 46520 21140 46572
rect 24860 46563 24912 46572
rect 24860 46529 24869 46563
rect 24869 46529 24903 46563
rect 24903 46529 24912 46563
rect 24860 46520 24912 46529
rect 1308 46452 1360 46504
rect 19708 46495 19760 46504
rect 19708 46461 19717 46495
rect 19717 46461 19751 46495
rect 19751 46461 19760 46495
rect 19708 46452 19760 46461
rect 21180 46452 21232 46504
rect 22836 46452 22888 46504
rect 25872 46452 25924 46504
rect 26148 46452 26200 46504
rect 27528 46427 27580 46436
rect 27528 46393 27537 46427
rect 27537 46393 27571 46427
rect 27571 46393 27580 46427
rect 27528 46384 27580 46393
rect 21640 46316 21692 46368
rect 22100 46316 22152 46368
rect 22652 46316 22704 46368
rect 25228 46316 25280 46368
rect 25320 46316 25372 46368
rect 29092 46452 29144 46504
rect 30012 46563 30064 46572
rect 30012 46529 30021 46563
rect 30021 46529 30055 46563
rect 30055 46529 30064 46563
rect 30012 46520 30064 46529
rect 31852 46520 31904 46572
rect 32496 46520 32548 46572
rect 28908 46316 28960 46368
rect 30840 46452 30892 46504
rect 31760 46495 31812 46504
rect 31760 46461 31769 46495
rect 31769 46461 31803 46495
rect 31803 46461 31812 46495
rect 31760 46452 31812 46461
rect 32772 46495 32824 46504
rect 32772 46461 32781 46495
rect 32781 46461 32815 46495
rect 32815 46461 32824 46495
rect 32772 46452 32824 46461
rect 34520 46563 34572 46572
rect 34520 46529 34529 46563
rect 34529 46529 34563 46563
rect 34563 46529 34572 46563
rect 34520 46520 34572 46529
rect 49056 46563 49108 46572
rect 49056 46529 49065 46563
rect 49065 46529 49099 46563
rect 49099 46529 49108 46563
rect 49056 46520 49108 46529
rect 34796 46495 34848 46504
rect 34796 46461 34805 46495
rect 34805 46461 34839 46495
rect 34839 46461 34848 46495
rect 34796 46452 34848 46461
rect 35348 46452 35400 46504
rect 30288 46316 30340 46368
rect 30472 46316 30524 46368
rect 32312 46359 32364 46368
rect 32312 46325 32321 46359
rect 32321 46325 32355 46359
rect 32355 46325 32364 46359
rect 32312 46316 32364 46325
rect 32588 46316 32640 46368
rect 34428 46316 34480 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 32950 46214 33002 46266
rect 33014 46214 33066 46266
rect 33078 46214 33130 46266
rect 33142 46214 33194 46266
rect 33206 46214 33258 46266
rect 42950 46214 43002 46266
rect 43014 46214 43066 46266
rect 43078 46214 43130 46266
rect 43142 46214 43194 46266
rect 43206 46214 43258 46266
rect 11060 46155 11112 46164
rect 11060 46121 11069 46155
rect 11069 46121 11103 46155
rect 11103 46121 11112 46155
rect 11060 46112 11112 46121
rect 19248 46112 19300 46164
rect 21732 46112 21784 46164
rect 1308 45976 1360 46028
rect 20996 46019 21048 46028
rect 20996 45985 21005 46019
rect 21005 45985 21039 46019
rect 21039 45985 21048 46019
rect 20996 45976 21048 45985
rect 21364 45976 21416 46028
rect 12256 45908 12308 45960
rect 19616 45951 19668 45960
rect 19616 45917 19625 45951
rect 19625 45917 19659 45951
rect 19659 45917 19668 45951
rect 19616 45908 19668 45917
rect 19708 45908 19760 45960
rect 22100 45976 22152 46028
rect 23296 45976 23348 46028
rect 23480 46155 23532 46164
rect 23480 46121 23489 46155
rect 23489 46121 23523 46155
rect 23523 46121 23532 46155
rect 23480 46112 23532 46121
rect 25044 46155 25096 46164
rect 25044 46121 25053 46155
rect 25053 46121 25087 46155
rect 25087 46121 25096 46155
rect 25044 46112 25096 46121
rect 25412 46112 25464 46164
rect 29920 46112 29972 46164
rect 30656 46112 30708 46164
rect 24308 46044 24360 46096
rect 26976 46044 27028 46096
rect 29000 46044 29052 46096
rect 32772 46112 32824 46164
rect 35440 46112 35492 46164
rect 31024 46087 31076 46096
rect 31024 46053 31033 46087
rect 31033 46053 31067 46087
rect 31067 46053 31076 46087
rect 31024 46044 31076 46053
rect 26700 46019 26752 46028
rect 26700 45985 26709 46019
rect 26709 45985 26743 46019
rect 26743 45985 26752 46019
rect 26700 45976 26752 45985
rect 26792 46019 26844 46028
rect 26792 45985 26801 46019
rect 26801 45985 26835 46019
rect 26835 45985 26844 46019
rect 26792 45976 26844 45985
rect 29460 45976 29512 46028
rect 30012 45976 30064 46028
rect 30196 45976 30248 46028
rect 30840 45976 30892 46028
rect 31576 46019 31628 46028
rect 31576 45985 31585 46019
rect 31585 45985 31619 46019
rect 31619 45985 31628 46019
rect 31576 45976 31628 45985
rect 34520 45976 34572 46028
rect 34888 45976 34940 46028
rect 35440 45976 35492 46028
rect 36820 45976 36872 46028
rect 25504 45908 25556 45960
rect 25964 45908 26016 45960
rect 27344 45908 27396 45960
rect 29184 45908 29236 45960
rect 29920 45908 29972 45960
rect 31668 45908 31720 45960
rect 32496 45908 32548 45960
rect 12532 45840 12584 45892
rect 13636 45840 13688 45892
rect 18604 45772 18656 45824
rect 23848 45840 23900 45892
rect 27712 45883 27764 45892
rect 27712 45849 27721 45883
rect 27721 45849 27755 45883
rect 27755 45849 27764 45883
rect 27712 45840 27764 45849
rect 31300 45840 31352 45892
rect 23388 45772 23440 45824
rect 23480 45772 23532 45824
rect 26700 45772 26752 45824
rect 26792 45772 26844 45824
rect 29276 45772 29328 45824
rect 32956 45840 33008 45892
rect 33232 45883 33284 45892
rect 33232 45849 33241 45883
rect 33241 45849 33275 45883
rect 33275 45849 33284 45883
rect 33232 45840 33284 45849
rect 34152 45951 34204 45960
rect 34152 45917 34161 45951
rect 34161 45917 34195 45951
rect 34195 45917 34204 45951
rect 34152 45908 34204 45917
rect 36544 45908 36596 45960
rect 37832 45951 37884 45960
rect 37832 45917 37841 45951
rect 37841 45917 37875 45951
rect 37875 45917 37884 45951
rect 37832 45908 37884 45917
rect 34244 45840 34296 45892
rect 35348 45840 35400 45892
rect 35532 45772 35584 45824
rect 37188 45772 37240 45824
rect 37740 45772 37792 45824
rect 49056 45951 49108 45960
rect 49056 45917 49065 45951
rect 49065 45917 49099 45951
rect 49099 45917 49108 45951
rect 49056 45908 49108 45917
rect 39120 45772 39172 45824
rect 48596 45772 48648 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 27950 45670 28002 45722
rect 28014 45670 28066 45722
rect 28078 45670 28130 45722
rect 28142 45670 28194 45722
rect 28206 45670 28258 45722
rect 37950 45670 38002 45722
rect 38014 45670 38066 45722
rect 38078 45670 38130 45722
rect 38142 45670 38194 45722
rect 38206 45670 38258 45722
rect 47950 45670 48002 45722
rect 48014 45670 48066 45722
rect 48078 45670 48130 45722
rect 48142 45670 48194 45722
rect 48206 45670 48258 45722
rect 7564 45500 7616 45552
rect 20812 45568 20864 45620
rect 12808 45432 12860 45484
rect 16580 45432 16632 45484
rect 23756 45500 23808 45552
rect 23940 45543 23992 45552
rect 23940 45509 23949 45543
rect 23949 45509 23983 45543
rect 23983 45509 23992 45543
rect 23940 45500 23992 45509
rect 25412 45568 25464 45620
rect 19708 45475 19760 45484
rect 19708 45441 19717 45475
rect 19717 45441 19751 45475
rect 19751 45441 19760 45475
rect 19708 45432 19760 45441
rect 21088 45432 21140 45484
rect 23848 45475 23900 45484
rect 23848 45441 23857 45475
rect 23857 45441 23891 45475
rect 23891 45441 23900 45475
rect 23848 45432 23900 45441
rect 25044 45475 25096 45484
rect 25044 45441 25053 45475
rect 25053 45441 25087 45475
rect 25087 45441 25096 45475
rect 25044 45432 25096 45441
rect 13820 45364 13872 45416
rect 19984 45407 20036 45416
rect 19984 45373 19993 45407
rect 19993 45373 20027 45407
rect 20027 45373 20036 45407
rect 19984 45364 20036 45373
rect 20720 45364 20772 45416
rect 9956 45296 10008 45348
rect 18328 45296 18380 45348
rect 20996 45296 21048 45348
rect 21548 45296 21600 45348
rect 22836 45407 22888 45416
rect 22836 45373 22845 45407
rect 22845 45373 22879 45407
rect 22879 45373 22888 45407
rect 22836 45364 22888 45373
rect 24032 45407 24084 45416
rect 24032 45373 24041 45407
rect 24041 45373 24075 45407
rect 24075 45373 24084 45407
rect 24032 45364 24084 45373
rect 24124 45364 24176 45416
rect 26424 45568 26476 45620
rect 26700 45568 26752 45620
rect 28172 45568 28224 45620
rect 28264 45568 28316 45620
rect 28632 45568 28684 45620
rect 32312 45568 32364 45620
rect 33416 45568 33468 45620
rect 34152 45611 34204 45620
rect 34152 45577 34161 45611
rect 34161 45577 34195 45611
rect 34195 45577 34204 45611
rect 34152 45568 34204 45577
rect 34244 45568 34296 45620
rect 38660 45568 38712 45620
rect 26332 45543 26384 45552
rect 26332 45509 26341 45543
rect 26341 45509 26375 45543
rect 26375 45509 26384 45543
rect 26332 45500 26384 45509
rect 27712 45500 27764 45552
rect 28448 45500 28500 45552
rect 29644 45500 29696 45552
rect 32496 45500 32548 45552
rect 32864 45500 32916 45552
rect 33232 45500 33284 45552
rect 34336 45500 34388 45552
rect 28632 45432 28684 45484
rect 29000 45432 29052 45484
rect 29736 45432 29788 45484
rect 30564 45432 30616 45484
rect 34060 45432 34112 45484
rect 39764 45500 39816 45552
rect 26608 45364 26660 45416
rect 26976 45364 27028 45416
rect 28724 45296 28776 45348
rect 29276 45364 29328 45416
rect 30288 45407 30340 45416
rect 30288 45373 30297 45407
rect 30297 45373 30331 45407
rect 30331 45373 30340 45407
rect 30288 45364 30340 45373
rect 30380 45364 30432 45416
rect 32036 45364 32088 45416
rect 32772 45364 32824 45416
rect 33508 45364 33560 45416
rect 34796 45364 34848 45416
rect 36452 45364 36504 45416
rect 30104 45296 30156 45348
rect 31116 45296 31168 45348
rect 31300 45296 31352 45348
rect 33232 45296 33284 45348
rect 34152 45296 34204 45348
rect 37464 45364 37516 45416
rect 38016 45407 38068 45416
rect 38016 45373 38025 45407
rect 38025 45373 38059 45407
rect 38059 45373 38068 45407
rect 38016 45364 38068 45373
rect 42800 45432 42852 45484
rect 39488 45364 39540 45416
rect 6828 45228 6880 45280
rect 20444 45228 20496 45280
rect 22192 45228 22244 45280
rect 23388 45228 23440 45280
rect 24768 45228 24820 45280
rect 28172 45228 28224 45280
rect 29276 45228 29328 45280
rect 29736 45271 29788 45280
rect 29736 45237 29745 45271
rect 29745 45237 29779 45271
rect 29779 45237 29788 45271
rect 29736 45228 29788 45237
rect 35256 45228 35308 45280
rect 36176 45271 36228 45280
rect 36176 45237 36185 45271
rect 36185 45237 36219 45271
rect 36219 45237 36228 45271
rect 36176 45228 36228 45237
rect 37372 45228 37424 45280
rect 46204 45228 46256 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 32950 45126 33002 45178
rect 33014 45126 33066 45178
rect 33078 45126 33130 45178
rect 33142 45126 33194 45178
rect 33206 45126 33258 45178
rect 42950 45126 43002 45178
rect 43014 45126 43066 45178
rect 43078 45126 43130 45178
rect 43142 45126 43194 45178
rect 43206 45126 43258 45178
rect 5632 45024 5684 45076
rect 11612 45024 11664 45076
rect 19800 45024 19852 45076
rect 18696 44956 18748 45008
rect 21824 45024 21876 45076
rect 1308 44888 1360 44940
rect 19524 44888 19576 44940
rect 20168 44888 20220 44940
rect 27068 45024 27120 45076
rect 31208 45024 31260 45076
rect 34152 45024 34204 45076
rect 34796 45024 34848 45076
rect 38016 45024 38068 45076
rect 25872 44956 25924 45008
rect 11060 44820 11112 44872
rect 15016 44820 15068 44872
rect 18512 44863 18564 44872
rect 18512 44829 18521 44863
rect 18521 44829 18555 44863
rect 18555 44829 18564 44863
rect 18512 44820 18564 44829
rect 19708 44820 19760 44872
rect 21456 44820 21508 44872
rect 23940 44931 23992 44940
rect 23940 44897 23949 44931
rect 23949 44897 23983 44931
rect 23983 44897 23992 44931
rect 23940 44888 23992 44897
rect 25596 44888 25648 44940
rect 28724 44956 28776 45008
rect 29276 44956 29328 45008
rect 33600 44956 33652 45008
rect 27252 44931 27304 44940
rect 27252 44897 27261 44931
rect 27261 44897 27295 44931
rect 27295 44897 27304 44931
rect 27252 44888 27304 44897
rect 27344 44931 27396 44940
rect 27344 44897 27353 44931
rect 27353 44897 27387 44931
rect 27387 44897 27396 44931
rect 27344 44888 27396 44897
rect 24032 44820 24084 44872
rect 13544 44752 13596 44804
rect 16304 44752 16356 44804
rect 20168 44795 20220 44804
rect 20168 44761 20177 44795
rect 20177 44761 20211 44795
rect 20211 44761 20220 44795
rect 20168 44752 20220 44761
rect 21180 44752 21232 44804
rect 21824 44752 21876 44804
rect 27528 44820 27580 44872
rect 28448 44820 28500 44872
rect 28724 44820 28776 44872
rect 31576 44888 31628 44940
rect 31760 44888 31812 44940
rect 32680 44888 32732 44940
rect 33140 44888 33192 44940
rect 33416 44931 33468 44940
rect 33416 44897 33425 44931
rect 33425 44897 33459 44931
rect 33459 44897 33468 44931
rect 33416 44888 33468 44897
rect 34060 44888 34112 44940
rect 34888 44931 34940 44940
rect 34888 44897 34897 44931
rect 34897 44897 34931 44931
rect 34931 44897 34940 44931
rect 34888 44888 34940 44897
rect 37372 44956 37424 45008
rect 47400 44956 47452 45008
rect 35900 44888 35952 44940
rect 36912 44888 36964 44940
rect 37740 44888 37792 44940
rect 38660 44888 38712 44940
rect 19064 44684 19116 44736
rect 19892 44684 19944 44736
rect 21732 44684 21784 44736
rect 24768 44752 24820 44804
rect 23664 44727 23716 44736
rect 23664 44693 23673 44727
rect 23673 44693 23707 44727
rect 23707 44693 23716 44727
rect 23664 44684 23716 44693
rect 24400 44684 24452 44736
rect 25044 44684 25096 44736
rect 25596 44752 25648 44804
rect 29092 44752 29144 44804
rect 33968 44820 34020 44872
rect 37096 44863 37148 44872
rect 37096 44829 37105 44863
rect 37105 44829 37139 44863
rect 37139 44829 37148 44863
rect 37096 44820 37148 44829
rect 33324 44752 33376 44804
rect 35164 44795 35216 44804
rect 35164 44761 35173 44795
rect 35173 44761 35207 44795
rect 35207 44761 35216 44795
rect 35164 44752 35216 44761
rect 36544 44752 36596 44804
rect 37004 44752 37056 44804
rect 26608 44684 26660 44736
rect 30840 44684 30892 44736
rect 31208 44684 31260 44736
rect 32496 44684 32548 44736
rect 35808 44684 35860 44736
rect 43352 44820 43404 44872
rect 49056 44863 49108 44872
rect 49056 44829 49065 44863
rect 49065 44829 49099 44863
rect 49099 44829 49108 44863
rect 49056 44820 49108 44829
rect 39672 44752 39724 44804
rect 37556 44727 37608 44736
rect 37556 44693 37565 44727
rect 37565 44693 37599 44727
rect 37599 44693 37608 44727
rect 37556 44684 37608 44693
rect 38384 44727 38436 44736
rect 38384 44693 38393 44727
rect 38393 44693 38427 44727
rect 38427 44693 38436 44727
rect 38384 44684 38436 44693
rect 38752 44727 38804 44736
rect 38752 44693 38761 44727
rect 38761 44693 38795 44727
rect 38795 44693 38804 44727
rect 38752 44684 38804 44693
rect 48596 44684 48648 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 27950 44582 28002 44634
rect 28014 44582 28066 44634
rect 28078 44582 28130 44634
rect 28142 44582 28194 44634
rect 28206 44582 28258 44634
rect 37950 44582 38002 44634
rect 38014 44582 38066 44634
rect 38078 44582 38130 44634
rect 38142 44582 38194 44634
rect 38206 44582 38258 44634
rect 47950 44582 48002 44634
rect 48014 44582 48066 44634
rect 48078 44582 48130 44634
rect 48142 44582 48194 44634
rect 48206 44582 48258 44634
rect 2044 44480 2096 44532
rect 9588 44480 9640 44532
rect 14924 44480 14976 44532
rect 17500 44480 17552 44532
rect 5540 44455 5592 44464
rect 5540 44421 5549 44455
rect 5549 44421 5583 44455
rect 5583 44421 5592 44455
rect 5540 44412 5592 44421
rect 6828 44455 6880 44464
rect 6828 44421 6837 44455
rect 6837 44421 6871 44455
rect 6871 44421 6880 44455
rect 6828 44412 6880 44421
rect 3424 44344 3476 44396
rect 5356 44387 5408 44396
rect 5356 44353 5365 44387
rect 5365 44353 5399 44387
rect 5399 44353 5408 44387
rect 5356 44344 5408 44353
rect 12440 44344 12492 44396
rect 2044 44319 2096 44328
rect 2044 44285 2053 44319
rect 2053 44285 2087 44319
rect 2087 44285 2096 44319
rect 2044 44276 2096 44285
rect 16304 44387 16356 44396
rect 16304 44353 16313 44387
rect 16313 44353 16347 44387
rect 16347 44353 16356 44387
rect 16304 44344 16356 44353
rect 20076 44480 20128 44532
rect 21456 44480 21508 44532
rect 22008 44523 22060 44532
rect 22008 44489 22017 44523
rect 22017 44489 22051 44523
rect 22051 44489 22060 44523
rect 22008 44480 22060 44489
rect 24492 44480 24544 44532
rect 27620 44480 27672 44532
rect 28724 44523 28776 44532
rect 28724 44489 28733 44523
rect 28733 44489 28767 44523
rect 28767 44489 28776 44523
rect 28724 44480 28776 44489
rect 30380 44480 30432 44532
rect 30748 44480 30800 44532
rect 37556 44480 37608 44532
rect 37648 44480 37700 44532
rect 38292 44480 38344 44532
rect 39672 44523 39724 44532
rect 39672 44489 39681 44523
rect 39681 44489 39715 44523
rect 39715 44489 39724 44523
rect 39672 44480 39724 44489
rect 20444 44412 20496 44464
rect 21088 44344 21140 44396
rect 22284 44344 22336 44396
rect 11888 44208 11940 44260
rect 14832 44208 14884 44260
rect 6920 44183 6972 44192
rect 6920 44149 6929 44183
rect 6929 44149 6963 44183
rect 6963 44149 6972 44183
rect 6920 44140 6972 44149
rect 17960 44208 18012 44260
rect 18328 44140 18380 44192
rect 19340 44276 19392 44328
rect 21272 44319 21324 44328
rect 21272 44285 21281 44319
rect 21281 44285 21315 44319
rect 21315 44285 21324 44319
rect 21272 44276 21324 44285
rect 22376 44276 22428 44328
rect 23572 44412 23624 44464
rect 27436 44412 27488 44464
rect 27804 44412 27856 44464
rect 28540 44412 28592 44464
rect 25596 44344 25648 44396
rect 26332 44344 26384 44396
rect 23296 44319 23348 44328
rect 23296 44285 23305 44319
rect 23305 44285 23339 44319
rect 23339 44285 23348 44319
rect 23296 44276 23348 44285
rect 20076 44208 20128 44260
rect 19708 44140 19760 44192
rect 20168 44183 20220 44192
rect 20168 44149 20177 44183
rect 20177 44149 20211 44183
rect 20211 44149 20220 44183
rect 20168 44140 20220 44149
rect 20260 44140 20312 44192
rect 21548 44208 21600 44260
rect 23940 44276 23992 44328
rect 24952 44276 25004 44328
rect 26148 44276 26200 44328
rect 27528 44276 27580 44328
rect 25872 44208 25924 44260
rect 28540 44276 28592 44328
rect 30104 44387 30156 44396
rect 30104 44353 30113 44387
rect 30113 44353 30147 44387
rect 30147 44353 30156 44387
rect 30104 44344 30156 44353
rect 30012 44276 30064 44328
rect 30472 44412 30524 44464
rect 32128 44344 32180 44396
rect 32220 44344 32272 44396
rect 32680 44344 32732 44396
rect 29000 44208 29052 44260
rect 29184 44208 29236 44260
rect 32404 44276 32456 44328
rect 32588 44276 32640 44328
rect 33324 44276 33376 44328
rect 33508 44276 33560 44328
rect 30840 44208 30892 44260
rect 23388 44140 23440 44192
rect 26516 44140 26568 44192
rect 28724 44140 28776 44192
rect 30288 44140 30340 44192
rect 33600 44140 33652 44192
rect 33692 44140 33744 44192
rect 35348 44387 35400 44396
rect 35348 44353 35357 44387
rect 35357 44353 35391 44387
rect 35391 44353 35400 44387
rect 35348 44344 35400 44353
rect 38384 44412 38436 44464
rect 37740 44344 37792 44396
rect 49332 44387 49384 44396
rect 49332 44353 49341 44387
rect 49341 44353 49375 44387
rect 49375 44353 49384 44387
rect 49332 44344 49384 44353
rect 34336 44319 34388 44328
rect 34336 44285 34345 44319
rect 34345 44285 34379 44319
rect 34379 44285 34388 44319
rect 34336 44276 34388 44285
rect 34428 44276 34480 44328
rect 35716 44276 35768 44328
rect 36176 44208 36228 44260
rect 34612 44140 34664 44192
rect 35624 44140 35676 44192
rect 35808 44183 35860 44192
rect 35808 44149 35817 44183
rect 35817 44149 35851 44183
rect 35851 44149 35860 44183
rect 35808 44140 35860 44149
rect 36820 44276 36872 44328
rect 37188 44276 37240 44328
rect 38016 44319 38068 44328
rect 38016 44285 38025 44319
rect 38025 44285 38059 44319
rect 38059 44285 38068 44319
rect 38016 44276 38068 44285
rect 39488 44276 39540 44328
rect 40132 44319 40184 44328
rect 40132 44285 40141 44319
rect 40141 44285 40175 44319
rect 40175 44285 40184 44319
rect 40132 44276 40184 44285
rect 37464 44251 37516 44260
rect 37464 44217 37473 44251
rect 37473 44217 37507 44251
rect 37507 44217 37516 44251
rect 37464 44208 37516 44217
rect 37556 44208 37608 44260
rect 38660 44140 38712 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 32950 44038 33002 44090
rect 33014 44038 33066 44090
rect 33078 44038 33130 44090
rect 33142 44038 33194 44090
rect 33206 44038 33258 44090
rect 42950 44038 43002 44090
rect 43014 44038 43066 44090
rect 43078 44038 43130 44090
rect 43142 44038 43194 44090
rect 43206 44038 43258 44090
rect 5816 43936 5868 43988
rect 11060 43936 11112 43988
rect 16120 43979 16172 43988
rect 16120 43945 16129 43979
rect 16129 43945 16163 43979
rect 16163 43945 16172 43979
rect 16120 43936 16172 43945
rect 4712 43911 4764 43920
rect 4712 43877 4721 43911
rect 4721 43877 4755 43911
rect 4755 43877 4764 43911
rect 4712 43868 4764 43877
rect 5724 43911 5776 43920
rect 5724 43877 5733 43911
rect 5733 43877 5767 43911
rect 5767 43877 5776 43911
rect 5724 43868 5776 43877
rect 12256 43911 12308 43920
rect 12256 43877 12265 43911
rect 12265 43877 12299 43911
rect 12299 43877 12308 43911
rect 12256 43868 12308 43877
rect 19984 43936 20036 43988
rect 20076 43936 20128 43988
rect 24124 43936 24176 43988
rect 26608 43979 26660 43988
rect 26608 43945 26617 43979
rect 26617 43945 26651 43979
rect 26651 43945 26660 43979
rect 26608 43936 26660 43945
rect 29552 43936 29604 43988
rect 31300 43936 31352 43988
rect 49240 43936 49292 43988
rect 9588 43732 9640 43784
rect 19248 43868 19300 43920
rect 32680 43868 32732 43920
rect 33968 43868 34020 43920
rect 38660 43868 38712 43920
rect 16856 43800 16908 43852
rect 17868 43800 17920 43852
rect 18420 43800 18472 43852
rect 18696 43800 18748 43852
rect 19340 43800 19392 43852
rect 21364 43800 21416 43852
rect 22468 43800 22520 43852
rect 23388 43843 23440 43852
rect 23388 43809 23397 43843
rect 23397 43809 23431 43843
rect 23431 43809 23440 43843
rect 23388 43800 23440 43809
rect 27436 43800 27488 43852
rect 29368 43800 29420 43852
rect 30012 43800 30064 43852
rect 31944 43800 31996 43852
rect 32220 43800 32272 43852
rect 32588 43800 32640 43852
rect 15936 43732 15988 43784
rect 16488 43732 16540 43784
rect 22652 43732 22704 43784
rect 24584 43732 24636 43784
rect 30932 43732 30984 43784
rect 33048 43800 33100 43852
rect 33692 43800 33744 43852
rect 33784 43800 33836 43852
rect 34888 43800 34940 43852
rect 35716 43800 35768 43852
rect 36544 43800 36596 43852
rect 4804 43664 4856 43716
rect 13636 43664 13688 43716
rect 14556 43596 14608 43648
rect 18420 43664 18472 43716
rect 19340 43664 19392 43716
rect 18328 43596 18380 43648
rect 19524 43639 19576 43648
rect 19524 43605 19533 43639
rect 19533 43605 19567 43639
rect 19567 43605 19576 43639
rect 19524 43596 19576 43605
rect 19892 43639 19944 43648
rect 19892 43605 19901 43639
rect 19901 43605 19935 43639
rect 19935 43605 19944 43639
rect 19892 43596 19944 43605
rect 20720 43596 20772 43648
rect 21272 43596 21324 43648
rect 24492 43664 24544 43716
rect 24676 43664 24728 43716
rect 24860 43596 24912 43648
rect 25044 43664 25096 43716
rect 25228 43664 25280 43716
rect 25596 43664 25648 43716
rect 27712 43664 27764 43716
rect 31024 43664 31076 43716
rect 31576 43707 31628 43716
rect 31576 43673 31585 43707
rect 31585 43673 31619 43707
rect 31619 43673 31628 43707
rect 31576 43664 31628 43673
rect 32864 43664 32916 43716
rect 33232 43664 33284 43716
rect 37280 43843 37332 43852
rect 37280 43809 37289 43843
rect 37289 43809 37323 43843
rect 37323 43809 37332 43843
rect 37280 43800 37332 43809
rect 30748 43596 30800 43648
rect 32588 43596 32640 43648
rect 33508 43596 33560 43648
rect 33968 43639 34020 43648
rect 33968 43605 33977 43639
rect 33977 43605 34011 43639
rect 34011 43605 34020 43639
rect 33968 43596 34020 43605
rect 36360 43596 36412 43648
rect 36820 43639 36872 43648
rect 36820 43605 36829 43639
rect 36829 43605 36863 43639
rect 36863 43605 36872 43639
rect 36820 43596 36872 43605
rect 37556 43707 37608 43716
rect 37556 43673 37565 43707
rect 37565 43673 37599 43707
rect 37599 43673 37608 43707
rect 37556 43664 37608 43673
rect 38844 43596 38896 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 27950 43494 28002 43546
rect 28014 43494 28066 43546
rect 28078 43494 28130 43546
rect 28142 43494 28194 43546
rect 28206 43494 28258 43546
rect 37950 43494 38002 43546
rect 38014 43494 38066 43546
rect 38078 43494 38130 43546
rect 38142 43494 38194 43546
rect 38206 43494 38258 43546
rect 47950 43494 48002 43546
rect 48014 43494 48066 43546
rect 48078 43494 48130 43546
rect 48142 43494 48194 43546
rect 48206 43494 48258 43546
rect 4068 43392 4120 43444
rect 8668 43435 8720 43444
rect 8668 43401 8677 43435
rect 8677 43401 8711 43435
rect 8711 43401 8720 43435
rect 8668 43392 8720 43401
rect 15108 43392 15160 43444
rect 15936 43435 15988 43444
rect 15936 43401 15945 43435
rect 15945 43401 15979 43435
rect 15979 43401 15988 43435
rect 15936 43392 15988 43401
rect 20260 43392 20312 43444
rect 21364 43392 21416 43444
rect 26424 43435 26476 43444
rect 6920 43324 6972 43376
rect 20076 43324 20128 43376
rect 1308 43188 1360 43240
rect 9496 43188 9548 43240
rect 17776 43256 17828 43308
rect 18880 43256 18932 43308
rect 19708 43299 19760 43308
rect 19708 43265 19717 43299
rect 19717 43265 19751 43299
rect 19751 43265 19760 43299
rect 19708 43256 19760 43265
rect 21088 43256 21140 43308
rect 18328 43188 18380 43240
rect 17040 43120 17092 43172
rect 18512 43095 18564 43104
rect 18512 43061 18521 43095
rect 18521 43061 18555 43095
rect 18555 43061 18564 43095
rect 18512 43052 18564 43061
rect 20628 43188 20680 43240
rect 22468 43324 22520 43376
rect 26424 43401 26433 43435
rect 26433 43401 26467 43435
rect 26467 43401 26476 43435
rect 26424 43392 26476 43401
rect 26700 43392 26752 43444
rect 27528 43392 27580 43444
rect 28264 43392 28316 43444
rect 31576 43392 31628 43444
rect 33232 43392 33284 43444
rect 22836 43324 22888 43376
rect 24952 43367 25004 43376
rect 24952 43333 24961 43367
rect 24961 43333 24995 43367
rect 24995 43333 25004 43367
rect 24952 43324 25004 43333
rect 25596 43324 25648 43376
rect 32864 43324 32916 43376
rect 35532 43392 35584 43444
rect 36268 43392 36320 43444
rect 49240 43435 49292 43444
rect 49240 43401 49249 43435
rect 49249 43401 49283 43435
rect 49283 43401 49292 43435
rect 49240 43392 49292 43401
rect 35164 43324 35216 43376
rect 27252 43256 27304 43308
rect 29460 43299 29512 43308
rect 29460 43265 29469 43299
rect 29469 43265 29503 43299
rect 29503 43265 29512 43299
rect 29460 43256 29512 43265
rect 31944 43256 31996 43308
rect 35348 43256 35400 43308
rect 49148 43299 49200 43308
rect 49148 43265 49157 43299
rect 49157 43265 49191 43299
rect 49191 43265 49200 43299
rect 49148 43256 49200 43265
rect 21640 43052 21692 43104
rect 22468 43231 22520 43240
rect 22468 43197 22477 43231
rect 22477 43197 22511 43231
rect 22511 43197 22520 43231
rect 22468 43188 22520 43197
rect 23296 43188 23348 43240
rect 29368 43188 29420 43240
rect 24400 43052 24452 43104
rect 31116 43052 31168 43104
rect 31300 43052 31352 43104
rect 33048 43188 33100 43240
rect 36176 43231 36228 43240
rect 36176 43197 36185 43231
rect 36185 43197 36219 43231
rect 36219 43197 36228 43231
rect 36176 43188 36228 43197
rect 34336 43052 34388 43104
rect 37004 43052 37056 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 32950 42950 33002 43002
rect 33014 42950 33066 43002
rect 33078 42950 33130 43002
rect 33142 42950 33194 43002
rect 33206 42950 33258 43002
rect 42950 42950 43002 43002
rect 43014 42950 43066 43002
rect 43078 42950 43130 43002
rect 43142 42950 43194 43002
rect 43206 42950 43258 43002
rect 21640 42848 21692 42900
rect 13360 42780 13412 42832
rect 1308 42712 1360 42764
rect 17500 42644 17552 42696
rect 15108 42619 15160 42628
rect 15108 42585 15117 42619
rect 15117 42585 15151 42619
rect 15151 42585 15160 42619
rect 15108 42576 15160 42585
rect 16672 42576 16724 42628
rect 18604 42755 18656 42764
rect 18604 42721 18613 42755
rect 18613 42721 18647 42755
rect 18647 42721 18656 42755
rect 18604 42712 18656 42721
rect 20168 42780 20220 42832
rect 25044 42848 25096 42900
rect 26700 42891 26752 42900
rect 26700 42857 26709 42891
rect 26709 42857 26743 42891
rect 26743 42857 26752 42891
rect 26700 42848 26752 42857
rect 27528 42848 27580 42900
rect 29276 42848 29328 42900
rect 30564 42848 30616 42900
rect 30840 42848 30892 42900
rect 31484 42848 31536 42900
rect 25136 42780 25188 42832
rect 19432 42712 19484 42764
rect 19708 42712 19760 42764
rect 20536 42712 20588 42764
rect 22560 42712 22612 42764
rect 22836 42712 22888 42764
rect 23296 42755 23348 42764
rect 23296 42721 23305 42755
rect 23305 42721 23339 42755
rect 23339 42721 23348 42755
rect 23296 42712 23348 42721
rect 26608 42780 26660 42832
rect 25596 42712 25648 42764
rect 19524 42644 19576 42696
rect 19984 42644 20036 42696
rect 21824 42644 21876 42696
rect 16396 42508 16448 42560
rect 18972 42508 19024 42560
rect 20628 42576 20680 42628
rect 21088 42576 21140 42628
rect 23572 42644 23624 42696
rect 25044 42644 25096 42696
rect 26884 42687 26936 42696
rect 26884 42653 26893 42687
rect 26893 42653 26927 42687
rect 26927 42653 26936 42687
rect 26884 42644 26936 42653
rect 27436 42755 27488 42764
rect 27436 42721 27445 42755
rect 27445 42721 27479 42755
rect 27479 42721 27488 42755
rect 27436 42712 27488 42721
rect 29460 42712 29512 42764
rect 31944 42712 31996 42764
rect 32772 42712 32824 42764
rect 33600 42712 33652 42764
rect 36820 42848 36872 42900
rect 34888 42712 34940 42764
rect 36544 42644 36596 42696
rect 49056 42687 49108 42696
rect 49056 42653 49065 42687
rect 49065 42653 49099 42687
rect 49099 42653 49108 42687
rect 49056 42644 49108 42653
rect 21548 42508 21600 42560
rect 21916 42508 21968 42560
rect 23756 42508 23808 42560
rect 25044 42551 25096 42560
rect 25044 42517 25053 42551
rect 25053 42517 25087 42551
rect 25087 42517 25096 42551
rect 25044 42508 25096 42517
rect 27160 42508 27212 42560
rect 27528 42508 27580 42560
rect 29184 42551 29236 42560
rect 29184 42517 29193 42551
rect 29193 42517 29227 42551
rect 29227 42517 29236 42551
rect 29184 42508 29236 42517
rect 31668 42576 31720 42628
rect 32864 42576 32916 42628
rect 32404 42508 32456 42560
rect 33600 42508 33652 42560
rect 33692 42551 33744 42560
rect 33692 42517 33701 42551
rect 33701 42517 33735 42551
rect 33735 42517 33744 42551
rect 33692 42508 33744 42517
rect 33784 42508 33836 42560
rect 37832 42508 37884 42560
rect 47216 42508 47268 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 27950 42406 28002 42458
rect 28014 42406 28066 42458
rect 28078 42406 28130 42458
rect 28142 42406 28194 42458
rect 28206 42406 28258 42458
rect 37950 42406 38002 42458
rect 38014 42406 38066 42458
rect 38078 42406 38130 42458
rect 38142 42406 38194 42458
rect 38206 42406 38258 42458
rect 47950 42406 48002 42458
rect 48014 42406 48066 42458
rect 48078 42406 48130 42458
rect 48142 42406 48194 42458
rect 48206 42406 48258 42458
rect 11888 42347 11940 42356
rect 11888 42313 11897 42347
rect 11897 42313 11931 42347
rect 11931 42313 11940 42347
rect 11888 42304 11940 42313
rect 15108 42304 15160 42356
rect 24400 42304 24452 42356
rect 24952 42304 25004 42356
rect 27804 42304 27856 42356
rect 29644 42304 29696 42356
rect 16304 42211 16356 42220
rect 16304 42177 16313 42211
rect 16313 42177 16347 42211
rect 16347 42177 16356 42211
rect 16304 42168 16356 42177
rect 16856 42211 16908 42220
rect 16856 42177 16865 42211
rect 16865 42177 16899 42211
rect 16899 42177 16908 42211
rect 16856 42168 16908 42177
rect 17132 42143 17184 42152
rect 17132 42109 17141 42143
rect 17141 42109 17175 42143
rect 17175 42109 17184 42143
rect 17132 42100 17184 42109
rect 17684 42100 17736 42152
rect 18420 42236 18472 42288
rect 21824 42236 21876 42288
rect 22560 42236 22612 42288
rect 23572 42236 23624 42288
rect 27160 42279 27212 42288
rect 27160 42245 27169 42279
rect 27169 42245 27203 42279
rect 27203 42245 27212 42279
rect 27160 42236 27212 42245
rect 31484 42304 31536 42356
rect 31668 42347 31720 42356
rect 31668 42313 31677 42347
rect 31677 42313 31711 42347
rect 31711 42313 31720 42347
rect 31668 42304 31720 42313
rect 31852 42236 31904 42288
rect 32864 42304 32916 42356
rect 34244 42304 34296 42356
rect 32772 42236 32824 42288
rect 35164 42236 35216 42288
rect 36268 42236 36320 42288
rect 19248 42168 19300 42220
rect 20352 42168 20404 42220
rect 20536 42211 20588 42220
rect 20536 42177 20545 42211
rect 20545 42177 20579 42211
rect 20579 42177 20588 42211
rect 20536 42168 20588 42177
rect 26884 42168 26936 42220
rect 29552 42168 29604 42220
rect 35256 42168 35308 42220
rect 21916 42100 21968 42152
rect 24768 42100 24820 42152
rect 25136 42100 25188 42152
rect 27068 42100 27120 42152
rect 29276 42143 29328 42152
rect 29276 42109 29285 42143
rect 29285 42109 29319 42143
rect 29319 42109 29328 42143
rect 29276 42100 29328 42109
rect 16856 42032 16908 42084
rect 18328 42032 18380 42084
rect 20444 42032 20496 42084
rect 21088 42032 21140 42084
rect 21548 42032 21600 42084
rect 21824 42032 21876 42084
rect 29644 42032 29696 42084
rect 15292 41964 15344 42016
rect 20812 41964 20864 42016
rect 23756 42007 23808 42016
rect 23756 41973 23765 42007
rect 23765 41973 23799 42007
rect 23799 41973 23808 42007
rect 23756 41964 23808 41973
rect 24216 41964 24268 42016
rect 26608 41964 26660 42016
rect 31944 42100 31996 42152
rect 32864 42100 32916 42152
rect 36084 42100 36136 42152
rect 36636 42143 36688 42152
rect 36636 42109 36645 42143
rect 36645 42109 36679 42143
rect 36679 42109 36688 42143
rect 36636 42100 36688 42109
rect 31300 42032 31352 42084
rect 35164 41964 35216 42016
rect 39488 41964 39540 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 32950 41862 33002 41914
rect 33014 41862 33066 41914
rect 33078 41862 33130 41914
rect 33142 41862 33194 41914
rect 33206 41862 33258 41914
rect 42950 41862 43002 41914
rect 43014 41862 43066 41914
rect 43078 41862 43130 41914
rect 43142 41862 43194 41914
rect 43206 41862 43258 41914
rect 11980 41803 12032 41812
rect 11980 41769 11989 41803
rect 11989 41769 12023 41803
rect 12023 41769 12032 41803
rect 11980 41760 12032 41769
rect 13728 41760 13780 41812
rect 16304 41760 16356 41812
rect 21640 41760 21692 41812
rect 21916 41760 21968 41812
rect 9496 41692 9548 41744
rect 1308 41624 1360 41676
rect 11060 41556 11112 41608
rect 14280 41624 14332 41676
rect 16028 41624 16080 41676
rect 21180 41692 21232 41744
rect 24492 41760 24544 41812
rect 13360 41488 13412 41540
rect 16120 41488 16172 41540
rect 3608 41420 3660 41472
rect 20628 41624 20680 41676
rect 21272 41667 21324 41676
rect 21272 41633 21281 41667
rect 21281 41633 21315 41667
rect 21315 41633 21324 41667
rect 21272 41624 21324 41633
rect 23756 41692 23808 41744
rect 26608 41735 26660 41744
rect 26608 41701 26617 41735
rect 26617 41701 26651 41735
rect 26651 41701 26660 41735
rect 26608 41692 26660 41701
rect 27344 41692 27396 41744
rect 22468 41624 22520 41676
rect 23296 41624 23348 41676
rect 24584 41624 24636 41676
rect 25136 41624 25188 41676
rect 26424 41624 26476 41676
rect 18512 41556 18564 41608
rect 18880 41599 18932 41608
rect 18880 41565 18889 41599
rect 18889 41565 18923 41599
rect 18923 41565 18932 41599
rect 18880 41556 18932 41565
rect 21088 41556 21140 41608
rect 24124 41556 24176 41608
rect 17040 41463 17092 41472
rect 17040 41429 17049 41463
rect 17049 41429 17083 41463
rect 17083 41429 17092 41463
rect 17040 41420 17092 41429
rect 17592 41420 17644 41472
rect 22008 41488 22060 41540
rect 22560 41488 22612 41540
rect 23756 41488 23808 41540
rect 20996 41420 21048 41472
rect 22744 41420 22796 41472
rect 25412 41488 25464 41540
rect 25596 41488 25648 41540
rect 26976 41556 27028 41608
rect 27344 41556 27396 41608
rect 26608 41420 26660 41472
rect 30104 41760 30156 41812
rect 31484 41803 31536 41812
rect 31484 41769 31493 41803
rect 31493 41769 31527 41803
rect 31527 41769 31536 41803
rect 31484 41760 31536 41769
rect 32588 41760 32640 41812
rect 32956 41760 33008 41812
rect 33416 41760 33468 41812
rect 36544 41760 36596 41812
rect 36728 41760 36780 41812
rect 36912 41760 36964 41812
rect 29184 41692 29236 41744
rect 29460 41624 29512 41676
rect 30380 41624 30432 41676
rect 30656 41624 30708 41676
rect 29000 41599 29052 41608
rect 29000 41565 29009 41599
rect 29009 41565 29043 41599
rect 29043 41565 29052 41599
rect 29000 41556 29052 41565
rect 31944 41667 31996 41676
rect 31944 41633 31953 41667
rect 31953 41633 31987 41667
rect 31987 41633 31996 41667
rect 31944 41624 31996 41633
rect 33876 41624 33928 41676
rect 34336 41624 34388 41676
rect 34888 41667 34940 41676
rect 34888 41633 34897 41667
rect 34897 41633 34931 41667
rect 34931 41633 34940 41667
rect 34888 41624 34940 41633
rect 35164 41624 35216 41676
rect 36912 41624 36964 41676
rect 49056 41599 49108 41608
rect 49056 41565 49065 41599
rect 49065 41565 49099 41599
rect 49099 41565 49108 41599
rect 49056 41556 49108 41565
rect 31852 41488 31904 41540
rect 35256 41488 35308 41540
rect 36452 41488 36504 41540
rect 27804 41420 27856 41472
rect 29552 41420 29604 41472
rect 32312 41420 32364 41472
rect 36084 41420 36136 41472
rect 49240 41463 49292 41472
rect 49240 41429 49249 41463
rect 49249 41429 49283 41463
rect 49283 41429 49292 41463
rect 49240 41420 49292 41429
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 27950 41318 28002 41370
rect 28014 41318 28066 41370
rect 28078 41318 28130 41370
rect 28142 41318 28194 41370
rect 28206 41318 28258 41370
rect 37950 41318 38002 41370
rect 38014 41318 38066 41370
rect 38078 41318 38130 41370
rect 38142 41318 38194 41370
rect 38206 41318 38258 41370
rect 47950 41318 48002 41370
rect 48014 41318 48066 41370
rect 48078 41318 48130 41370
rect 48142 41318 48194 41370
rect 48206 41318 48258 41370
rect 11060 41216 11112 41268
rect 22100 41216 22152 41268
rect 18788 41148 18840 41200
rect 12256 41080 12308 41132
rect 19432 41148 19484 41200
rect 20444 41148 20496 41200
rect 21364 41148 21416 41200
rect 22008 41148 22060 41200
rect 23664 41216 23716 41268
rect 24768 41259 24820 41268
rect 24768 41225 24777 41259
rect 24777 41225 24811 41259
rect 24811 41225 24820 41259
rect 24768 41216 24820 41225
rect 25228 41259 25280 41268
rect 25228 41225 25237 41259
rect 25237 41225 25271 41259
rect 25271 41225 25280 41259
rect 25228 41216 25280 41225
rect 27712 41259 27764 41268
rect 27712 41225 27721 41259
rect 27721 41225 27755 41259
rect 27755 41225 27764 41259
rect 27712 41216 27764 41225
rect 29000 41216 29052 41268
rect 29736 41216 29788 41268
rect 28908 41148 28960 41200
rect 30840 41216 30892 41268
rect 1308 41012 1360 41064
rect 13820 40944 13872 40996
rect 15108 40944 15160 40996
rect 21088 41080 21140 41132
rect 18788 41012 18840 41064
rect 13544 40876 13596 40928
rect 20996 40944 21048 40996
rect 22376 41012 22428 41064
rect 23572 41080 23624 41132
rect 23296 40944 23348 40996
rect 23940 41012 23992 41064
rect 24032 41055 24084 41064
rect 24032 41021 24041 41055
rect 24041 41021 24075 41055
rect 24075 41021 24084 41055
rect 24032 41012 24084 41021
rect 24216 41055 24268 41064
rect 24216 41021 24225 41055
rect 24225 41021 24259 41055
rect 24259 41021 24268 41055
rect 24216 41012 24268 41021
rect 27712 41012 27764 41064
rect 28356 41080 28408 41132
rect 28448 41012 28500 41064
rect 28816 41012 28868 41064
rect 30840 41055 30892 41064
rect 30840 41021 30849 41055
rect 30849 41021 30883 41055
rect 30883 41021 30892 41055
rect 30840 41012 30892 41021
rect 31024 41012 31076 41064
rect 31392 41012 31444 41064
rect 24860 40944 24912 40996
rect 25504 40944 25556 40996
rect 29000 40944 29052 40996
rect 29184 40987 29236 40996
rect 29184 40953 29193 40987
rect 29193 40953 29227 40987
rect 29227 40953 29236 40987
rect 29184 40944 29236 40953
rect 33416 41216 33468 41268
rect 36544 41259 36596 41268
rect 36544 41225 36553 41259
rect 36553 41225 36587 41259
rect 36587 41225 36596 41259
rect 36544 41216 36596 41225
rect 32496 41080 32548 41132
rect 34244 41148 34296 41200
rect 35256 41148 35308 41200
rect 36084 41148 36136 41200
rect 33324 41080 33376 41132
rect 35440 41080 35492 41132
rect 37188 41080 37240 41132
rect 37280 41080 37332 41132
rect 38844 41080 38896 41132
rect 49332 41123 49384 41132
rect 49332 41089 49341 41123
rect 49341 41089 49375 41123
rect 49375 41089 49384 41123
rect 49332 41080 49384 41089
rect 32956 41055 33008 41064
rect 32956 41021 32965 41055
rect 32965 41021 32999 41055
rect 32999 41021 33008 41055
rect 32956 41012 33008 41021
rect 34520 41012 34572 41064
rect 35992 41012 36044 41064
rect 36728 41012 36780 41064
rect 37740 41055 37792 41064
rect 37740 41021 37749 41055
rect 37749 41021 37783 41055
rect 37783 41021 37792 41055
rect 37740 41012 37792 41021
rect 35072 40944 35124 40996
rect 20628 40919 20680 40928
rect 20628 40885 20637 40919
rect 20637 40885 20671 40919
rect 20671 40885 20680 40919
rect 20628 40876 20680 40885
rect 20904 40876 20956 40928
rect 22376 40876 22428 40928
rect 28356 40876 28408 40928
rect 28724 40876 28776 40928
rect 29736 40876 29788 40928
rect 31392 40876 31444 40928
rect 32496 40876 32548 40928
rect 34612 40876 34664 40928
rect 38752 40876 38804 40928
rect 39212 40919 39264 40928
rect 39212 40885 39221 40919
rect 39221 40885 39255 40919
rect 39255 40885 39264 40919
rect 39212 40876 39264 40885
rect 49148 40919 49200 40928
rect 49148 40885 49157 40919
rect 49157 40885 49191 40919
rect 49191 40885 49200 40919
rect 49148 40876 49200 40885
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 32950 40774 33002 40826
rect 33014 40774 33066 40826
rect 33078 40774 33130 40826
rect 33142 40774 33194 40826
rect 33206 40774 33258 40826
rect 42950 40774 43002 40826
rect 43014 40774 43066 40826
rect 43078 40774 43130 40826
rect 43142 40774 43194 40826
rect 43206 40774 43258 40826
rect 12256 40715 12308 40724
rect 12256 40681 12265 40715
rect 12265 40681 12299 40715
rect 12299 40681 12308 40715
rect 12256 40672 12308 40681
rect 17132 40672 17184 40724
rect 17868 40715 17920 40724
rect 17868 40681 17877 40715
rect 17877 40681 17911 40715
rect 17911 40681 17920 40715
rect 17868 40672 17920 40681
rect 19892 40672 19944 40724
rect 9588 40604 9640 40656
rect 20904 40672 20956 40724
rect 20996 40672 21048 40724
rect 23572 40672 23624 40724
rect 24952 40672 25004 40724
rect 29092 40672 29144 40724
rect 16948 40536 17000 40588
rect 17132 40536 17184 40588
rect 22100 40604 22152 40656
rect 25504 40604 25556 40656
rect 35072 40672 35124 40724
rect 15660 40511 15712 40520
rect 15660 40477 15669 40511
rect 15669 40477 15703 40511
rect 15703 40477 15712 40511
rect 15660 40468 15712 40477
rect 15936 40468 15988 40520
rect 19248 40468 19300 40520
rect 16028 40400 16080 40452
rect 16672 40400 16724 40452
rect 16856 40400 16908 40452
rect 18696 40400 18748 40452
rect 18420 40332 18472 40384
rect 20076 40536 20128 40588
rect 20536 40536 20588 40588
rect 22560 40536 22612 40588
rect 23848 40579 23900 40588
rect 23848 40545 23857 40579
rect 23857 40545 23891 40579
rect 23891 40545 23900 40579
rect 23848 40536 23900 40545
rect 27344 40579 27396 40588
rect 27344 40545 27353 40579
rect 27353 40545 27387 40579
rect 27387 40545 27396 40579
rect 27344 40536 27396 40545
rect 24308 40468 24360 40520
rect 20812 40400 20864 40452
rect 20904 40443 20956 40452
rect 20904 40409 20913 40443
rect 20913 40409 20947 40443
rect 20947 40409 20956 40443
rect 20904 40400 20956 40409
rect 21364 40400 21416 40452
rect 26240 40443 26292 40452
rect 26240 40409 26249 40443
rect 26249 40409 26283 40443
rect 26283 40409 26292 40443
rect 26240 40400 26292 40409
rect 29828 40604 29880 40656
rect 29368 40536 29420 40588
rect 29644 40536 29696 40588
rect 28632 40468 28684 40520
rect 30288 40579 30340 40588
rect 30288 40545 30297 40579
rect 30297 40545 30331 40579
rect 30331 40545 30340 40579
rect 30288 40536 30340 40545
rect 31484 40579 31536 40588
rect 31484 40545 31493 40579
rect 31493 40545 31527 40579
rect 31527 40545 31536 40579
rect 31484 40536 31536 40545
rect 34336 40604 34388 40656
rect 37096 40672 37148 40724
rect 37188 40672 37240 40724
rect 47400 40672 47452 40724
rect 32864 40536 32916 40588
rect 33324 40536 33376 40588
rect 37096 40536 37148 40588
rect 37648 40579 37700 40588
rect 37648 40545 37657 40579
rect 37657 40545 37691 40579
rect 37691 40545 37700 40579
rect 37648 40536 37700 40545
rect 37832 40536 37884 40588
rect 30564 40468 30616 40520
rect 30932 40468 30984 40520
rect 32404 40511 32456 40520
rect 32404 40477 32413 40511
rect 32413 40477 32447 40511
rect 32447 40477 32456 40511
rect 32404 40468 32456 40477
rect 32772 40468 32824 40520
rect 34520 40468 34572 40520
rect 35164 40511 35216 40520
rect 35164 40477 35173 40511
rect 35173 40477 35207 40511
rect 35207 40477 35216 40511
rect 35164 40468 35216 40477
rect 49148 40468 49200 40520
rect 20996 40332 21048 40384
rect 22468 40332 22520 40384
rect 25872 40332 25924 40384
rect 26424 40332 26476 40384
rect 28724 40332 28776 40384
rect 33692 40400 33744 40452
rect 30104 40332 30156 40384
rect 31760 40332 31812 40384
rect 33968 40332 34020 40384
rect 36084 40400 36136 40452
rect 39212 40400 39264 40452
rect 37648 40332 37700 40384
rect 47216 40400 47268 40452
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 27950 40230 28002 40282
rect 28014 40230 28066 40282
rect 28078 40230 28130 40282
rect 28142 40230 28194 40282
rect 28206 40230 28258 40282
rect 37950 40230 38002 40282
rect 38014 40230 38066 40282
rect 38078 40230 38130 40282
rect 38142 40230 38194 40282
rect 38206 40230 38258 40282
rect 47950 40230 48002 40282
rect 48014 40230 48066 40282
rect 48078 40230 48130 40282
rect 48142 40230 48194 40282
rect 48206 40230 48258 40282
rect 12808 40128 12860 40180
rect 17316 40128 17368 40180
rect 18880 40128 18932 40180
rect 8392 40060 8444 40112
rect 9312 40060 9364 40112
rect 9588 40060 9640 40112
rect 16856 40060 16908 40112
rect 17684 40060 17736 40112
rect 19524 40060 19576 40112
rect 20628 40128 20680 40180
rect 20812 40128 20864 40180
rect 21824 40128 21876 40180
rect 22284 40171 22336 40180
rect 22284 40137 22293 40171
rect 22293 40137 22327 40171
rect 22327 40137 22336 40171
rect 22284 40128 22336 40137
rect 23756 40128 23808 40180
rect 26700 40128 26752 40180
rect 27804 40128 27856 40180
rect 29736 40128 29788 40180
rect 31484 40128 31536 40180
rect 22468 40060 22520 40112
rect 22836 40060 22888 40112
rect 24952 40060 25004 40112
rect 25504 40060 25556 40112
rect 27436 40060 27488 40112
rect 14648 40035 14700 40044
rect 14648 40001 14657 40035
rect 14657 40001 14691 40035
rect 14691 40001 14700 40035
rect 14648 39992 14700 40001
rect 15476 39992 15528 40044
rect 16304 39992 16356 40044
rect 2044 39967 2096 39976
rect 2044 39933 2053 39967
rect 2053 39933 2087 39967
rect 2087 39933 2096 39967
rect 2044 39924 2096 39933
rect 14924 39967 14976 39976
rect 14924 39933 14933 39967
rect 14933 39933 14967 39967
rect 14967 39933 14976 39967
rect 14924 39924 14976 39933
rect 19432 39992 19484 40044
rect 20996 39992 21048 40044
rect 21364 39992 21416 40044
rect 21732 39992 21784 40044
rect 3332 39856 3384 39908
rect 18788 39967 18840 39976
rect 18788 39933 18797 39967
rect 18797 39933 18831 39967
rect 18831 39933 18840 39967
rect 18788 39924 18840 39933
rect 19616 39967 19668 39976
rect 19616 39933 19625 39967
rect 19625 39933 19659 39967
rect 19659 39933 19668 39967
rect 19616 39924 19668 39933
rect 17684 39856 17736 39908
rect 22192 39924 22244 39976
rect 22560 39924 22612 39976
rect 24584 40035 24636 40044
rect 24584 40001 24593 40035
rect 24593 40001 24627 40035
rect 24627 40001 24636 40035
rect 24584 39992 24636 40001
rect 23756 39856 23808 39908
rect 7564 39788 7616 39840
rect 12716 39788 12768 39840
rect 14372 39788 14424 39840
rect 22744 39788 22796 39840
rect 23940 39788 23992 39840
rect 24492 39788 24544 39840
rect 26884 39924 26936 39976
rect 27344 39924 27396 39976
rect 30656 40060 30708 40112
rect 31760 40060 31812 40112
rect 31116 39992 31168 40044
rect 26516 39856 26568 39908
rect 30196 39924 30248 39976
rect 31576 39967 31628 39976
rect 31576 39933 31585 39967
rect 31585 39933 31619 39967
rect 31619 39933 31628 39967
rect 31576 39924 31628 39933
rect 25964 39788 26016 39840
rect 34428 40128 34480 40180
rect 35440 40128 35492 40180
rect 36176 40128 36228 40180
rect 38752 40128 38804 40180
rect 32864 40060 32916 40112
rect 33876 40060 33928 40112
rect 35256 40060 35308 40112
rect 32312 40035 32364 40044
rect 32312 40001 32321 40035
rect 32321 40001 32355 40035
rect 32355 40001 32364 40035
rect 32312 39992 32364 40001
rect 34520 40035 34572 40044
rect 34520 40001 34529 40035
rect 34529 40001 34563 40035
rect 34563 40001 34572 40035
rect 34520 39992 34572 40001
rect 33600 39924 33652 39976
rect 33876 39924 33928 39976
rect 34428 39924 34480 39976
rect 35348 39924 35400 39976
rect 39120 40035 39172 40044
rect 39120 40001 39129 40035
rect 39129 40001 39163 40035
rect 39163 40001 39172 40035
rect 39120 39992 39172 40001
rect 49056 40035 49108 40044
rect 49056 40001 49065 40035
rect 49065 40001 49099 40035
rect 49099 40001 49108 40035
rect 49056 39992 49108 40001
rect 27160 39831 27212 39840
rect 27160 39797 27169 39831
rect 27169 39797 27203 39831
rect 27203 39797 27212 39831
rect 27160 39788 27212 39797
rect 27804 39788 27856 39840
rect 28908 39788 28960 39840
rect 34060 39831 34112 39840
rect 34060 39797 34069 39831
rect 34069 39797 34103 39831
rect 34103 39797 34112 39831
rect 34060 39788 34112 39797
rect 37556 39788 37608 39840
rect 38476 39788 38528 39840
rect 39396 39924 39448 39976
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 32950 39686 33002 39738
rect 33014 39686 33066 39738
rect 33078 39686 33130 39738
rect 33142 39686 33194 39738
rect 33206 39686 33258 39738
rect 42950 39686 43002 39738
rect 43014 39686 43066 39738
rect 43078 39686 43130 39738
rect 43142 39686 43194 39738
rect 43206 39686 43258 39738
rect 1676 39584 1728 39636
rect 7564 39584 7616 39636
rect 14648 39584 14700 39636
rect 16672 39584 16724 39636
rect 17776 39584 17828 39636
rect 14464 39448 14516 39500
rect 15936 39448 15988 39500
rect 16304 39448 16356 39500
rect 21548 39516 21600 39568
rect 21732 39584 21784 39636
rect 22468 39584 22520 39636
rect 24400 39584 24452 39636
rect 25044 39584 25096 39636
rect 25872 39627 25924 39636
rect 25872 39593 25881 39627
rect 25881 39593 25915 39627
rect 25915 39593 25924 39627
rect 25872 39584 25924 39593
rect 28632 39584 28684 39636
rect 29092 39627 29144 39636
rect 29092 39593 29101 39627
rect 29101 39593 29135 39627
rect 29135 39593 29144 39627
rect 29092 39584 29144 39593
rect 30012 39584 30064 39636
rect 31760 39584 31812 39636
rect 31944 39584 31996 39636
rect 34060 39584 34112 39636
rect 23020 39559 23072 39568
rect 23020 39525 23029 39559
rect 23029 39525 23063 39559
rect 23063 39525 23072 39559
rect 23020 39516 23072 39525
rect 12716 39423 12768 39432
rect 12716 39389 12725 39423
rect 12725 39389 12759 39423
rect 12759 39389 12768 39423
rect 12716 39380 12768 39389
rect 13636 39380 13688 39432
rect 17868 39380 17920 39432
rect 20904 39448 20956 39500
rect 21456 39491 21508 39500
rect 21456 39457 21465 39491
rect 21465 39457 21499 39491
rect 21499 39457 21508 39491
rect 21456 39448 21508 39457
rect 22652 39448 22704 39500
rect 25136 39491 25188 39500
rect 25136 39457 25145 39491
rect 25145 39457 25179 39491
rect 25179 39457 25188 39491
rect 25136 39448 25188 39457
rect 26884 39448 26936 39500
rect 27068 39448 27120 39500
rect 28632 39448 28684 39500
rect 25412 39380 25464 39432
rect 28954 39448 29006 39500
rect 32772 39516 32824 39568
rect 29828 39380 29880 39432
rect 1308 39312 1360 39364
rect 12624 39244 12676 39296
rect 15844 39312 15896 39364
rect 16212 39312 16264 39364
rect 18696 39312 18748 39364
rect 16580 39244 16632 39296
rect 16856 39244 16908 39296
rect 18604 39287 18656 39296
rect 18604 39253 18613 39287
rect 18613 39253 18647 39287
rect 18647 39253 18656 39287
rect 18604 39244 18656 39253
rect 22744 39312 22796 39364
rect 23296 39312 23348 39364
rect 26976 39312 27028 39364
rect 27620 39355 27672 39364
rect 27620 39321 27629 39355
rect 27629 39321 27663 39355
rect 27663 39321 27672 39355
rect 27620 39312 27672 39321
rect 28632 39312 28684 39364
rect 28908 39312 28960 39364
rect 32312 39448 32364 39500
rect 33692 39448 33744 39500
rect 34060 39448 34112 39500
rect 34336 39516 34388 39568
rect 37372 39584 37424 39636
rect 39304 39584 39356 39636
rect 33140 39380 33192 39432
rect 34888 39448 34940 39500
rect 35348 39448 35400 39500
rect 41328 39516 41380 39568
rect 38936 39448 38988 39500
rect 39212 39448 39264 39500
rect 34520 39380 34572 39432
rect 20168 39287 20220 39296
rect 20168 39253 20177 39287
rect 20177 39253 20211 39287
rect 20211 39253 20220 39287
rect 20168 39244 20220 39253
rect 20904 39287 20956 39296
rect 20904 39253 20913 39287
rect 20913 39253 20947 39287
rect 20947 39253 20956 39287
rect 20904 39244 20956 39253
rect 22468 39244 22520 39296
rect 22652 39244 22704 39296
rect 26056 39244 26108 39296
rect 26332 39287 26384 39296
rect 26332 39253 26341 39287
rect 26341 39253 26375 39287
rect 26375 39253 26384 39287
rect 26332 39244 26384 39253
rect 27252 39244 27304 39296
rect 29920 39244 29972 39296
rect 31760 39244 31812 39296
rect 33416 39312 33468 39364
rect 34152 39312 34204 39364
rect 49240 39380 49292 39432
rect 35164 39312 35216 39364
rect 35256 39355 35308 39364
rect 35256 39321 35265 39355
rect 35265 39321 35299 39355
rect 35299 39321 35308 39355
rect 35256 39312 35308 39321
rect 36268 39312 36320 39364
rect 32312 39244 32364 39296
rect 33600 39287 33652 39296
rect 33600 39253 33609 39287
rect 33609 39253 33643 39287
rect 33643 39253 33652 39287
rect 33600 39244 33652 39253
rect 33968 39287 34020 39296
rect 33968 39253 33977 39287
rect 33977 39253 34011 39287
rect 34011 39253 34020 39287
rect 33968 39244 34020 39253
rect 36084 39244 36136 39296
rect 36912 39244 36964 39296
rect 37464 39355 37516 39364
rect 37464 39321 37473 39355
rect 37473 39321 37507 39355
rect 37507 39321 37516 39355
rect 37464 39312 37516 39321
rect 39120 39312 39172 39364
rect 39304 39355 39356 39364
rect 39304 39321 39313 39355
rect 39313 39321 39347 39355
rect 39347 39321 39356 39355
rect 39304 39312 39356 39321
rect 49148 39355 49200 39364
rect 49148 39321 49157 39355
rect 49157 39321 49191 39355
rect 49191 39321 49200 39355
rect 49148 39312 49200 39321
rect 38476 39287 38528 39296
rect 38476 39253 38485 39287
rect 38485 39253 38519 39287
rect 38519 39253 38528 39287
rect 38476 39244 38528 39253
rect 39212 39287 39264 39296
rect 39212 39253 39221 39287
rect 39221 39253 39255 39287
rect 39255 39253 39264 39287
rect 39212 39244 39264 39253
rect 49240 39287 49292 39296
rect 49240 39253 49249 39287
rect 49249 39253 49283 39287
rect 49283 39253 49292 39287
rect 49240 39244 49292 39253
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 27950 39142 28002 39194
rect 28014 39142 28066 39194
rect 28078 39142 28130 39194
rect 28142 39142 28194 39194
rect 28206 39142 28258 39194
rect 37950 39142 38002 39194
rect 38014 39142 38066 39194
rect 38078 39142 38130 39194
rect 38142 39142 38194 39194
rect 38206 39142 38258 39194
rect 47950 39142 48002 39194
rect 48014 39142 48066 39194
rect 48078 39142 48130 39194
rect 48142 39142 48194 39194
rect 48206 39142 48258 39194
rect 15016 39040 15068 39092
rect 15660 39040 15712 39092
rect 16948 39083 17000 39092
rect 16948 39049 16957 39083
rect 16957 39049 16991 39083
rect 16991 39049 17000 39083
rect 16948 39040 17000 39049
rect 17316 39083 17368 39092
rect 17316 39049 17325 39083
rect 17325 39049 17359 39083
rect 17359 39049 17368 39083
rect 17316 39040 17368 39049
rect 17776 39040 17828 39092
rect 18420 39083 18472 39092
rect 18420 39049 18429 39083
rect 18429 39049 18463 39083
rect 18463 39049 18472 39083
rect 18420 39040 18472 39049
rect 14648 38972 14700 39024
rect 17132 38972 17184 39024
rect 19340 38972 19392 39024
rect 17684 38904 17736 38956
rect 18328 38947 18380 38956
rect 18328 38913 18337 38947
rect 18337 38913 18371 38947
rect 18371 38913 18380 38947
rect 18328 38904 18380 38913
rect 16028 38836 16080 38888
rect 16120 38879 16172 38888
rect 16120 38845 16129 38879
rect 16129 38845 16163 38879
rect 16163 38845 16172 38879
rect 16120 38836 16172 38845
rect 19524 38904 19576 38956
rect 19616 38904 19668 38956
rect 20996 38972 21048 39024
rect 21456 39083 21508 39092
rect 21456 39049 21465 39083
rect 21465 39049 21499 39083
rect 21499 39049 21508 39083
rect 21456 39040 21508 39049
rect 21548 39040 21600 39092
rect 23756 39083 23808 39092
rect 23756 39049 23765 39083
rect 23765 39049 23799 39083
rect 23799 39049 23808 39083
rect 23756 39040 23808 39049
rect 24032 39040 24084 39092
rect 24676 39083 24728 39092
rect 24676 39049 24685 39083
rect 24685 39049 24719 39083
rect 24719 39049 24728 39083
rect 24676 39040 24728 39049
rect 26332 39040 26384 39092
rect 27620 39040 27672 39092
rect 21364 38972 21416 39024
rect 22744 38972 22796 39024
rect 21456 38904 21508 38956
rect 16212 38768 16264 38820
rect 21548 38836 21600 38888
rect 21824 38768 21876 38820
rect 25780 38972 25832 39024
rect 24584 38947 24636 38956
rect 24584 38913 24593 38947
rect 24593 38913 24627 38947
rect 24627 38913 24636 38947
rect 24584 38904 24636 38913
rect 27804 38972 27856 39024
rect 30196 39083 30248 39092
rect 30196 39049 30205 39083
rect 30205 39049 30239 39083
rect 30239 39049 30248 39083
rect 30196 39040 30248 39049
rect 31300 39040 31352 39092
rect 31760 39040 31812 39092
rect 30932 38972 30984 39024
rect 31576 38972 31628 39024
rect 31852 38972 31904 39024
rect 33600 39040 33652 39092
rect 35256 39040 35308 39092
rect 37832 39040 37884 39092
rect 38660 39040 38712 39092
rect 34612 38972 34664 39024
rect 36176 38972 36228 39024
rect 37648 38972 37700 39024
rect 27252 38904 27304 38956
rect 15108 38700 15160 38752
rect 15844 38700 15896 38752
rect 21088 38700 21140 38752
rect 24768 38879 24820 38888
rect 24768 38845 24777 38879
rect 24777 38845 24811 38879
rect 24811 38845 24820 38879
rect 24768 38836 24820 38845
rect 27344 38836 27396 38888
rect 29828 38904 29880 38956
rect 30656 38904 30708 38956
rect 32220 38904 32272 38956
rect 33600 38904 33652 38956
rect 33968 38904 34020 38956
rect 35164 38947 35216 38956
rect 35164 38913 35173 38947
rect 35173 38913 35207 38947
rect 35207 38913 35216 38947
rect 35164 38904 35216 38913
rect 38108 38947 38160 38956
rect 38108 38913 38117 38947
rect 38117 38913 38151 38947
rect 38151 38913 38160 38947
rect 38108 38904 38160 38913
rect 39304 38904 39356 38956
rect 49240 38904 49292 38956
rect 28448 38879 28500 38888
rect 28448 38845 28457 38879
rect 28457 38845 28491 38879
rect 28491 38845 28500 38879
rect 28448 38836 28500 38845
rect 29184 38836 29236 38888
rect 29276 38836 29328 38888
rect 32680 38836 32732 38888
rect 24492 38768 24544 38820
rect 24584 38700 24636 38752
rect 24768 38700 24820 38752
rect 26240 38700 26292 38752
rect 27344 38700 27396 38752
rect 33140 38768 33192 38820
rect 33692 38836 33744 38888
rect 33876 38836 33928 38888
rect 35440 38879 35492 38888
rect 35440 38845 35449 38879
rect 35449 38845 35483 38879
rect 35483 38845 35492 38879
rect 35440 38836 35492 38845
rect 36912 38836 36964 38888
rect 35072 38768 35124 38820
rect 29920 38700 29972 38752
rect 38844 38768 38896 38820
rect 38660 38743 38712 38752
rect 38660 38709 38669 38743
rect 38669 38709 38703 38743
rect 38703 38709 38712 38743
rect 38660 38700 38712 38709
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 32950 38598 33002 38650
rect 33014 38598 33066 38650
rect 33078 38598 33130 38650
rect 33142 38598 33194 38650
rect 33206 38598 33258 38650
rect 42950 38598 43002 38650
rect 43014 38598 43066 38650
rect 43078 38598 43130 38650
rect 43142 38598 43194 38650
rect 43206 38598 43258 38650
rect 8392 38539 8444 38548
rect 8392 38505 8401 38539
rect 8401 38505 8435 38539
rect 8435 38505 8444 38539
rect 8392 38496 8444 38505
rect 12440 38539 12492 38548
rect 12440 38505 12449 38539
rect 12449 38505 12483 38539
rect 12483 38505 12492 38539
rect 12440 38496 12492 38505
rect 12716 38496 12768 38548
rect 14372 38496 14424 38548
rect 1768 38428 1820 38480
rect 17868 38496 17920 38548
rect 18972 38496 19024 38548
rect 20168 38496 20220 38548
rect 21272 38496 21324 38548
rect 24952 38496 25004 38548
rect 25688 38496 25740 38548
rect 1308 38360 1360 38412
rect 16212 38471 16264 38480
rect 16212 38437 16221 38471
rect 16221 38437 16255 38471
rect 16255 38437 16264 38471
rect 16212 38428 16264 38437
rect 17040 38428 17092 38480
rect 20076 38428 20128 38480
rect 12716 38292 12768 38344
rect 12808 38292 12860 38344
rect 14464 38403 14516 38412
rect 14464 38369 14473 38403
rect 14473 38369 14507 38403
rect 14507 38369 14516 38403
rect 14464 38360 14516 38369
rect 18880 38360 18932 38412
rect 21824 38428 21876 38480
rect 22744 38403 22796 38412
rect 22744 38369 22753 38403
rect 22753 38369 22787 38403
rect 22787 38369 22796 38403
rect 22744 38360 22796 38369
rect 16856 38292 16908 38344
rect 19432 38292 19484 38344
rect 19984 38335 20036 38344
rect 19984 38301 19993 38335
rect 19993 38301 20027 38335
rect 20027 38301 20036 38335
rect 19984 38292 20036 38301
rect 21732 38292 21784 38344
rect 25596 38428 25648 38480
rect 28540 38496 28592 38548
rect 24676 38360 24728 38412
rect 25780 38403 25832 38412
rect 25780 38369 25789 38403
rect 25789 38369 25823 38403
rect 25823 38369 25832 38403
rect 25780 38360 25832 38369
rect 26884 38360 26936 38412
rect 27160 38292 27212 38344
rect 27436 38360 27488 38412
rect 29644 38428 29696 38480
rect 32128 38496 32180 38548
rect 39212 38496 39264 38548
rect 31944 38360 31996 38412
rect 35440 38360 35492 38412
rect 36820 38403 36872 38412
rect 36820 38369 36829 38403
rect 36829 38369 36863 38403
rect 36863 38369 36872 38403
rect 36820 38360 36872 38369
rect 37740 38360 37792 38412
rect 39672 38428 39724 38480
rect 38936 38403 38988 38412
rect 38936 38369 38945 38403
rect 38945 38369 38979 38403
rect 38979 38369 38988 38403
rect 38936 38360 38988 38369
rect 12900 38156 12952 38208
rect 14832 38224 14884 38276
rect 16672 38224 16724 38276
rect 15108 38156 15160 38208
rect 17408 38199 17460 38208
rect 17408 38165 17417 38199
rect 17417 38165 17451 38199
rect 17451 38165 17460 38199
rect 17408 38156 17460 38165
rect 18604 38224 18656 38276
rect 21456 38267 21508 38276
rect 21456 38233 21465 38267
rect 21465 38233 21499 38267
rect 21499 38233 21508 38267
rect 21456 38224 21508 38233
rect 20904 38156 20956 38208
rect 22560 38199 22612 38208
rect 22560 38165 22569 38199
rect 22569 38165 22603 38199
rect 22603 38165 22612 38199
rect 22560 38156 22612 38165
rect 23296 38224 23348 38276
rect 23572 38156 23624 38208
rect 23664 38199 23716 38208
rect 23664 38165 23673 38199
rect 23673 38165 23707 38199
rect 23707 38165 23716 38199
rect 23664 38156 23716 38165
rect 25320 38156 25372 38208
rect 25688 38156 25740 38208
rect 26424 38224 26476 38276
rect 27620 38224 27672 38276
rect 28448 38292 28500 38344
rect 32220 38335 32272 38344
rect 32220 38301 32229 38335
rect 32229 38301 32263 38335
rect 32263 38301 32272 38335
rect 32220 38292 32272 38301
rect 27436 38199 27488 38208
rect 27436 38165 27445 38199
rect 27445 38165 27479 38199
rect 27479 38165 27488 38199
rect 27436 38156 27488 38165
rect 31300 38224 31352 38276
rect 31576 38224 31628 38276
rect 31484 38199 31536 38208
rect 31484 38165 31493 38199
rect 31493 38165 31527 38199
rect 31527 38165 31536 38199
rect 36636 38292 36688 38344
rect 38660 38292 38712 38344
rect 31484 38156 31536 38165
rect 33416 38199 33468 38208
rect 33416 38165 33425 38199
rect 33425 38165 33459 38199
rect 33459 38165 33468 38199
rect 33416 38156 33468 38165
rect 33876 38156 33928 38208
rect 34244 38156 34296 38208
rect 34888 38267 34940 38276
rect 34888 38233 34897 38267
rect 34897 38233 34931 38267
rect 34931 38233 34940 38267
rect 34888 38224 34940 38233
rect 35164 38224 35216 38276
rect 36176 38224 36228 38276
rect 36452 38156 36504 38208
rect 36636 38199 36688 38208
rect 36636 38165 36645 38199
rect 36645 38165 36679 38199
rect 36679 38165 36688 38199
rect 36636 38156 36688 38165
rect 36728 38199 36780 38208
rect 36728 38165 36737 38199
rect 36737 38165 36771 38199
rect 36771 38165 36780 38199
rect 36728 38156 36780 38165
rect 38844 38224 38896 38276
rect 49148 38267 49200 38276
rect 49148 38233 49157 38267
rect 49157 38233 49191 38267
rect 49191 38233 49200 38267
rect 49148 38224 49200 38233
rect 49240 38199 49292 38208
rect 49240 38165 49249 38199
rect 49249 38165 49283 38199
rect 49283 38165 49292 38199
rect 49240 38156 49292 38165
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 27950 38054 28002 38106
rect 28014 38054 28066 38106
rect 28078 38054 28130 38106
rect 28142 38054 28194 38106
rect 28206 38054 28258 38106
rect 37950 38054 38002 38106
rect 38014 38054 38066 38106
rect 38078 38054 38130 38106
rect 38142 38054 38194 38106
rect 38206 38054 38258 38106
rect 47950 38054 48002 38106
rect 48014 38054 48066 38106
rect 48078 38054 48130 38106
rect 48142 38054 48194 38106
rect 48206 38054 48258 38106
rect 15200 37952 15252 38004
rect 18512 37952 18564 38004
rect 20720 37995 20772 38004
rect 20720 37961 20729 37995
rect 20729 37961 20763 37995
rect 20763 37961 20772 37995
rect 20720 37952 20772 37961
rect 16672 37884 16724 37936
rect 1768 37859 1820 37868
rect 1768 37825 1777 37859
rect 1777 37825 1811 37859
rect 1811 37825 1820 37859
rect 1768 37816 1820 37825
rect 12900 37816 12952 37868
rect 14464 37816 14516 37868
rect 21640 37952 21692 38004
rect 22560 37952 22612 38004
rect 21548 37884 21600 37936
rect 26240 37884 26292 37936
rect 28448 37952 28500 38004
rect 28816 37952 28868 38004
rect 30932 37952 30984 38004
rect 28172 37884 28224 37936
rect 20996 37816 21048 37868
rect 21456 37816 21508 37868
rect 22008 37859 22060 37868
rect 22008 37825 22017 37859
rect 22017 37825 22051 37859
rect 22051 37825 22060 37859
rect 22008 37816 22060 37825
rect 23388 37816 23440 37868
rect 23756 37816 23808 37868
rect 24768 37816 24820 37868
rect 24860 37859 24912 37868
rect 24860 37825 24869 37859
rect 24869 37825 24903 37859
rect 24903 37825 24912 37859
rect 24860 37816 24912 37825
rect 25872 37816 25924 37868
rect 27160 37859 27212 37868
rect 27160 37825 27169 37859
rect 27169 37825 27203 37859
rect 27203 37825 27212 37859
rect 27160 37816 27212 37825
rect 29920 37884 29972 37936
rect 31300 37884 31352 37936
rect 32036 37816 32088 37868
rect 35164 37952 35216 38004
rect 36728 37952 36780 38004
rect 39120 37995 39172 38004
rect 39120 37961 39129 37995
rect 39129 37961 39163 37995
rect 39163 37961 39172 37995
rect 39120 37952 39172 37961
rect 34428 37884 34480 37936
rect 36452 37884 36504 37936
rect 1308 37748 1360 37800
rect 16120 37748 16172 37800
rect 19340 37748 19392 37800
rect 19432 37791 19484 37800
rect 19432 37757 19441 37791
rect 19441 37757 19475 37791
rect 19475 37757 19484 37791
rect 19432 37748 19484 37757
rect 19524 37791 19576 37800
rect 19524 37757 19533 37791
rect 19533 37757 19567 37791
rect 19567 37757 19576 37791
rect 19524 37748 19576 37757
rect 20444 37748 20496 37800
rect 20076 37680 20128 37732
rect 8576 37655 8628 37664
rect 8576 37621 8585 37655
rect 8585 37621 8619 37655
rect 8619 37621 8628 37655
rect 8576 37612 8628 37621
rect 13820 37612 13872 37664
rect 14924 37612 14976 37664
rect 16488 37612 16540 37664
rect 25044 37791 25096 37800
rect 25044 37757 25053 37791
rect 25053 37757 25087 37791
rect 25087 37757 25096 37791
rect 25044 37748 25096 37757
rect 25228 37748 25280 37800
rect 23388 37680 23440 37732
rect 23480 37680 23532 37732
rect 23848 37612 23900 37664
rect 25872 37680 25924 37732
rect 27068 37748 27120 37800
rect 28172 37748 28224 37800
rect 28632 37748 28684 37800
rect 31852 37748 31904 37800
rect 33784 37748 33836 37800
rect 31116 37612 31168 37664
rect 35440 37748 35492 37800
rect 37004 37816 37056 37868
rect 35716 37791 35768 37800
rect 35716 37757 35725 37791
rect 35725 37757 35759 37791
rect 35759 37757 35768 37791
rect 35716 37748 35768 37757
rect 35808 37791 35860 37800
rect 35808 37757 35817 37791
rect 35817 37757 35851 37791
rect 35851 37757 35860 37791
rect 35808 37748 35860 37757
rect 37832 37748 37884 37800
rect 49240 37884 49292 37936
rect 38568 37748 38620 37800
rect 49332 37859 49384 37868
rect 49332 37825 49341 37859
rect 49341 37825 49375 37859
rect 49375 37825 49384 37859
rect 49332 37816 49384 37825
rect 34244 37655 34296 37664
rect 34244 37621 34253 37655
rect 34253 37621 34287 37655
rect 34287 37621 34296 37655
rect 34244 37612 34296 37621
rect 34704 37655 34756 37664
rect 34704 37621 34713 37655
rect 34713 37621 34747 37655
rect 34747 37621 34756 37655
rect 34704 37612 34756 37621
rect 35716 37612 35768 37664
rect 39856 37612 39908 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 32950 37510 33002 37562
rect 33014 37510 33066 37562
rect 33078 37510 33130 37562
rect 33142 37510 33194 37562
rect 33206 37510 33258 37562
rect 42950 37510 43002 37562
rect 43014 37510 43066 37562
rect 43078 37510 43130 37562
rect 43142 37510 43194 37562
rect 43206 37510 43258 37562
rect 14372 37408 14424 37460
rect 12992 37272 13044 37324
rect 12532 37204 12584 37256
rect 14648 37272 14700 37324
rect 15108 37315 15160 37324
rect 15108 37281 15117 37315
rect 15117 37281 15151 37315
rect 15151 37281 15160 37315
rect 15108 37272 15160 37281
rect 16212 37272 16264 37324
rect 18420 37272 18472 37324
rect 20996 37408 21048 37460
rect 18880 37340 18932 37392
rect 28264 37408 28316 37460
rect 31116 37408 31168 37460
rect 31300 37408 31352 37460
rect 19248 37272 19300 37324
rect 22376 37272 22428 37324
rect 23940 37272 23992 37324
rect 24032 37272 24084 37324
rect 27068 37272 27120 37324
rect 28356 37272 28408 37324
rect 13912 37204 13964 37256
rect 14464 37204 14516 37256
rect 15844 37247 15896 37256
rect 15844 37213 15853 37247
rect 15853 37213 15887 37247
rect 15887 37213 15896 37247
rect 15844 37204 15896 37213
rect 17592 37204 17644 37256
rect 23296 37204 23348 37256
rect 27620 37204 27672 37256
rect 5356 37136 5408 37188
rect 15752 37136 15804 37188
rect 16672 37136 16724 37188
rect 19892 37136 19944 37188
rect 14740 37068 14792 37120
rect 15016 37068 15068 37120
rect 16212 37068 16264 37120
rect 17684 37068 17736 37120
rect 18788 37068 18840 37120
rect 19800 37068 19852 37120
rect 21732 37068 21784 37120
rect 26056 37136 26108 37188
rect 27528 37136 27580 37188
rect 30012 37272 30064 37324
rect 30932 37315 30984 37324
rect 30932 37281 30941 37315
rect 30941 37281 30975 37315
rect 30975 37281 30984 37315
rect 30932 37272 30984 37281
rect 33416 37408 33468 37460
rect 29920 37204 29972 37256
rect 30472 37136 30524 37188
rect 23296 37111 23348 37120
rect 23296 37077 23305 37111
rect 23305 37077 23339 37111
rect 23339 37077 23348 37111
rect 23296 37068 23348 37077
rect 26240 37111 26292 37120
rect 26240 37077 26249 37111
rect 26249 37077 26283 37111
rect 26283 37077 26292 37111
rect 26240 37068 26292 37077
rect 26516 37068 26568 37120
rect 30380 37068 30432 37120
rect 32312 37204 32364 37256
rect 33324 37272 33376 37324
rect 36820 37272 36872 37324
rect 36912 37272 36964 37324
rect 33140 37204 33192 37256
rect 34152 37204 34204 37256
rect 37648 37204 37700 37256
rect 32312 37068 32364 37120
rect 32772 37136 32824 37188
rect 33416 37136 33468 37188
rect 36360 37136 36412 37188
rect 32496 37068 32548 37120
rect 35808 37068 35860 37120
rect 38660 37136 38712 37188
rect 39396 37136 39448 37188
rect 37556 37111 37608 37120
rect 37556 37077 37565 37111
rect 37565 37077 37599 37111
rect 37599 37077 37608 37111
rect 37556 37068 37608 37077
rect 37648 37068 37700 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 27950 36966 28002 37018
rect 28014 36966 28066 37018
rect 28078 36966 28130 37018
rect 28142 36966 28194 37018
rect 28206 36966 28258 37018
rect 37950 36966 38002 37018
rect 38014 36966 38066 37018
rect 38078 36966 38130 37018
rect 38142 36966 38194 37018
rect 38206 36966 38258 37018
rect 47950 36966 48002 37018
rect 48014 36966 48066 37018
rect 48078 36966 48130 37018
rect 48142 36966 48194 37018
rect 48206 36966 48258 37018
rect 12716 36864 12768 36916
rect 13452 36864 13504 36916
rect 14464 36864 14516 36916
rect 18512 36864 18564 36916
rect 19064 36864 19116 36916
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 4896 36728 4948 36780
rect 5356 36728 5408 36780
rect 13452 36728 13504 36780
rect 13820 36839 13872 36848
rect 13820 36805 13829 36839
rect 13829 36805 13863 36839
rect 13863 36805 13872 36839
rect 13820 36796 13872 36805
rect 14924 36728 14976 36780
rect 16672 36796 16724 36848
rect 19616 36864 19668 36916
rect 22192 36864 22244 36916
rect 26240 36864 26292 36916
rect 16764 36728 16816 36780
rect 18512 36728 18564 36780
rect 20812 36796 20864 36848
rect 22008 36796 22060 36848
rect 21824 36728 21876 36780
rect 24400 36796 24452 36848
rect 1308 36660 1360 36712
rect 12992 36703 13044 36712
rect 12992 36669 13001 36703
rect 13001 36669 13035 36703
rect 13035 36669 13044 36703
rect 12992 36660 13044 36669
rect 13360 36660 13412 36712
rect 15844 36660 15896 36712
rect 16856 36703 16908 36712
rect 16856 36669 16865 36703
rect 16865 36669 16899 36703
rect 16899 36669 16908 36703
rect 16856 36660 16908 36669
rect 17132 36703 17184 36712
rect 17132 36669 17141 36703
rect 17141 36669 17175 36703
rect 17175 36669 17184 36703
rect 17132 36660 17184 36669
rect 19248 36660 19300 36712
rect 19800 36660 19852 36712
rect 21180 36703 21232 36712
rect 21180 36669 21189 36703
rect 21189 36669 21223 36703
rect 21223 36669 21232 36703
rect 21180 36660 21232 36669
rect 21364 36703 21416 36712
rect 21364 36669 21373 36703
rect 21373 36669 21407 36703
rect 21407 36669 21416 36703
rect 21364 36660 21416 36669
rect 22652 36703 22704 36712
rect 22652 36669 22661 36703
rect 22661 36669 22695 36703
rect 22695 36669 22704 36703
rect 22652 36660 22704 36669
rect 22744 36660 22796 36712
rect 23848 36703 23900 36712
rect 23848 36669 23857 36703
rect 23857 36669 23891 36703
rect 23891 36669 23900 36703
rect 23848 36660 23900 36669
rect 24584 36660 24636 36712
rect 25228 36728 25280 36780
rect 27712 36796 27764 36848
rect 28172 36796 28224 36848
rect 30748 36864 30800 36916
rect 32680 36864 32732 36916
rect 33508 36864 33560 36916
rect 25136 36660 25188 36712
rect 25964 36660 26016 36712
rect 26056 36660 26108 36712
rect 27160 36771 27212 36780
rect 27160 36737 27169 36771
rect 27169 36737 27203 36771
rect 27203 36737 27212 36771
rect 27160 36728 27212 36737
rect 29920 36796 29972 36848
rect 31300 36796 31352 36848
rect 35348 36864 35400 36916
rect 36820 36864 36872 36916
rect 38752 36907 38804 36916
rect 38752 36873 38761 36907
rect 38761 36873 38795 36907
rect 38795 36873 38804 36907
rect 38752 36864 38804 36873
rect 36544 36796 36596 36848
rect 49240 36796 49292 36848
rect 15200 36524 15252 36576
rect 15292 36567 15344 36576
rect 15292 36533 15301 36567
rect 15301 36533 15335 36567
rect 15335 36533 15344 36567
rect 15292 36524 15344 36533
rect 16488 36524 16540 36576
rect 26148 36592 26200 36644
rect 27804 36660 27856 36712
rect 30288 36660 30340 36712
rect 30472 36660 30524 36712
rect 32404 36703 32456 36712
rect 32404 36669 32413 36703
rect 32413 36669 32447 36703
rect 32447 36669 32456 36703
rect 32404 36660 32456 36669
rect 32772 36660 32824 36712
rect 33140 36660 33192 36712
rect 34428 36728 34480 36780
rect 36360 36728 36412 36780
rect 47400 36728 47452 36780
rect 49056 36771 49108 36780
rect 49056 36737 49065 36771
rect 49065 36737 49099 36771
rect 49099 36737 49108 36771
rect 49056 36728 49108 36737
rect 34152 36660 34204 36712
rect 38844 36703 38896 36712
rect 38844 36669 38853 36703
rect 38853 36669 38887 36703
rect 38887 36669 38896 36703
rect 38844 36660 38896 36669
rect 48320 36592 48372 36644
rect 19248 36524 19300 36576
rect 21916 36524 21968 36576
rect 22560 36524 22612 36576
rect 22744 36524 22796 36576
rect 30104 36524 30156 36576
rect 32220 36524 32272 36576
rect 34704 36524 34756 36576
rect 35072 36524 35124 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 32950 36422 33002 36474
rect 33014 36422 33066 36474
rect 33078 36422 33130 36474
rect 33142 36422 33194 36474
rect 33206 36422 33258 36474
rect 42950 36422 43002 36474
rect 43014 36422 43066 36474
rect 43078 36422 43130 36474
rect 43142 36422 43194 36474
rect 43206 36422 43258 36474
rect 1768 36320 1820 36372
rect 11796 36320 11848 36372
rect 13452 36320 13504 36372
rect 14648 36320 14700 36372
rect 15476 36320 15528 36372
rect 17408 36320 17460 36372
rect 18512 36320 18564 36372
rect 19340 36320 19392 36372
rect 17224 36252 17276 36304
rect 20720 36252 20772 36304
rect 23756 36320 23808 36372
rect 23848 36320 23900 36372
rect 24676 36320 24728 36372
rect 27712 36320 27764 36372
rect 32312 36320 32364 36372
rect 33508 36320 33560 36372
rect 38568 36320 38620 36372
rect 49240 36363 49292 36372
rect 49240 36329 49249 36363
rect 49249 36329 49283 36363
rect 49283 36329 49292 36363
rect 49240 36320 49292 36329
rect 28816 36252 28868 36304
rect 29184 36295 29236 36304
rect 29184 36261 29193 36295
rect 29193 36261 29227 36295
rect 29227 36261 29236 36295
rect 29184 36252 29236 36261
rect 31852 36252 31904 36304
rect 32864 36252 32916 36304
rect 9588 36184 9640 36236
rect 12440 36184 12492 36236
rect 13452 36227 13504 36236
rect 13452 36193 13461 36227
rect 13461 36193 13495 36227
rect 13495 36193 13504 36227
rect 13452 36184 13504 36193
rect 14372 36184 14424 36236
rect 15108 36227 15160 36236
rect 15108 36193 15117 36227
rect 15117 36193 15151 36227
rect 15151 36193 15160 36227
rect 15108 36184 15160 36193
rect 16120 36227 16172 36236
rect 16120 36193 16129 36227
rect 16129 36193 16163 36227
rect 16163 36193 16172 36227
rect 16120 36184 16172 36193
rect 16856 36227 16908 36236
rect 16856 36193 16865 36227
rect 16865 36193 16899 36227
rect 16899 36193 16908 36227
rect 16856 36184 16908 36193
rect 16948 36227 17000 36236
rect 16948 36193 16957 36227
rect 16957 36193 16991 36227
rect 16991 36193 17000 36227
rect 16948 36184 17000 36193
rect 18880 36184 18932 36236
rect 20444 36184 20496 36236
rect 22008 36184 22060 36236
rect 24584 36227 24636 36236
rect 24584 36193 24593 36227
rect 24593 36193 24627 36227
rect 24627 36193 24636 36227
rect 27436 36227 27488 36236
rect 24584 36184 24636 36193
rect 27436 36193 27445 36227
rect 27445 36193 27479 36227
rect 27479 36193 27488 36227
rect 27436 36184 27488 36193
rect 28356 36184 28408 36236
rect 29920 36184 29972 36236
rect 30288 36184 30340 36236
rect 9496 36159 9548 36168
rect 9496 36125 9505 36159
rect 9505 36125 9539 36159
rect 9539 36125 9548 36159
rect 9496 36116 9548 36125
rect 11980 36159 12032 36168
rect 11980 36125 11989 36159
rect 11989 36125 12023 36159
rect 12023 36125 12032 36159
rect 11980 36116 12032 36125
rect 15016 36116 15068 36168
rect 16764 36116 16816 36168
rect 19064 36116 19116 36168
rect 20812 36116 20864 36168
rect 32312 36116 32364 36168
rect 34888 36116 34940 36168
rect 38660 36184 38712 36236
rect 2780 36091 2832 36100
rect 2780 36057 2789 36091
rect 2789 36057 2823 36091
rect 2823 36057 2832 36091
rect 2780 36048 2832 36057
rect 11060 36048 11112 36100
rect 14648 36048 14700 36100
rect 15476 36048 15528 36100
rect 16304 36048 16356 36100
rect 19156 36048 19208 36100
rect 19708 36091 19760 36100
rect 19708 36057 19717 36091
rect 19717 36057 19751 36091
rect 19751 36057 19760 36091
rect 19708 36048 19760 36057
rect 4804 35980 4856 36032
rect 14188 35980 14240 36032
rect 14556 36023 14608 36032
rect 14556 35989 14565 36023
rect 14565 35989 14599 36023
rect 14599 35989 14608 36023
rect 14556 35980 14608 35989
rect 15108 35980 15160 36032
rect 16396 36023 16448 36032
rect 16396 35989 16405 36023
rect 16405 35989 16439 36023
rect 16439 35989 16448 36023
rect 16396 35980 16448 35989
rect 17040 35980 17092 36032
rect 23848 36048 23900 36100
rect 24492 36048 24544 36100
rect 25136 36048 25188 36100
rect 25504 36048 25556 36100
rect 27712 36048 27764 36100
rect 28172 36048 28224 36100
rect 25872 35980 25924 36032
rect 27896 35980 27948 36032
rect 28540 35980 28592 36032
rect 31300 36048 31352 36100
rect 31024 35980 31076 36032
rect 31208 35980 31260 36032
rect 32680 36091 32732 36100
rect 32680 36057 32689 36091
rect 32689 36057 32723 36091
rect 32723 36057 32732 36091
rect 32680 36048 32732 36057
rect 34152 36091 34204 36100
rect 34152 36057 34161 36091
rect 34161 36057 34195 36091
rect 34195 36057 34204 36091
rect 36360 36116 36412 36168
rect 37096 36116 37148 36168
rect 48320 36116 48372 36168
rect 34152 36048 34204 36057
rect 35348 36048 35400 36100
rect 37372 36048 37424 36100
rect 37464 36048 37516 36100
rect 37096 35980 37148 36032
rect 38844 35980 38896 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 27950 35878 28002 35930
rect 28014 35878 28066 35930
rect 28078 35878 28130 35930
rect 28142 35878 28194 35930
rect 28206 35878 28258 35930
rect 37950 35878 38002 35930
rect 38014 35878 38066 35930
rect 38078 35878 38130 35930
rect 38142 35878 38194 35930
rect 38206 35878 38258 35930
rect 47950 35878 48002 35930
rect 48014 35878 48066 35930
rect 48078 35878 48130 35930
rect 48142 35878 48194 35930
rect 48206 35878 48258 35930
rect 3424 35776 3476 35828
rect 12624 35776 12676 35828
rect 9312 35751 9364 35760
rect 9312 35717 9321 35751
rect 9321 35717 9355 35751
rect 9355 35717 9364 35751
rect 9312 35708 9364 35717
rect 14648 35708 14700 35760
rect 14832 35819 14884 35828
rect 14832 35785 14841 35819
rect 14841 35785 14875 35819
rect 14875 35785 14884 35819
rect 14832 35776 14884 35785
rect 15200 35776 15252 35828
rect 16028 35776 16080 35828
rect 17960 35776 18012 35828
rect 19156 35776 19208 35828
rect 20720 35776 20772 35828
rect 15660 35708 15712 35760
rect 15752 35708 15804 35760
rect 17132 35708 17184 35760
rect 9588 35615 9640 35624
rect 9588 35581 9597 35615
rect 9597 35581 9631 35615
rect 9631 35581 9640 35615
rect 9588 35572 9640 35581
rect 10784 35436 10836 35488
rect 13728 35572 13780 35624
rect 15292 35572 15344 35624
rect 14096 35436 14148 35488
rect 14464 35436 14516 35488
rect 17960 35640 18012 35692
rect 18236 35683 18288 35692
rect 18236 35649 18245 35683
rect 18245 35649 18279 35683
rect 18279 35649 18288 35683
rect 18236 35640 18288 35649
rect 19340 35708 19392 35760
rect 20812 35708 20864 35760
rect 22100 35708 22152 35760
rect 17776 35572 17828 35624
rect 22192 35683 22244 35692
rect 22192 35649 22201 35683
rect 22201 35649 22235 35683
rect 22235 35649 22244 35683
rect 22192 35640 22244 35649
rect 23848 35708 23900 35760
rect 28448 35708 28500 35760
rect 28632 35708 28684 35760
rect 30380 35708 30432 35760
rect 31576 35708 31628 35760
rect 32036 35776 32088 35828
rect 33876 35776 33928 35828
rect 34060 35776 34112 35828
rect 32220 35708 32272 35760
rect 32312 35751 32364 35760
rect 32312 35717 32321 35751
rect 32321 35717 32355 35751
rect 32355 35717 32364 35751
rect 32312 35708 32364 35717
rect 19064 35572 19116 35624
rect 34704 35708 34756 35760
rect 35992 35776 36044 35828
rect 36912 35776 36964 35828
rect 16120 35436 16172 35488
rect 21272 35479 21324 35488
rect 21272 35445 21281 35479
rect 21281 35445 21315 35479
rect 21315 35445 21324 35479
rect 21272 35436 21324 35445
rect 21456 35436 21508 35488
rect 23388 35615 23440 35624
rect 23388 35581 23397 35615
rect 23397 35581 23431 35615
rect 23431 35581 23440 35615
rect 23388 35572 23440 35581
rect 23388 35436 23440 35488
rect 24952 35572 25004 35624
rect 25872 35615 25924 35624
rect 25872 35581 25881 35615
rect 25881 35581 25915 35615
rect 25915 35581 25924 35615
rect 25872 35572 25924 35581
rect 29092 35572 29144 35624
rect 30196 35572 30248 35624
rect 31024 35615 31076 35624
rect 31024 35581 31033 35615
rect 31033 35581 31067 35615
rect 31067 35581 31076 35615
rect 31024 35572 31076 35581
rect 31484 35572 31536 35624
rect 32496 35572 32548 35624
rect 33692 35572 33744 35624
rect 30288 35504 30340 35556
rect 31116 35504 31168 35556
rect 33968 35504 34020 35556
rect 34152 35615 34204 35624
rect 34152 35581 34161 35615
rect 34161 35581 34195 35615
rect 34195 35581 34204 35615
rect 34152 35572 34204 35581
rect 35164 35572 35216 35624
rect 24584 35436 24636 35488
rect 25044 35436 25096 35488
rect 27252 35436 27304 35488
rect 33784 35436 33836 35488
rect 34428 35436 34480 35488
rect 36360 35572 36412 35624
rect 39948 35436 40000 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 32950 35334 33002 35386
rect 33014 35334 33066 35386
rect 33078 35334 33130 35386
rect 33142 35334 33194 35386
rect 33206 35334 33258 35386
rect 42950 35334 43002 35386
rect 43014 35334 43066 35386
rect 43078 35334 43130 35386
rect 43142 35334 43194 35386
rect 43206 35334 43258 35386
rect 1308 35096 1360 35148
rect 12624 35096 12676 35148
rect 13544 35139 13596 35148
rect 13544 35105 13553 35139
rect 13553 35105 13587 35139
rect 13587 35105 13596 35139
rect 13544 35096 13596 35105
rect 10876 35071 10928 35080
rect 10876 35037 10885 35071
rect 10885 35037 10919 35071
rect 10919 35037 10928 35071
rect 10876 35028 10928 35037
rect 18788 35232 18840 35284
rect 21456 35232 21508 35284
rect 22376 35275 22428 35284
rect 22376 35241 22385 35275
rect 22385 35241 22419 35275
rect 22419 35241 22428 35275
rect 22376 35232 22428 35241
rect 23664 35232 23716 35284
rect 24952 35232 25004 35284
rect 29092 35232 29144 35284
rect 30288 35232 30340 35284
rect 31116 35232 31168 35284
rect 15660 35164 15712 35216
rect 16212 35164 16264 35216
rect 14096 35096 14148 35148
rect 15292 35096 15344 35148
rect 16396 35096 16448 35148
rect 15844 35028 15896 35080
rect 17500 35096 17552 35148
rect 18328 35139 18380 35148
rect 18328 35105 18337 35139
rect 18337 35105 18371 35139
rect 18371 35105 18380 35139
rect 18328 35096 18380 35105
rect 19616 35096 19668 35148
rect 20444 35096 20496 35148
rect 21272 35096 21324 35148
rect 22560 35096 22612 35148
rect 23756 35139 23808 35148
rect 23756 35105 23765 35139
rect 23765 35105 23799 35139
rect 23799 35105 23808 35139
rect 23756 35096 23808 35105
rect 24492 35096 24544 35148
rect 24584 35096 24636 35148
rect 29276 35164 29328 35216
rect 31024 35164 31076 35216
rect 17868 35028 17920 35080
rect 20352 35028 20404 35080
rect 27988 35139 28040 35148
rect 27988 35105 27997 35139
rect 27997 35105 28031 35139
rect 28031 35105 28040 35139
rect 27988 35096 28040 35105
rect 14464 34960 14516 35012
rect 14832 34960 14884 35012
rect 16028 34960 16080 35012
rect 20536 34960 20588 35012
rect 20812 34960 20864 35012
rect 10968 34935 11020 34944
rect 10968 34901 10977 34935
rect 10977 34901 11011 34935
rect 11011 34901 11020 34935
rect 10968 34892 11020 34901
rect 12992 34935 13044 34944
rect 12992 34901 13001 34935
rect 13001 34901 13035 34935
rect 13035 34901 13044 34935
rect 12992 34892 13044 34901
rect 13452 34935 13504 34944
rect 13452 34901 13461 34935
rect 13461 34901 13495 34935
rect 13495 34901 13504 34935
rect 13452 34892 13504 34901
rect 17868 34935 17920 34944
rect 17868 34901 17877 34935
rect 17877 34901 17911 34935
rect 17911 34901 17920 34935
rect 17868 34892 17920 34901
rect 18420 34892 18472 34944
rect 19892 34935 19944 34944
rect 19892 34901 19901 34935
rect 19901 34901 19935 34935
rect 19935 34901 19944 34935
rect 19892 34892 19944 34901
rect 20444 34892 20496 34944
rect 22468 34892 22520 34944
rect 25044 34960 25096 35012
rect 25688 34960 25740 35012
rect 29184 35096 29236 35148
rect 30288 35139 30340 35148
rect 30288 35105 30297 35139
rect 30297 35105 30331 35139
rect 30331 35105 30340 35139
rect 30288 35096 30340 35105
rect 32036 35028 32088 35080
rect 32588 35139 32640 35148
rect 32588 35105 32597 35139
rect 32597 35105 32631 35139
rect 32631 35105 32640 35139
rect 32588 35096 32640 35105
rect 37188 35232 37240 35284
rect 34796 35164 34848 35216
rect 32864 35096 32916 35148
rect 35164 35096 35216 35148
rect 33784 35071 33836 35080
rect 33784 35037 33793 35071
rect 33793 35037 33827 35071
rect 33827 35037 33836 35071
rect 33784 35028 33836 35037
rect 34152 35028 34204 35080
rect 34428 35028 34480 35080
rect 36268 35028 36320 35080
rect 39488 35028 39540 35080
rect 49056 35071 49108 35080
rect 49056 35037 49065 35071
rect 49065 35037 49099 35071
rect 49099 35037 49108 35071
rect 49056 35028 49108 35037
rect 30380 34960 30432 35012
rect 33692 34960 33744 35012
rect 34244 34960 34296 35012
rect 25964 34892 26016 34944
rect 29460 34892 29512 34944
rect 31484 34892 31536 34944
rect 32220 34892 32272 34944
rect 34980 34892 35032 34944
rect 37096 34892 37148 34944
rect 42616 34892 42668 34944
rect 48320 34892 48372 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 27950 34790 28002 34842
rect 28014 34790 28066 34842
rect 28078 34790 28130 34842
rect 28142 34790 28194 34842
rect 28206 34790 28258 34842
rect 37950 34790 38002 34842
rect 38014 34790 38066 34842
rect 38078 34790 38130 34842
rect 38142 34790 38194 34842
rect 38206 34790 38258 34842
rect 47950 34790 48002 34842
rect 48014 34790 48066 34842
rect 48078 34790 48130 34842
rect 48142 34790 48194 34842
rect 48206 34790 48258 34842
rect 13452 34688 13504 34740
rect 14556 34688 14608 34740
rect 14740 34731 14792 34740
rect 14740 34697 14749 34731
rect 14749 34697 14783 34731
rect 14783 34697 14792 34731
rect 14740 34688 14792 34697
rect 15384 34688 15436 34740
rect 12992 34620 13044 34672
rect 13912 34620 13964 34672
rect 16212 34620 16264 34672
rect 23204 34688 23256 34740
rect 23664 34688 23716 34740
rect 24032 34688 24084 34740
rect 24400 34688 24452 34740
rect 20720 34620 20772 34672
rect 22376 34620 22428 34672
rect 22928 34620 22980 34672
rect 24676 34663 24728 34672
rect 24676 34629 24685 34663
rect 24685 34629 24719 34663
rect 24719 34629 24728 34663
rect 24676 34620 24728 34629
rect 25596 34688 25648 34740
rect 10968 34552 11020 34604
rect 14372 34552 14424 34604
rect 16304 34552 16356 34604
rect 16672 34552 16724 34604
rect 17500 34552 17552 34604
rect 2044 34527 2096 34536
rect 2044 34493 2053 34527
rect 2053 34493 2087 34527
rect 2087 34493 2096 34527
rect 2044 34484 2096 34493
rect 9588 34484 9640 34536
rect 13636 34527 13688 34536
rect 13636 34493 13645 34527
rect 13645 34493 13679 34527
rect 13679 34493 13688 34527
rect 13636 34484 13688 34493
rect 14832 34484 14884 34536
rect 15844 34484 15896 34536
rect 15568 34459 15620 34468
rect 15568 34425 15577 34459
rect 15577 34425 15611 34459
rect 15611 34425 15620 34459
rect 15568 34416 15620 34425
rect 16396 34484 16448 34536
rect 13360 34348 13412 34400
rect 14556 34348 14608 34400
rect 18236 34595 18288 34604
rect 18236 34561 18245 34595
rect 18245 34561 18279 34595
rect 18279 34561 18288 34595
rect 18236 34552 18288 34561
rect 19064 34595 19116 34604
rect 19064 34561 19073 34595
rect 19073 34561 19107 34595
rect 19107 34561 19116 34595
rect 19064 34552 19116 34561
rect 25688 34552 25740 34604
rect 27712 34688 27764 34740
rect 27804 34688 27856 34740
rect 30380 34688 30432 34740
rect 27436 34620 27488 34672
rect 27896 34620 27948 34672
rect 27160 34595 27212 34604
rect 27160 34561 27169 34595
rect 27169 34561 27203 34595
rect 27203 34561 27212 34595
rect 27160 34552 27212 34561
rect 19340 34484 19392 34536
rect 19708 34484 19760 34536
rect 20628 34484 20680 34536
rect 22008 34527 22060 34536
rect 22008 34493 22017 34527
rect 22017 34493 22051 34527
rect 22051 34493 22060 34527
rect 22008 34484 22060 34493
rect 26332 34484 26384 34536
rect 31208 34620 31260 34672
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 29920 34552 29972 34561
rect 32864 34688 32916 34740
rect 36636 34688 36688 34740
rect 37556 34688 37608 34740
rect 44180 34688 44232 34740
rect 47400 34688 47452 34740
rect 32128 34552 32180 34604
rect 28816 34484 28868 34536
rect 18880 34348 18932 34400
rect 19524 34348 19576 34400
rect 21640 34348 21692 34400
rect 22100 34348 22152 34400
rect 22928 34348 22980 34400
rect 23848 34348 23900 34400
rect 24400 34348 24452 34400
rect 29368 34348 29420 34400
rect 29828 34348 29880 34400
rect 31668 34527 31720 34536
rect 31668 34493 31677 34527
rect 31677 34493 31711 34527
rect 31711 34493 31720 34527
rect 31668 34484 31720 34493
rect 31576 34416 31628 34468
rect 32220 34484 32272 34536
rect 34060 34620 34112 34672
rect 36268 34620 36320 34672
rect 34336 34552 34388 34604
rect 38568 34552 38620 34604
rect 41328 34595 41380 34604
rect 41328 34561 41337 34595
rect 41337 34561 41371 34595
rect 41371 34561 41380 34595
rect 41328 34552 41380 34561
rect 49332 34595 49384 34604
rect 49332 34561 49341 34595
rect 49341 34561 49375 34595
rect 49375 34561 49384 34595
rect 49332 34552 49384 34561
rect 32772 34484 32824 34536
rect 33508 34484 33560 34536
rect 34428 34484 34480 34536
rect 35808 34484 35860 34536
rect 32588 34416 32640 34468
rect 33692 34391 33744 34400
rect 33692 34357 33701 34391
rect 33701 34357 33735 34391
rect 33735 34357 33744 34391
rect 33692 34348 33744 34357
rect 35992 34348 36044 34400
rect 36268 34391 36320 34400
rect 36268 34357 36277 34391
rect 36277 34357 36311 34391
rect 36311 34357 36320 34391
rect 36268 34348 36320 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 32950 34246 33002 34298
rect 33014 34246 33066 34298
rect 33078 34246 33130 34298
rect 33142 34246 33194 34298
rect 33206 34246 33258 34298
rect 42950 34246 43002 34298
rect 43014 34246 43066 34298
rect 43078 34246 43130 34298
rect 43142 34246 43194 34298
rect 43206 34246 43258 34298
rect 14280 34187 14332 34196
rect 14280 34153 14289 34187
rect 14289 34153 14323 34187
rect 14323 34153 14332 34187
rect 14280 34144 14332 34153
rect 10784 34008 10836 34060
rect 12532 34008 12584 34060
rect 11796 33983 11848 33992
rect 11796 33949 11805 33983
rect 11805 33949 11839 33983
rect 11839 33949 11848 33983
rect 11796 33940 11848 33949
rect 15292 34008 15344 34060
rect 17132 34144 17184 34196
rect 19064 34144 19116 34196
rect 19248 34144 19300 34196
rect 21456 34144 21508 34196
rect 21640 34144 21692 34196
rect 23572 34144 23624 34196
rect 25964 34187 26016 34196
rect 25964 34153 25973 34187
rect 25973 34153 26007 34187
rect 26007 34153 26016 34187
rect 25964 34144 26016 34153
rect 28908 34144 28960 34196
rect 17684 34076 17736 34128
rect 17592 34008 17644 34060
rect 24124 34076 24176 34128
rect 34336 34144 34388 34196
rect 18788 33940 18840 33992
rect 25872 34008 25924 34060
rect 30012 34008 30064 34060
rect 34612 34076 34664 34128
rect 34704 34076 34756 34128
rect 31116 34008 31168 34060
rect 32404 34008 32456 34060
rect 33324 34008 33376 34060
rect 34336 34008 34388 34060
rect 22008 33940 22060 33992
rect 25228 33940 25280 33992
rect 27620 33983 27672 33992
rect 27620 33949 27629 33983
rect 27629 33949 27663 33983
rect 27663 33949 27672 33983
rect 27620 33940 27672 33949
rect 27712 33940 27764 33992
rect 28816 33940 28868 33992
rect 14464 33804 14516 33856
rect 15384 33804 15436 33856
rect 16028 33872 16080 33924
rect 16580 33804 16632 33856
rect 20168 33872 20220 33924
rect 20720 33872 20772 33924
rect 18788 33804 18840 33856
rect 29552 33872 29604 33924
rect 32496 33940 32548 33992
rect 34152 33940 34204 33992
rect 36084 33940 36136 33992
rect 30104 33804 30156 33856
rect 30840 33804 30892 33856
rect 31024 33804 31076 33856
rect 32404 33872 32456 33924
rect 33140 33872 33192 33924
rect 33048 33804 33100 33856
rect 33232 33804 33284 33856
rect 35532 33804 35584 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 27950 33702 28002 33754
rect 28014 33702 28066 33754
rect 28078 33702 28130 33754
rect 28142 33702 28194 33754
rect 28206 33702 28258 33754
rect 37950 33702 38002 33754
rect 38014 33702 38066 33754
rect 38078 33702 38130 33754
rect 38142 33702 38194 33754
rect 38206 33702 38258 33754
rect 47950 33702 48002 33754
rect 48014 33702 48066 33754
rect 48078 33702 48130 33754
rect 48142 33702 48194 33754
rect 48206 33702 48258 33754
rect 14372 33643 14424 33652
rect 14372 33609 14381 33643
rect 14381 33609 14415 33643
rect 14415 33609 14424 33643
rect 14372 33600 14424 33609
rect 16396 33600 16448 33652
rect 17868 33600 17920 33652
rect 20536 33600 20588 33652
rect 21088 33643 21140 33652
rect 21088 33609 21097 33643
rect 21097 33609 21131 33643
rect 21131 33609 21140 33643
rect 21088 33600 21140 33609
rect 22100 33600 22152 33652
rect 14188 33532 14240 33584
rect 17684 33532 17736 33584
rect 8576 33464 8628 33516
rect 13544 33464 13596 33516
rect 1308 33396 1360 33448
rect 14648 33396 14700 33448
rect 16488 33464 16540 33516
rect 18420 33464 18472 33516
rect 18604 33575 18656 33584
rect 18604 33541 18613 33575
rect 18613 33541 18647 33575
rect 18647 33541 18656 33575
rect 18604 33532 18656 33541
rect 18788 33532 18840 33584
rect 19064 33532 19116 33584
rect 19248 33532 19300 33584
rect 21272 33532 21324 33584
rect 21364 33532 21416 33584
rect 22284 33532 22336 33584
rect 23940 33600 23992 33652
rect 20996 33464 21048 33516
rect 24584 33532 24636 33584
rect 24676 33532 24728 33584
rect 31116 33600 31168 33652
rect 31208 33600 31260 33652
rect 33140 33600 33192 33652
rect 27896 33532 27948 33584
rect 30748 33532 30800 33584
rect 33692 33600 33744 33652
rect 36268 33600 36320 33652
rect 33784 33532 33836 33584
rect 27160 33507 27212 33516
rect 27160 33473 27169 33507
rect 27169 33473 27203 33507
rect 27203 33473 27212 33507
rect 27160 33464 27212 33473
rect 29552 33507 29604 33516
rect 29552 33473 29561 33507
rect 29561 33473 29595 33507
rect 29595 33473 29604 33507
rect 29552 33464 29604 33473
rect 29736 33464 29788 33516
rect 30012 33507 30064 33516
rect 30012 33473 30021 33507
rect 30021 33473 30055 33507
rect 30055 33473 30064 33507
rect 30012 33464 30064 33473
rect 32404 33464 32456 33516
rect 39672 33507 39724 33516
rect 39672 33473 39681 33507
rect 39681 33473 39715 33507
rect 39715 33473 39724 33507
rect 39672 33464 39724 33473
rect 39856 33464 39908 33516
rect 49148 33507 49200 33516
rect 49148 33473 49157 33507
rect 49157 33473 49191 33507
rect 49191 33473 49200 33507
rect 49148 33464 49200 33473
rect 17684 33396 17736 33448
rect 17776 33396 17828 33448
rect 18788 33396 18840 33448
rect 19248 33328 19300 33380
rect 17408 33303 17460 33312
rect 17408 33269 17417 33303
rect 17417 33269 17451 33303
rect 17451 33269 17460 33303
rect 17408 33260 17460 33269
rect 17868 33260 17920 33312
rect 21364 33396 21416 33448
rect 22008 33439 22060 33448
rect 22008 33405 22017 33439
rect 22017 33405 22051 33439
rect 22051 33405 22060 33439
rect 22008 33396 22060 33405
rect 22284 33439 22336 33448
rect 22284 33405 22293 33439
rect 22293 33405 22327 33439
rect 22327 33405 22336 33439
rect 22284 33396 22336 33405
rect 24032 33396 24084 33448
rect 25228 33396 25280 33448
rect 25596 33396 25648 33448
rect 31668 33396 31720 33448
rect 32588 33396 32640 33448
rect 33692 33396 33744 33448
rect 34060 33396 34112 33448
rect 34336 33328 34388 33380
rect 44088 33328 44140 33380
rect 21456 33260 21508 33312
rect 21640 33260 21692 33312
rect 27252 33260 27304 33312
rect 30472 33260 30524 33312
rect 30748 33260 30800 33312
rect 30840 33260 30892 33312
rect 33048 33260 33100 33312
rect 36176 33260 36228 33312
rect 45836 33260 45888 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 32950 33158 33002 33210
rect 33014 33158 33066 33210
rect 33078 33158 33130 33210
rect 33142 33158 33194 33210
rect 33206 33158 33258 33210
rect 42950 33158 43002 33210
rect 43014 33158 43066 33210
rect 43078 33158 43130 33210
rect 43142 33158 43194 33210
rect 43206 33158 43258 33210
rect 1308 32920 1360 32972
rect 16672 33056 16724 33108
rect 18420 33056 18472 33108
rect 18696 33056 18748 33108
rect 18972 33056 19024 33108
rect 15292 32920 15344 32972
rect 16212 32920 16264 32972
rect 20076 32988 20128 33040
rect 22928 33056 22980 33108
rect 24860 33056 24912 33108
rect 31576 33056 31628 33108
rect 23572 32988 23624 33040
rect 31300 32988 31352 33040
rect 20628 32920 20680 32972
rect 23664 32920 23716 32972
rect 27252 32920 27304 32972
rect 13544 32852 13596 32904
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 21364 32895 21416 32904
rect 21364 32861 21373 32895
rect 21373 32861 21407 32895
rect 21407 32861 21416 32895
rect 21364 32852 21416 32861
rect 15936 32784 15988 32836
rect 20076 32784 20128 32836
rect 20720 32784 20772 32836
rect 22100 32784 22152 32836
rect 23572 32784 23624 32836
rect 25412 32852 25464 32904
rect 27620 32852 27672 32904
rect 25320 32784 25372 32836
rect 28356 32920 28408 32972
rect 28632 32920 28684 32972
rect 30104 32920 30156 32972
rect 30472 32920 30524 32972
rect 31208 32920 31260 32972
rect 32588 32963 32640 32972
rect 32588 32929 32597 32963
rect 32597 32929 32631 32963
rect 32631 32929 32640 32963
rect 32588 32920 32640 32929
rect 33508 32920 33560 32972
rect 29184 32895 29236 32904
rect 29184 32861 29193 32895
rect 29193 32861 29227 32895
rect 29227 32861 29236 32895
rect 29184 32852 29236 32861
rect 29736 32895 29788 32904
rect 29736 32861 29745 32895
rect 29745 32861 29779 32895
rect 29779 32861 29788 32895
rect 29736 32852 29788 32861
rect 49056 32895 49108 32904
rect 49056 32861 49065 32895
rect 49065 32861 49099 32895
rect 49099 32861 49108 32895
rect 49056 32852 49108 32861
rect 30288 32784 30340 32836
rect 30472 32784 30524 32836
rect 31852 32784 31904 32836
rect 16396 32716 16448 32768
rect 17132 32716 17184 32768
rect 17500 32716 17552 32768
rect 19340 32716 19392 32768
rect 20444 32716 20496 32768
rect 20628 32759 20680 32768
rect 20628 32725 20637 32759
rect 20637 32725 20671 32759
rect 20671 32725 20680 32759
rect 20628 32716 20680 32725
rect 23848 32716 23900 32768
rect 27620 32716 27672 32768
rect 28540 32716 28592 32768
rect 32128 32716 32180 32768
rect 33140 32784 33192 32836
rect 33876 32784 33928 32836
rect 36728 32716 36780 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 27950 32614 28002 32666
rect 28014 32614 28066 32666
rect 28078 32614 28130 32666
rect 28142 32614 28194 32666
rect 28206 32614 28258 32666
rect 37950 32614 38002 32666
rect 38014 32614 38066 32666
rect 38078 32614 38130 32666
rect 38142 32614 38194 32666
rect 38206 32614 38258 32666
rect 47950 32614 48002 32666
rect 48014 32614 48066 32666
rect 48078 32614 48130 32666
rect 48142 32614 48194 32666
rect 48206 32614 48258 32666
rect 12808 32512 12860 32564
rect 1860 32172 1912 32224
rect 16212 32512 16264 32564
rect 14556 32487 14608 32496
rect 14556 32453 14565 32487
rect 14565 32453 14599 32487
rect 14599 32453 14608 32487
rect 14556 32444 14608 32453
rect 16028 32444 16080 32496
rect 16396 32444 16448 32496
rect 13728 32308 13780 32360
rect 15292 32308 15344 32360
rect 20260 32512 20312 32564
rect 20996 32555 21048 32564
rect 20996 32521 21005 32555
rect 21005 32521 21039 32555
rect 21039 32521 21048 32555
rect 20996 32512 21048 32521
rect 21732 32512 21784 32564
rect 22836 32512 22888 32564
rect 17684 32444 17736 32496
rect 19800 32444 19852 32496
rect 20076 32444 20128 32496
rect 22284 32444 22336 32496
rect 17316 32376 17368 32428
rect 19064 32376 19116 32428
rect 22192 32376 22244 32428
rect 17500 32351 17552 32360
rect 17500 32317 17509 32351
rect 17509 32317 17543 32351
rect 17543 32317 17552 32351
rect 17500 32308 17552 32317
rect 17684 32351 17736 32360
rect 17684 32317 17693 32351
rect 17693 32317 17727 32351
rect 17727 32317 17736 32351
rect 17684 32308 17736 32317
rect 18052 32308 18104 32360
rect 22560 32351 22612 32360
rect 22560 32317 22569 32351
rect 22569 32317 22603 32351
rect 22603 32317 22612 32351
rect 22560 32308 22612 32317
rect 22836 32376 22888 32428
rect 23848 32444 23900 32496
rect 23940 32487 23992 32496
rect 23940 32453 23949 32487
rect 23949 32453 23983 32487
rect 23983 32453 23992 32487
rect 23940 32444 23992 32453
rect 24400 32444 24452 32496
rect 28540 32487 28592 32496
rect 28540 32453 28549 32487
rect 28549 32453 28583 32487
rect 28583 32453 28592 32487
rect 28540 32444 28592 32453
rect 30564 32512 30616 32564
rect 33600 32512 33652 32564
rect 35440 32512 35492 32564
rect 31300 32444 31352 32496
rect 31668 32444 31720 32496
rect 30472 32376 30524 32428
rect 30840 32419 30892 32428
rect 30840 32385 30849 32419
rect 30849 32385 30883 32419
rect 30883 32385 30892 32419
rect 30840 32376 30892 32385
rect 32680 32419 32732 32428
rect 32680 32385 32689 32419
rect 32689 32385 32723 32419
rect 32723 32385 32732 32419
rect 32680 32376 32732 32385
rect 32864 32376 32916 32428
rect 12716 32215 12768 32224
rect 12716 32181 12725 32215
rect 12725 32181 12759 32215
rect 12759 32181 12768 32215
rect 12716 32172 12768 32181
rect 17316 32240 17368 32292
rect 19064 32240 19116 32292
rect 22284 32240 22336 32292
rect 16028 32215 16080 32224
rect 16028 32181 16037 32215
rect 16037 32181 16071 32215
rect 16071 32181 16080 32215
rect 16028 32172 16080 32181
rect 19708 32172 19760 32224
rect 20720 32172 20772 32224
rect 21548 32172 21600 32224
rect 29092 32308 29144 32360
rect 29276 32308 29328 32360
rect 30380 32308 30432 32360
rect 32772 32351 32824 32360
rect 32772 32317 32781 32351
rect 32781 32317 32815 32351
rect 32815 32317 32824 32351
rect 32772 32308 32824 32317
rect 33324 32376 33376 32428
rect 33784 32376 33836 32428
rect 33876 32419 33928 32428
rect 33876 32385 33885 32419
rect 33885 32385 33919 32419
rect 33919 32385 33928 32419
rect 33876 32376 33928 32385
rect 36544 32419 36596 32428
rect 36544 32385 36553 32419
rect 36553 32385 36587 32419
rect 36587 32385 36596 32419
rect 36544 32376 36596 32385
rect 32036 32240 32088 32292
rect 23940 32172 23992 32224
rect 28540 32172 28592 32224
rect 28724 32172 28776 32224
rect 30104 32172 30156 32224
rect 31944 32172 31996 32224
rect 36728 32351 36780 32360
rect 36728 32317 36737 32351
rect 36737 32317 36771 32351
rect 36771 32317 36780 32351
rect 36728 32308 36780 32317
rect 37832 32240 37884 32292
rect 34244 32172 34296 32224
rect 34612 32172 34664 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 32950 32070 33002 32122
rect 33014 32070 33066 32122
rect 33078 32070 33130 32122
rect 33142 32070 33194 32122
rect 33206 32070 33258 32122
rect 42950 32070 43002 32122
rect 43014 32070 43066 32122
rect 43078 32070 43130 32122
rect 43142 32070 43194 32122
rect 43206 32070 43258 32122
rect 1308 31832 1360 31884
rect 12716 31900 12768 31952
rect 7380 31764 7432 31816
rect 13636 31832 13688 31884
rect 16580 32011 16632 32020
rect 16580 31977 16589 32011
rect 16589 31977 16623 32011
rect 16623 31977 16632 32011
rect 16580 31968 16632 31977
rect 17316 31968 17368 32020
rect 17500 31968 17552 32020
rect 18052 31968 18104 32020
rect 18788 32011 18840 32020
rect 18788 31977 18797 32011
rect 18797 31977 18831 32011
rect 18831 31977 18840 32011
rect 18788 31968 18840 31977
rect 19432 31968 19484 32020
rect 22652 31968 22704 32020
rect 23664 31968 23716 32020
rect 24032 32011 24084 32020
rect 24032 31977 24041 32011
rect 24041 31977 24075 32011
rect 24075 31977 24084 32011
rect 24032 31968 24084 31977
rect 30104 31968 30156 32020
rect 19064 31900 19116 31952
rect 20720 31900 20772 31952
rect 15200 31832 15252 31884
rect 19248 31832 19300 31884
rect 21456 31900 21508 31952
rect 21364 31832 21416 31884
rect 21640 31875 21692 31884
rect 21640 31841 21649 31875
rect 21649 31841 21683 31875
rect 21683 31841 21692 31875
rect 21640 31832 21692 31841
rect 22284 31875 22336 31884
rect 19616 31764 19668 31816
rect 11060 31671 11112 31680
rect 11060 31637 11069 31671
rect 11069 31637 11103 31671
rect 11103 31637 11112 31671
rect 11060 31628 11112 31637
rect 16396 31696 16448 31748
rect 16856 31696 16908 31748
rect 19064 31696 19116 31748
rect 20076 31696 20128 31748
rect 20168 31739 20220 31748
rect 20168 31705 20177 31739
rect 20177 31705 20211 31739
rect 20211 31705 20220 31739
rect 20168 31696 20220 31705
rect 20812 31764 20864 31816
rect 22284 31841 22293 31875
rect 22293 31841 22327 31875
rect 22327 31841 22336 31875
rect 22284 31832 22336 31841
rect 23940 31832 23992 31884
rect 26332 31875 26384 31884
rect 26332 31841 26341 31875
rect 26341 31841 26375 31875
rect 26375 31841 26384 31875
rect 26332 31832 26384 31841
rect 26976 31832 27028 31884
rect 27804 31807 27856 31816
rect 27804 31773 27813 31807
rect 27813 31773 27847 31807
rect 27847 31773 27856 31807
rect 27804 31764 27856 31773
rect 21088 31696 21140 31748
rect 22008 31696 22060 31748
rect 28724 31875 28776 31884
rect 28724 31841 28733 31875
rect 28733 31841 28767 31875
rect 28767 31841 28776 31875
rect 28724 31832 28776 31841
rect 29460 31900 29512 31952
rect 28908 31875 28960 31884
rect 28908 31841 28917 31875
rect 28917 31841 28951 31875
rect 28951 31841 28960 31875
rect 28908 31832 28960 31841
rect 29092 31832 29144 31884
rect 29736 31875 29788 31884
rect 29736 31841 29745 31875
rect 29745 31841 29779 31875
rect 29779 31841 29788 31875
rect 29736 31832 29788 31841
rect 30012 31832 30064 31884
rect 31852 31968 31904 32020
rect 31116 31900 31168 31952
rect 32128 31900 32180 31952
rect 33416 31968 33468 32020
rect 33784 31968 33836 32020
rect 29000 31764 29052 31816
rect 31208 31832 31260 31884
rect 31392 31832 31444 31884
rect 31300 31764 31352 31816
rect 33692 31875 33744 31884
rect 33692 31841 33701 31875
rect 33701 31841 33735 31875
rect 33735 31841 33744 31875
rect 33692 31832 33744 31841
rect 33600 31807 33652 31816
rect 33600 31773 33609 31807
rect 33609 31773 33643 31807
rect 33643 31773 33652 31807
rect 33600 31764 33652 31773
rect 49056 31807 49108 31816
rect 49056 31773 49065 31807
rect 49065 31773 49099 31807
rect 49099 31773 49108 31807
rect 49056 31764 49108 31773
rect 30012 31739 30064 31748
rect 30012 31705 30021 31739
rect 30021 31705 30055 31739
rect 30055 31705 30064 31739
rect 30012 31696 30064 31705
rect 33508 31739 33560 31748
rect 33508 31705 33517 31739
rect 33517 31705 33551 31739
rect 33551 31705 33560 31739
rect 33508 31696 33560 31705
rect 16488 31628 16540 31680
rect 19524 31628 19576 31680
rect 19800 31671 19852 31680
rect 19800 31637 19809 31671
rect 19809 31637 19843 31671
rect 19843 31637 19852 31671
rect 19800 31628 19852 31637
rect 21364 31628 21416 31680
rect 21640 31628 21692 31680
rect 22192 31628 22244 31680
rect 28724 31628 28776 31680
rect 32312 31671 32364 31680
rect 32312 31637 32321 31671
rect 32321 31637 32355 31671
rect 32355 31637 32364 31671
rect 32312 31628 32364 31637
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 27950 31526 28002 31578
rect 28014 31526 28066 31578
rect 28078 31526 28130 31578
rect 28142 31526 28194 31578
rect 28206 31526 28258 31578
rect 37950 31526 38002 31578
rect 38014 31526 38066 31578
rect 38078 31526 38130 31578
rect 38142 31526 38194 31578
rect 38206 31526 38258 31578
rect 47950 31526 48002 31578
rect 48014 31526 48066 31578
rect 48078 31526 48130 31578
rect 48142 31526 48194 31578
rect 48206 31526 48258 31578
rect 11060 31356 11112 31408
rect 13544 31467 13596 31476
rect 13544 31433 13553 31467
rect 13553 31433 13587 31467
rect 13587 31433 13596 31467
rect 13544 31424 13596 31433
rect 13636 31467 13688 31476
rect 13636 31433 13645 31467
rect 13645 31433 13679 31467
rect 13679 31433 13688 31467
rect 13636 31424 13688 31433
rect 14740 31467 14792 31476
rect 14740 31433 14749 31467
rect 14749 31433 14783 31467
rect 14783 31433 14792 31467
rect 14740 31424 14792 31433
rect 15660 31424 15712 31476
rect 17224 31424 17276 31476
rect 17408 31467 17460 31476
rect 17408 31433 17417 31467
rect 17417 31433 17451 31467
rect 17451 31433 17460 31467
rect 17408 31424 17460 31433
rect 15752 31356 15804 31408
rect 16120 31356 16172 31408
rect 10692 31331 10744 31340
rect 10692 31297 10701 31331
rect 10701 31297 10735 31331
rect 10735 31297 10744 31331
rect 10692 31288 10744 31297
rect 1308 31220 1360 31272
rect 12532 31220 12584 31272
rect 13728 31263 13780 31272
rect 13728 31229 13737 31263
rect 13737 31229 13771 31263
rect 13771 31229 13780 31263
rect 13728 31220 13780 31229
rect 14740 31220 14792 31272
rect 15476 31288 15528 31340
rect 20812 31424 20864 31476
rect 27804 31424 27856 31476
rect 29184 31424 29236 31476
rect 19064 31356 19116 31408
rect 20904 31356 20956 31408
rect 21640 31356 21692 31408
rect 31484 31356 31536 31408
rect 21272 31288 21324 31340
rect 33600 31356 33652 31408
rect 39948 31356 40000 31408
rect 32680 31288 32732 31340
rect 37188 31288 37240 31340
rect 49332 31331 49384 31340
rect 49332 31297 49341 31331
rect 49341 31297 49375 31331
rect 49375 31297 49384 31331
rect 49332 31288 49384 31297
rect 15844 31220 15896 31272
rect 16028 31152 16080 31204
rect 16212 31263 16264 31272
rect 16212 31229 16221 31263
rect 16221 31229 16255 31263
rect 16255 31229 16264 31263
rect 16212 31220 16264 31229
rect 17408 31220 17460 31272
rect 17868 31152 17920 31204
rect 19524 31152 19576 31204
rect 20904 31263 20956 31272
rect 20904 31229 20913 31263
rect 20913 31229 20947 31263
rect 20947 31229 20956 31263
rect 20904 31220 20956 31229
rect 21088 31263 21140 31272
rect 21088 31229 21097 31263
rect 21097 31229 21131 31263
rect 21131 31229 21140 31263
rect 21088 31220 21140 31229
rect 21916 31220 21968 31272
rect 22560 31220 22612 31272
rect 26516 31220 26568 31272
rect 27620 31220 27672 31272
rect 29276 31220 29328 31272
rect 29828 31263 29880 31272
rect 29828 31229 29837 31263
rect 29837 31229 29871 31263
rect 29871 31229 29880 31263
rect 29828 31220 29880 31229
rect 38568 31220 38620 31272
rect 22376 31152 22428 31204
rect 8668 31084 8720 31136
rect 14832 31084 14884 31136
rect 15936 31084 15988 31136
rect 16212 31084 16264 31136
rect 18512 31084 18564 31136
rect 20444 31127 20496 31136
rect 20444 31093 20453 31127
rect 20453 31093 20487 31127
rect 20487 31093 20496 31127
rect 20444 31084 20496 31093
rect 20904 31084 20956 31136
rect 21732 31084 21784 31136
rect 25136 31152 25188 31204
rect 30840 31152 30892 31204
rect 46756 31152 46808 31204
rect 23388 31127 23440 31136
rect 23388 31093 23397 31127
rect 23397 31093 23431 31127
rect 23431 31093 23440 31127
rect 23388 31084 23440 31093
rect 24952 31084 25004 31136
rect 33876 31084 33928 31136
rect 44548 31084 44600 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 32950 30982 33002 31034
rect 33014 30982 33066 31034
rect 33078 30982 33130 31034
rect 33142 30982 33194 31034
rect 33206 30982 33258 31034
rect 42950 30982 43002 31034
rect 43014 30982 43066 31034
rect 43078 30982 43130 31034
rect 43142 30982 43194 31034
rect 43206 30982 43258 31034
rect 10692 30880 10744 30932
rect 14464 30744 14516 30796
rect 15016 30787 15068 30796
rect 15016 30753 15025 30787
rect 15025 30753 15059 30787
rect 15059 30753 15068 30787
rect 15016 30744 15068 30753
rect 16672 30744 16724 30796
rect 16856 30744 16908 30796
rect 19064 30812 19116 30864
rect 19340 30812 19392 30864
rect 11152 30676 11204 30728
rect 14832 30719 14884 30728
rect 14832 30685 14841 30719
rect 14841 30685 14875 30719
rect 14875 30685 14884 30719
rect 14832 30676 14884 30685
rect 15200 30676 15252 30728
rect 17868 30787 17920 30796
rect 17868 30753 17877 30787
rect 17877 30753 17911 30787
rect 17911 30753 17920 30787
rect 17868 30744 17920 30753
rect 22560 30880 22612 30932
rect 23296 30880 23348 30932
rect 30196 30880 30248 30932
rect 20168 30812 20220 30864
rect 12808 30651 12860 30660
rect 12808 30617 12817 30651
rect 12817 30617 12851 30651
rect 12851 30617 12860 30651
rect 12808 30608 12860 30617
rect 11060 30540 11112 30592
rect 15844 30540 15896 30592
rect 16396 30608 16448 30660
rect 20720 30744 20772 30796
rect 18788 30676 18840 30728
rect 23572 30744 23624 30796
rect 23940 30787 23992 30796
rect 23940 30753 23949 30787
rect 23949 30753 23983 30787
rect 23983 30753 23992 30787
rect 23940 30744 23992 30753
rect 24952 30719 25004 30728
rect 24952 30685 24961 30719
rect 24961 30685 24995 30719
rect 24995 30685 25004 30719
rect 24952 30676 25004 30685
rect 25228 30787 25280 30796
rect 25228 30753 25237 30787
rect 25237 30753 25271 30787
rect 25271 30753 25280 30787
rect 25228 30744 25280 30753
rect 26884 30744 26936 30796
rect 42616 30676 42668 30728
rect 22192 30608 22244 30660
rect 28724 30608 28776 30660
rect 46480 30608 46532 30660
rect 18972 30540 19024 30592
rect 21180 30540 21232 30592
rect 23664 30583 23716 30592
rect 23664 30549 23673 30583
rect 23673 30549 23707 30583
rect 23707 30549 23716 30583
rect 23664 30540 23716 30549
rect 26700 30540 26752 30592
rect 27712 30540 27764 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 27950 30438 28002 30490
rect 28014 30438 28066 30490
rect 28078 30438 28130 30490
rect 28142 30438 28194 30490
rect 28206 30438 28258 30490
rect 37950 30438 38002 30490
rect 38014 30438 38066 30490
rect 38078 30438 38130 30490
rect 38142 30438 38194 30490
rect 38206 30438 38258 30490
rect 47950 30438 48002 30490
rect 48014 30438 48066 30490
rect 48078 30438 48130 30490
rect 48142 30438 48194 30490
rect 48206 30438 48258 30490
rect 12808 30336 12860 30388
rect 16672 30268 16724 30320
rect 7380 30200 7432 30252
rect 18604 30200 18656 30252
rect 19524 30200 19576 30252
rect 19892 30268 19944 30320
rect 20628 30268 20680 30320
rect 22192 30243 22244 30252
rect 22192 30209 22201 30243
rect 22201 30209 22235 30243
rect 22235 30209 22244 30243
rect 22192 30200 22244 30209
rect 22744 30336 22796 30388
rect 23388 30336 23440 30388
rect 23664 30336 23716 30388
rect 31024 30336 31076 30388
rect 33600 30336 33652 30388
rect 40132 30336 40184 30388
rect 23572 30268 23624 30320
rect 30012 30200 30064 30252
rect 37372 30200 37424 30252
rect 49056 30243 49108 30252
rect 49056 30209 49065 30243
rect 49065 30209 49099 30243
rect 49099 30209 49108 30243
rect 49056 30200 49108 30209
rect 1308 30132 1360 30184
rect 14096 30175 14148 30184
rect 14096 30141 14105 30175
rect 14105 30141 14139 30175
rect 14139 30141 14148 30175
rect 14096 30132 14148 30141
rect 13728 30064 13780 30116
rect 16212 30132 16264 30184
rect 17132 30132 17184 30184
rect 20352 30132 20404 30184
rect 20996 30132 21048 30184
rect 21456 30175 21508 30184
rect 21456 30141 21465 30175
rect 21465 30141 21499 30175
rect 21499 30141 21508 30175
rect 21456 30132 21508 30141
rect 15936 29996 15988 30048
rect 16304 29996 16356 30048
rect 22008 29996 22060 30048
rect 22284 29996 22336 30048
rect 29092 29996 29144 30048
rect 39396 29996 39448 30048
rect 49240 30039 49292 30048
rect 49240 30005 49249 30039
rect 49249 30005 49283 30039
rect 49283 30005 49292 30039
rect 49240 29996 49292 30005
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 32950 29894 33002 29946
rect 33014 29894 33066 29946
rect 33078 29894 33130 29946
rect 33142 29894 33194 29946
rect 33206 29894 33258 29946
rect 42950 29894 43002 29946
rect 43014 29894 43066 29946
rect 43078 29894 43130 29946
rect 43142 29894 43194 29946
rect 43206 29894 43258 29946
rect 19524 29792 19576 29844
rect 27528 29792 27580 29844
rect 49240 29792 49292 29844
rect 1308 29656 1360 29708
rect 8668 29588 8720 29640
rect 14096 29588 14148 29640
rect 15016 29656 15068 29708
rect 17132 29656 17184 29708
rect 18880 29699 18932 29708
rect 18880 29665 18889 29699
rect 18889 29665 18923 29699
rect 18923 29665 18932 29699
rect 18880 29656 18932 29665
rect 21456 29656 21508 29708
rect 21916 29699 21968 29708
rect 21916 29665 21925 29699
rect 21925 29665 21959 29699
rect 21959 29665 21968 29699
rect 21916 29656 21968 29665
rect 16856 29631 16908 29640
rect 16856 29597 16865 29631
rect 16865 29597 16899 29631
rect 16899 29597 16908 29631
rect 16856 29588 16908 29597
rect 19892 29631 19944 29640
rect 19892 29597 19901 29631
rect 19901 29597 19935 29631
rect 19935 29597 19944 29631
rect 19892 29588 19944 29597
rect 14924 29563 14976 29572
rect 14924 29529 14933 29563
rect 14933 29529 14967 29563
rect 14967 29529 14976 29563
rect 14924 29520 14976 29529
rect 16672 29520 16724 29572
rect 15936 29452 15988 29504
rect 16396 29495 16448 29504
rect 16396 29461 16405 29495
rect 16405 29461 16439 29495
rect 16439 29461 16448 29495
rect 16396 29452 16448 29461
rect 19064 29520 19116 29572
rect 20628 29520 20680 29572
rect 28632 29656 28684 29708
rect 22376 29588 22428 29640
rect 30012 29588 30064 29640
rect 18788 29452 18840 29504
rect 20536 29452 20588 29504
rect 25872 29563 25924 29572
rect 25872 29529 25881 29563
rect 25881 29529 25915 29563
rect 25915 29529 25924 29563
rect 25872 29520 25924 29529
rect 22008 29452 22060 29504
rect 24492 29452 24544 29504
rect 32312 29520 32364 29572
rect 29184 29452 29236 29504
rect 44180 29452 44232 29504
rect 45836 29563 45888 29572
rect 45836 29529 45845 29563
rect 45845 29529 45879 29563
rect 45879 29529 45888 29563
rect 45836 29520 45888 29529
rect 47768 29520 47820 29572
rect 49148 29563 49200 29572
rect 49148 29529 49157 29563
rect 49157 29529 49191 29563
rect 49191 29529 49200 29563
rect 49148 29520 49200 29529
rect 45928 29495 45980 29504
rect 45928 29461 45937 29495
rect 45937 29461 45971 29495
rect 45971 29461 45980 29495
rect 45928 29452 45980 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 27950 29350 28002 29402
rect 28014 29350 28066 29402
rect 28078 29350 28130 29402
rect 28142 29350 28194 29402
rect 28206 29350 28258 29402
rect 37950 29350 38002 29402
rect 38014 29350 38066 29402
rect 38078 29350 38130 29402
rect 38142 29350 38194 29402
rect 38206 29350 38258 29402
rect 47950 29350 48002 29402
rect 48014 29350 48066 29402
rect 48078 29350 48130 29402
rect 48142 29350 48194 29402
rect 48206 29350 48258 29402
rect 14648 29248 14700 29300
rect 16028 29291 16080 29300
rect 16028 29257 16037 29291
rect 16037 29257 16071 29291
rect 16071 29257 16080 29291
rect 16028 29248 16080 29257
rect 16120 29248 16172 29300
rect 16304 29248 16356 29300
rect 16856 29248 16908 29300
rect 16028 29112 16080 29164
rect 19064 29180 19116 29232
rect 21456 29291 21508 29300
rect 21456 29257 21465 29291
rect 21465 29257 21499 29291
rect 21499 29257 21508 29291
rect 21456 29248 21508 29257
rect 21824 29248 21876 29300
rect 22376 29291 22428 29300
rect 22376 29257 22385 29291
rect 22385 29257 22419 29291
rect 22419 29257 22428 29291
rect 22376 29248 22428 29257
rect 25320 29248 25372 29300
rect 28816 29248 28868 29300
rect 29092 29291 29144 29300
rect 29092 29257 29101 29291
rect 29101 29257 29135 29291
rect 29135 29257 29144 29291
rect 29092 29248 29144 29257
rect 19892 29180 19944 29232
rect 20260 29180 20312 29232
rect 20628 29180 20680 29232
rect 24492 29223 24544 29232
rect 24492 29189 24501 29223
rect 24501 29189 24535 29223
rect 24535 29189 24544 29223
rect 24492 29180 24544 29189
rect 32404 29180 32456 29232
rect 32772 29180 32824 29232
rect 25320 29155 25372 29164
rect 25320 29121 25329 29155
rect 25329 29121 25363 29155
rect 25363 29121 25372 29155
rect 25320 29112 25372 29121
rect 28908 29112 28960 29164
rect 17224 29044 17276 29096
rect 17592 29087 17644 29096
rect 17592 29053 17601 29087
rect 17601 29053 17635 29087
rect 17635 29053 17644 29087
rect 17592 29044 17644 29053
rect 17684 29044 17736 29096
rect 18604 29044 18656 29096
rect 22652 29087 22704 29096
rect 22652 29053 22661 29087
rect 22661 29053 22695 29087
rect 22695 29053 22704 29087
rect 22652 29044 22704 29053
rect 27068 29044 27120 29096
rect 29184 29087 29236 29096
rect 29184 29053 29193 29087
rect 29193 29053 29227 29087
rect 29227 29053 29236 29087
rect 29184 29044 29236 29053
rect 17408 28908 17460 28960
rect 17684 28908 17736 28960
rect 21548 28908 21600 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 32950 28806 33002 28858
rect 33014 28806 33066 28858
rect 33078 28806 33130 28858
rect 33142 28806 33194 28858
rect 33206 28806 33258 28858
rect 42950 28806 43002 28858
rect 43014 28806 43066 28858
rect 43078 28806 43130 28858
rect 43142 28806 43194 28858
rect 43206 28806 43258 28858
rect 17592 28704 17644 28756
rect 18696 28704 18748 28756
rect 18788 28704 18840 28756
rect 19892 28704 19944 28756
rect 28448 28704 28500 28756
rect 19248 28636 19300 28688
rect 23756 28636 23808 28688
rect 1308 28568 1360 28620
rect 15936 28611 15988 28620
rect 15936 28577 15945 28611
rect 15945 28577 15979 28611
rect 15979 28577 15988 28611
rect 15936 28568 15988 28577
rect 17132 28611 17184 28620
rect 17132 28577 17141 28611
rect 17141 28577 17175 28611
rect 17175 28577 17184 28611
rect 17132 28568 17184 28577
rect 17408 28611 17460 28620
rect 17408 28577 17417 28611
rect 17417 28577 17451 28611
rect 17451 28577 17460 28611
rect 17408 28568 17460 28577
rect 21548 28611 21600 28620
rect 21548 28577 21557 28611
rect 21557 28577 21591 28611
rect 21591 28577 21600 28611
rect 21548 28568 21600 28577
rect 11060 28500 11112 28552
rect 15752 28543 15804 28552
rect 15752 28509 15761 28543
rect 15761 28509 15795 28543
rect 15795 28509 15804 28543
rect 15752 28500 15804 28509
rect 19524 28543 19576 28552
rect 19524 28509 19533 28543
rect 19533 28509 19567 28543
rect 19567 28509 19576 28543
rect 19524 28500 19576 28509
rect 22284 28500 22336 28552
rect 34796 28500 34848 28552
rect 49056 28543 49108 28552
rect 49056 28509 49065 28543
rect 49065 28509 49099 28543
rect 49099 28509 49108 28543
rect 49056 28500 49108 28509
rect 19064 28432 19116 28484
rect 20260 28475 20312 28484
rect 20260 28441 20269 28475
rect 20269 28441 20303 28475
rect 20303 28441 20312 28475
rect 20260 28432 20312 28441
rect 26516 28432 26568 28484
rect 15384 28407 15436 28416
rect 15384 28373 15393 28407
rect 15393 28373 15427 28407
rect 15427 28373 15436 28407
rect 15384 28364 15436 28373
rect 16948 28364 17000 28416
rect 17316 28364 17368 28416
rect 20168 28364 20220 28416
rect 20904 28407 20956 28416
rect 20904 28373 20913 28407
rect 20913 28373 20947 28407
rect 20947 28373 20956 28407
rect 20904 28364 20956 28373
rect 21364 28407 21416 28416
rect 21364 28373 21373 28407
rect 21373 28373 21407 28407
rect 21407 28373 21416 28407
rect 21364 28364 21416 28373
rect 43904 28364 43956 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 27950 28262 28002 28314
rect 28014 28262 28066 28314
rect 28078 28262 28130 28314
rect 28142 28262 28194 28314
rect 28206 28262 28258 28314
rect 37950 28262 38002 28314
rect 38014 28262 38066 28314
rect 38078 28262 38130 28314
rect 38142 28262 38194 28314
rect 38206 28262 38258 28314
rect 47950 28262 48002 28314
rect 48014 28262 48066 28314
rect 48078 28262 48130 28314
rect 48142 28262 48194 28314
rect 48206 28262 48258 28314
rect 15292 28203 15344 28212
rect 15292 28169 15301 28203
rect 15301 28169 15335 28203
rect 15335 28169 15344 28203
rect 15292 28160 15344 28169
rect 16948 28203 17000 28212
rect 16948 28169 16957 28203
rect 16957 28169 16991 28203
rect 16991 28169 17000 28203
rect 16948 28160 17000 28169
rect 19156 28160 19208 28212
rect 21364 28160 21416 28212
rect 31760 28092 31812 28144
rect 44088 28092 44140 28144
rect 11152 28024 11204 28076
rect 14740 28024 14792 28076
rect 16212 28024 16264 28076
rect 1308 27956 1360 28008
rect 16488 27956 16540 28008
rect 17316 28067 17368 28076
rect 17316 28033 17325 28067
rect 17325 28033 17359 28067
rect 17359 28033 17368 28067
rect 17316 28024 17368 28033
rect 18880 28024 18932 28076
rect 20076 28067 20128 28076
rect 20076 28033 20085 28067
rect 20085 28033 20119 28067
rect 20119 28033 20128 28067
rect 20076 28024 20128 28033
rect 21640 28024 21692 28076
rect 49332 28067 49384 28076
rect 49332 28033 49341 28067
rect 49341 28033 49375 28067
rect 49375 28033 49384 28067
rect 49332 28024 49384 28033
rect 18880 27888 18932 27940
rect 19708 27956 19760 28008
rect 20352 27999 20404 28008
rect 20352 27965 20361 27999
rect 20361 27965 20395 27999
rect 20395 27965 20404 27999
rect 20352 27956 20404 27965
rect 19248 27888 19300 27940
rect 36544 27888 36596 27940
rect 14740 27863 14792 27872
rect 14740 27829 14749 27863
rect 14749 27829 14783 27863
rect 14783 27829 14792 27863
rect 14740 27820 14792 27829
rect 45284 27863 45336 27872
rect 45284 27829 45293 27863
rect 45293 27829 45327 27863
rect 45327 27829 45336 27863
rect 45284 27820 45336 27829
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 32950 27718 33002 27770
rect 33014 27718 33066 27770
rect 33078 27718 33130 27770
rect 33142 27718 33194 27770
rect 33206 27718 33258 27770
rect 42950 27718 43002 27770
rect 43014 27718 43066 27770
rect 43078 27718 43130 27770
rect 43142 27718 43194 27770
rect 43206 27718 43258 27770
rect 16856 27548 16908 27600
rect 15844 27523 15896 27532
rect 15844 27489 15853 27523
rect 15853 27489 15887 27523
rect 15887 27489 15896 27523
rect 15844 27480 15896 27489
rect 16396 27480 16448 27532
rect 18420 27548 18472 27600
rect 19156 27548 19208 27600
rect 20444 27548 20496 27600
rect 17592 27480 17644 27532
rect 18604 27480 18656 27532
rect 15384 27412 15436 27464
rect 16948 27455 17000 27464
rect 16948 27421 16957 27455
rect 16957 27421 16991 27455
rect 16991 27421 17000 27455
rect 16948 27412 17000 27421
rect 18972 27412 19024 27464
rect 28356 27344 28408 27396
rect 46848 27344 46900 27396
rect 18420 27276 18472 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 27950 27174 28002 27226
rect 28014 27174 28066 27226
rect 28078 27174 28130 27226
rect 28142 27174 28194 27226
rect 28206 27174 28258 27226
rect 37950 27174 38002 27226
rect 38014 27174 38066 27226
rect 38078 27174 38130 27226
rect 38142 27174 38194 27226
rect 38206 27174 38258 27226
rect 47950 27174 48002 27226
rect 48014 27174 48066 27226
rect 48078 27174 48130 27226
rect 48142 27174 48194 27226
rect 48206 27174 48258 27226
rect 20904 27072 20956 27124
rect 19800 27004 19852 27056
rect 44548 27047 44600 27056
rect 44548 27013 44557 27047
rect 44557 27013 44591 27047
rect 44591 27013 44600 27047
rect 44548 27004 44600 27013
rect 940 26936 992 26988
rect 46756 26936 46808 26988
rect 21456 26868 21508 26920
rect 49148 26911 49200 26920
rect 49148 26877 49157 26911
rect 49157 26877 49191 26911
rect 49191 26877 49200 26911
rect 49148 26868 49200 26877
rect 44732 26843 44784 26852
rect 44732 26809 44741 26843
rect 44741 26809 44775 26843
rect 44775 26809 44784 26843
rect 44732 26800 44784 26809
rect 12440 26732 12492 26784
rect 22284 26732 22336 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 32950 26630 33002 26682
rect 33014 26630 33066 26682
rect 33078 26630 33130 26682
rect 33142 26630 33194 26682
rect 33206 26630 33258 26682
rect 42950 26630 43002 26682
rect 43014 26630 43066 26682
rect 43078 26630 43130 26682
rect 43142 26630 43194 26682
rect 43206 26630 43258 26682
rect 20168 26460 20220 26512
rect 18604 26435 18656 26444
rect 18604 26401 18613 26435
rect 18613 26401 18647 26435
rect 18647 26401 18656 26435
rect 18604 26392 18656 26401
rect 18788 26435 18840 26444
rect 18788 26401 18797 26435
rect 18797 26401 18831 26435
rect 18831 26401 18840 26435
rect 18788 26392 18840 26401
rect 48228 26392 48280 26444
rect 12624 26324 12676 26376
rect 18420 26324 18472 26376
rect 46480 26324 46532 26376
rect 1676 26299 1728 26308
rect 1676 26265 1685 26299
rect 1685 26265 1719 26299
rect 1719 26265 1728 26299
rect 1676 26256 1728 26265
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 27950 26086 28002 26138
rect 28014 26086 28066 26138
rect 28078 26086 28130 26138
rect 28142 26086 28194 26138
rect 28206 26086 28258 26138
rect 37950 26086 38002 26138
rect 38014 26086 38066 26138
rect 38078 26086 38130 26138
rect 38142 26086 38194 26138
rect 38206 26086 38258 26138
rect 47950 26086 48002 26138
rect 48014 26086 48066 26138
rect 48078 26086 48130 26138
rect 48142 26086 48194 26138
rect 48206 26086 48258 26138
rect 29644 25916 29696 25968
rect 37832 25848 37884 25900
rect 44272 25712 44324 25764
rect 39948 25644 40000 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 32950 25542 33002 25594
rect 33014 25542 33066 25594
rect 33078 25542 33130 25594
rect 33142 25542 33194 25594
rect 33206 25542 33258 25594
rect 42950 25542 43002 25594
rect 43014 25542 43066 25594
rect 43078 25542 43130 25594
rect 43142 25542 43194 25594
rect 43206 25542 43258 25594
rect 3424 25304 3476 25356
rect 940 25236 992 25288
rect 45928 25236 45980 25288
rect 49148 25279 49200 25288
rect 49148 25245 49157 25279
rect 49157 25245 49191 25279
rect 49191 25245 49200 25279
rect 49148 25236 49200 25245
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 27950 24998 28002 25050
rect 28014 24998 28066 25050
rect 28078 24998 28130 25050
rect 28142 24998 28194 25050
rect 28206 24998 28258 25050
rect 37950 24998 38002 25050
rect 38014 24998 38066 25050
rect 38078 24998 38130 25050
rect 38142 24998 38194 25050
rect 38206 24998 38258 25050
rect 47950 24998 48002 25050
rect 48014 24998 48066 25050
rect 48078 24998 48130 25050
rect 48142 24998 48194 25050
rect 48206 24998 48258 25050
rect 940 24760 992 24812
rect 28448 24760 28500 24812
rect 39304 24735 39356 24744
rect 39304 24701 39313 24735
rect 39313 24701 39347 24735
rect 39347 24701 39356 24735
rect 47768 24760 47820 24812
rect 39304 24692 39356 24701
rect 49148 24735 49200 24744
rect 49148 24701 49157 24735
rect 49157 24701 49191 24735
rect 49191 24701 49200 24735
rect 49148 24692 49200 24701
rect 44180 24624 44232 24676
rect 14832 24556 14884 24608
rect 46940 24556 46992 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 13360 24148 13412 24200
rect 33784 24148 33836 24200
rect 39396 24148 39448 24200
rect 45100 24080 45152 24132
rect 15660 24055 15712 24064
rect 15660 24021 15669 24055
rect 15669 24021 15703 24055
rect 15703 24021 15712 24055
rect 15660 24012 15712 24021
rect 43444 24012 43496 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 4896 23740 4948 23792
rect 33416 23740 33468 23792
rect 940 23672 992 23724
rect 32036 23672 32088 23724
rect 46848 23672 46900 23724
rect 49148 23647 49200 23656
rect 49148 23613 49157 23647
rect 49157 23613 49191 23647
rect 49191 23613 49200 23647
rect 49148 23604 49200 23613
rect 47032 23536 47084 23588
rect 36728 23511 36780 23520
rect 36728 23477 36737 23511
rect 36737 23477 36771 23511
rect 36771 23477 36780 23511
rect 36728 23468 36780 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 4804 23128 4856 23180
rect 940 23060 992 23112
rect 45284 23060 45336 23112
rect 49148 23035 49200 23044
rect 49148 23001 49157 23035
rect 49157 23001 49191 23035
rect 49191 23001 49200 23035
rect 49148 22992 49200 23001
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 43904 22015 43956 22024
rect 43904 21981 43913 22015
rect 43913 21981 43947 22015
rect 43947 21981 43956 22015
rect 43904 21972 43956 21981
rect 44732 21972 44784 22024
rect 49148 22015 49200 22024
rect 49148 21981 49157 22015
rect 49157 21981 49191 22015
rect 49191 21981 49200 22015
rect 49148 21972 49200 21981
rect 940 21904 992 21956
rect 44824 21904 44876 21956
rect 19156 21836 19208 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 940 21496 992 21548
rect 26700 21496 26752 21548
rect 44272 21496 44324 21548
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 42800 21360 42852 21412
rect 19892 21292 19944 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 32220 20816 32272 20868
rect 47768 20816 47820 20868
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 940 20408 992 20460
rect 44180 20408 44232 20460
rect 49148 20383 49200 20392
rect 49148 20349 49157 20383
rect 49157 20349 49191 20383
rect 49191 20349 49200 20383
rect 49148 20340 49200 20349
rect 16764 20204 16816 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 46940 19796 46992 19848
rect 940 19728 992 19780
rect 49148 19771 49200 19780
rect 49148 19737 49157 19771
rect 49157 19737 49191 19771
rect 49191 19737 49200 19771
rect 49148 19728 49200 19737
rect 17040 19660 17092 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 19984 19456 20036 19508
rect 22192 19456 22244 19508
rect 39948 19388 40000 19440
rect 16856 19320 16908 19372
rect 22284 19363 22336 19372
rect 22284 19329 22293 19363
rect 22293 19329 22327 19363
rect 22327 19329 22336 19363
rect 22284 19320 22336 19329
rect 32404 19320 32456 19372
rect 44272 19184 44324 19236
rect 46940 19184 46992 19236
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 940 18708 992 18760
rect 20168 18751 20220 18760
rect 20168 18717 20177 18751
rect 20177 18717 20211 18751
rect 20211 18717 20220 18751
rect 20168 18708 20220 18717
rect 40132 18751 40184 18760
rect 40132 18717 40141 18751
rect 40141 18717 40175 18751
rect 40175 18717 40184 18751
rect 40132 18708 40184 18717
rect 45100 18708 45152 18760
rect 49148 18751 49200 18760
rect 49148 18717 49157 18751
rect 49157 18717 49191 18751
rect 49191 18717 49200 18751
rect 49148 18708 49200 18717
rect 33416 18640 33468 18692
rect 47860 18640 47912 18692
rect 21916 18572 21968 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 47032 18232 47084 18284
rect 49148 18207 49200 18216
rect 49148 18173 49157 18207
rect 49157 18173 49191 18207
rect 49191 18173 49200 18207
rect 49148 18164 49200 18173
rect 26700 18028 26752 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 29184 17620 29236 17672
rect 43352 17552 43404 17604
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 940 17144 992 17196
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 27712 17144 27764 17196
rect 42800 17144 42852 17196
rect 49148 17119 49200 17128
rect 49148 17085 49157 17119
rect 49157 17085 49191 17119
rect 49191 17085 49200 17119
rect 49148 17076 49200 17085
rect 38292 17051 38344 17060
rect 38292 17017 38301 17051
rect 38301 17017 38335 17051
rect 38335 17017 38344 17051
rect 38292 17008 38344 17017
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 18328 16600 18380 16652
rect 38568 16600 38620 16652
rect 46204 16600 46256 16652
rect 43444 16532 43496 16584
rect 47768 16532 47820 16584
rect 940 16464 992 16516
rect 21824 16464 21876 16516
rect 49148 16507 49200 16516
rect 49148 16473 49157 16507
rect 49157 16473 49191 16507
rect 49191 16473 49200 16507
rect 49148 16464 49200 16473
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 23572 16124 23624 16176
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 22836 15920 22888 15972
rect 18972 15852 19024 15904
rect 38476 15920 38528 15972
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 25596 15512 25648 15564
rect 26240 15487 26292 15496
rect 26240 15453 26249 15487
rect 26249 15453 26283 15487
rect 26283 15453 26292 15487
rect 26240 15444 26292 15453
rect 44824 15444 44876 15496
rect 49148 15487 49200 15496
rect 49148 15453 49157 15487
rect 49157 15453 49191 15487
rect 49191 15453 49200 15487
rect 49148 15444 49200 15453
rect 940 15376 992 15428
rect 24676 15376 24728 15428
rect 15844 15308 15896 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 22652 15104 22704 15156
rect 25504 15036 25556 15088
rect 940 14968 992 15020
rect 28356 14900 28408 14952
rect 36728 15036 36780 15088
rect 44272 14968 44324 15020
rect 49148 14943 49200 14952
rect 49148 14909 49157 14943
rect 49157 14909 49191 14943
rect 49191 14909 49200 14943
rect 49148 14900 49200 14909
rect 21548 14764 21600 14816
rect 43812 14807 43864 14816
rect 43812 14773 43821 14807
rect 43821 14773 43855 14807
rect 43855 14773 43864 14807
rect 43812 14764 43864 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 30380 14467 30432 14476
rect 30380 14433 30389 14467
rect 30389 14433 30423 14467
rect 30423 14433 30432 14467
rect 30380 14424 30432 14433
rect 29828 14399 29880 14408
rect 29828 14365 29837 14399
rect 29837 14365 29871 14399
rect 29871 14365 29880 14399
rect 29828 14356 29880 14365
rect 27160 14288 27212 14340
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 940 13880 992 13932
rect 28632 13880 28684 13932
rect 47860 13880 47912 13932
rect 29184 13812 29236 13864
rect 37740 13855 37792 13864
rect 37740 13821 37749 13855
rect 37749 13821 37783 13855
rect 37783 13821 37792 13855
rect 37740 13812 37792 13821
rect 49148 13855 49200 13864
rect 49148 13821 49157 13855
rect 49157 13821 49191 13855
rect 49191 13821 49200 13855
rect 49148 13812 49200 13821
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 1860 13379 1912 13388
rect 1860 13345 1869 13379
rect 1869 13345 1903 13379
rect 1903 13345 1912 13379
rect 1860 13336 1912 13345
rect 15660 13336 15712 13388
rect 940 13268 992 13320
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 31024 13268 31076 13320
rect 43352 13268 43404 13320
rect 38568 13200 38620 13252
rect 49148 13243 49200 13252
rect 49148 13209 49157 13243
rect 49157 13209 49191 13243
rect 49191 13209 49200 13243
rect 49148 13200 49200 13209
rect 19524 13132 19576 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 23572 12928 23624 12980
rect 18420 12792 18472 12844
rect 24860 12792 24912 12844
rect 20076 12724 20128 12776
rect 38384 12631 38436 12640
rect 38384 12597 38393 12631
rect 38393 12597 38427 12631
rect 38427 12597 38436 12631
rect 38384 12588 38436 12597
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 24676 12384 24728 12436
rect 25504 12384 25556 12436
rect 27160 12384 27212 12436
rect 20168 12180 20220 12232
rect 27528 12248 27580 12300
rect 25320 12223 25372 12232
rect 25320 12189 25364 12223
rect 25364 12189 25372 12223
rect 25320 12180 25372 12189
rect 25504 12180 25556 12232
rect 46940 12180 46992 12232
rect 49148 12223 49200 12232
rect 49148 12189 49157 12223
rect 49157 12189 49191 12223
rect 49191 12189 49200 12223
rect 49148 12180 49200 12189
rect 940 12112 992 12164
rect 17500 12044 17552 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 940 11704 992 11756
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 37832 11704 37884 11756
rect 18604 11636 18656 11688
rect 20168 11679 20220 11688
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 49148 11679 49200 11688
rect 49148 11645 49157 11679
rect 49157 11645 49191 11679
rect 49191 11645 49200 11679
rect 49148 11636 49200 11645
rect 21824 11568 21876 11620
rect 21364 11500 21416 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 17316 11296 17368 11348
rect 21916 11203 21968 11212
rect 21916 11169 21925 11203
rect 21925 11169 21959 11203
rect 21959 11169 21968 11203
rect 21916 11160 21968 11169
rect 25320 11228 25372 11280
rect 22192 11160 22244 11212
rect 23388 11092 23440 11144
rect 25504 11160 25556 11212
rect 24584 11024 24636 11076
rect 26608 11024 26660 11076
rect 37464 11024 37516 11076
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 940 10616 992 10668
rect 15844 10480 15896 10532
rect 16396 10480 16448 10532
rect 38292 10616 38344 10668
rect 49148 10591 49200 10600
rect 49148 10557 49157 10591
rect 49157 10557 49191 10591
rect 49191 10557 49200 10591
rect 49148 10548 49200 10557
rect 37832 10480 37884 10532
rect 18972 10412 19024 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 27068 10072 27120 10124
rect 38476 10004 38528 10056
rect 940 9936 992 9988
rect 25412 9936 25464 9988
rect 14648 9868 14700 9920
rect 22376 9868 22428 9920
rect 33324 9936 33376 9988
rect 49148 9979 49200 9988
rect 49148 9945 49157 9979
rect 49157 9945 49191 9979
rect 49191 9945 49200 9979
rect 49148 9936 49200 9945
rect 27804 9911 27856 9920
rect 27804 9877 27813 9911
rect 27813 9877 27847 9911
rect 27847 9877 27856 9911
rect 27804 9868 27856 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 22376 9596 22428 9648
rect 20260 9528 20312 9580
rect 25228 9528 25280 9580
rect 22284 9503 22336 9512
rect 22284 9469 22293 9503
rect 22293 9469 22327 9503
rect 22327 9469 22336 9503
rect 22284 9460 22336 9469
rect 36452 9435 36504 9444
rect 36452 9401 36461 9435
rect 36461 9401 36495 9435
rect 36495 9401 36504 9435
rect 36452 9392 36504 9401
rect 25412 9324 25464 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 940 8916 992 8968
rect 46204 8916 46256 8968
rect 49148 8959 49200 8968
rect 49148 8925 49157 8959
rect 49157 8925 49191 8959
rect 49191 8925 49200 8959
rect 49148 8916 49200 8925
rect 28632 8780 28684 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 25320 8576 25372 8628
rect 25596 8619 25648 8628
rect 25596 8585 25605 8619
rect 25605 8585 25639 8619
rect 25639 8585 25648 8619
rect 25596 8576 25648 8585
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 24676 8440 24728 8492
rect 30748 8576 30800 8628
rect 33324 8576 33376 8628
rect 31024 8440 31076 8492
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 37740 8440 37792 8492
rect 27804 8372 27856 8424
rect 49148 8415 49200 8424
rect 49148 8381 49157 8415
rect 49157 8381 49191 8415
rect 49191 8381 49200 8415
rect 49148 8372 49200 8381
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 27620 8279 27672 8288
rect 27620 8245 27629 8279
rect 27629 8245 27663 8279
rect 27663 8245 27672 8279
rect 27620 8236 27672 8245
rect 34428 8279 34480 8288
rect 34428 8245 34437 8279
rect 34437 8245 34471 8279
rect 34471 8245 34480 8279
rect 34428 8236 34480 8245
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 22284 8032 22336 8084
rect 23388 8075 23440 8084
rect 23388 8041 23397 8075
rect 23397 8041 23431 8075
rect 23431 8041 23440 8075
rect 23388 8032 23440 8041
rect 24676 7828 24728 7880
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 940 7352 992 7404
rect 30748 7395 30800 7404
rect 30748 7361 30757 7395
rect 30757 7361 30791 7395
rect 30791 7361 30800 7395
rect 30748 7352 30800 7361
rect 38568 7352 38620 7404
rect 49148 7327 49200 7336
rect 49148 7293 49157 7327
rect 49157 7293 49191 7327
rect 49191 7293 49200 7327
rect 49148 7284 49200 7293
rect 18420 7216 18472 7268
rect 24860 7216 24912 7268
rect 20076 7148 20128 7200
rect 34428 7148 34480 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 38384 6740 38436 6792
rect 940 6672 992 6724
rect 49148 6715 49200 6724
rect 49148 6681 49157 6715
rect 49157 6681 49191 6715
rect 49191 6681 49200 6715
rect 49148 6672 49200 6681
rect 16948 6604 17000 6656
rect 19616 6647 19668 6656
rect 19616 6613 19625 6647
rect 19625 6613 19659 6647
rect 19659 6613 19668 6647
rect 19616 6604 19668 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 22284 5788 22336 5840
rect 14096 5720 14148 5772
rect 21364 5695 21416 5704
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 940 5584 992 5636
rect 9680 5584 9732 5636
rect 22376 5652 22428 5704
rect 24676 5695 24728 5704
rect 24676 5661 24685 5695
rect 24685 5661 24719 5695
rect 24719 5661 24728 5695
rect 24676 5652 24728 5661
rect 26608 5695 26660 5704
rect 26608 5661 26617 5695
rect 26617 5661 26651 5695
rect 26651 5661 26660 5695
rect 26608 5652 26660 5661
rect 43812 5652 43864 5704
rect 49148 5695 49200 5704
rect 49148 5661 49157 5695
rect 49157 5661 49191 5695
rect 49191 5661 49200 5695
rect 49148 5652 49200 5661
rect 22192 5584 22244 5636
rect 25228 5584 25280 5636
rect 28816 5584 28868 5636
rect 17224 5516 17276 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 18420 5244 18472 5296
rect 940 5176 992 5228
rect 37464 5176 37516 5228
rect 49148 5151 49200 5160
rect 49148 5117 49157 5151
rect 49157 5117 49191 5151
rect 49191 5117 49200 5151
rect 49148 5108 49200 5117
rect 15844 5040 15896 5092
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 14188 4632 14240 4684
rect 18604 4564 18656 4616
rect 23388 4564 23440 4616
rect 25596 4496 25648 4548
rect 11060 4428 11112 4480
rect 17868 4428 17920 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 940 4088 992 4140
rect 37832 4088 37884 4140
rect 49148 4063 49200 4072
rect 49148 4029 49157 4063
rect 49157 4029 49191 4063
rect 49191 4029 49200 4063
rect 49148 4020 49200 4029
rect 25320 3884 25372 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 36452 3476 36504 3528
rect 940 3408 992 3460
rect 25872 3408 25924 3460
rect 48596 3408 48648 3460
rect 49148 3451 49200 3460
rect 49148 3417 49157 3451
rect 49157 3417 49191 3451
rect 49191 3417 49200 3451
rect 49148 3408 49200 3417
rect 14740 3340 14792 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 28816 3043 28868 3052
rect 28816 3009 28825 3043
rect 28825 3009 28859 3043
rect 28859 3009 28868 3043
rect 28816 3000 28868 3009
rect 28724 2932 28776 2984
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 34428 2592 34480 2644
rect 28356 2524 28408 2576
rect 5540 2456 5592 2508
rect 8852 2456 8904 2508
rect 12164 2456 12216 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 18788 2456 18840 2508
rect 22100 2456 22152 2508
rect 25412 2456 25464 2508
rect 29828 2456 29880 2508
rect 2228 2388 2280 2440
rect 11060 2388 11112 2440
rect 14188 2388 14240 2440
rect 17868 2388 17920 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 32036 2388 32088 2440
rect 35348 2388 35400 2440
rect 13636 2320 13688 2372
rect 26240 2320 26292 2372
rect 38660 2431 38712 2440
rect 38660 2397 38669 2431
rect 38669 2397 38703 2431
rect 38703 2397 38712 2431
rect 38660 2388 38712 2397
rect 41972 2388 42024 2440
rect 45284 2320 45336 2372
rect 49148 2363 49200 2372
rect 49148 2329 49157 2363
rect 49157 2329 49191 2363
rect 49191 2329 49200 2363
rect 49148 2320 49200 2329
rect 9680 2252 9732 2304
rect 24768 2252 24820 2304
rect 45560 2295 45612 2304
rect 45560 2261 45569 2295
rect 45569 2261 45603 2295
rect 45603 2261 45612 2295
rect 45560 2252 45612 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 30748 2048 30800 2100
rect 45560 2048 45612 2100
<< metal2 >>
rect 1582 56200 1638 57000
rect 2226 56200 2282 57000
rect 2870 56200 2926 57000
rect 3514 56200 3570 57000
rect 4158 56200 4214 57000
rect 4802 56200 4858 57000
rect 5446 56200 5502 57000
rect 6090 56200 6146 57000
rect 6734 56200 6790 57000
rect 7378 56200 7434 57000
rect 8022 56200 8078 57000
rect 8666 56200 8722 57000
rect 9310 56200 9366 57000
rect 9954 56200 10010 57000
rect 10598 56200 10654 57000
rect 11242 56200 11298 57000
rect 11886 56200 11942 57000
rect 12530 56200 12586 57000
rect 13174 56200 13230 57000
rect 13818 56200 13874 57000
rect 14462 56200 14518 57000
rect 15106 56200 15162 57000
rect 15750 56200 15806 57000
rect 16394 56200 16450 57000
rect 17038 56200 17094 57000
rect 17682 56200 17738 57000
rect 18326 56200 18382 57000
rect 18970 56200 19026 57000
rect 19614 56200 19670 57000
rect 20258 56200 20314 57000
rect 20902 56200 20958 57000
rect 21546 56200 21602 57000
rect 22190 56200 22246 57000
rect 22834 56200 22890 57000
rect 23478 56200 23534 57000
rect 24122 56200 24178 57000
rect 24766 56200 24822 57000
rect 25410 56200 25466 57000
rect 26054 56200 26110 57000
rect 26698 56200 26754 57000
rect 27342 56200 27398 57000
rect 27986 56200 28042 57000
rect 28092 56222 28396 56250
rect 1596 52562 1624 56200
rect 2044 53576 2096 53582
rect 2044 53518 2096 53524
rect 1584 52556 1636 52562
rect 1584 52498 1636 52504
rect 1676 52488 1728 52494
rect 1676 52430 1728 52436
rect 1308 51468 1360 51474
rect 1308 51410 1360 51416
rect 1320 51377 1348 51410
rect 1306 51368 1362 51377
rect 1306 51303 1362 51312
rect 1308 50856 1360 50862
rect 1308 50798 1360 50804
rect 1320 50561 1348 50798
rect 1306 50552 1362 50561
rect 1306 50487 1362 50496
rect 1308 49768 1360 49774
rect 1306 49736 1308 49745
rect 1360 49736 1362 49745
rect 1306 49671 1362 49680
rect 1308 49292 1360 49298
rect 1308 49234 1360 49240
rect 1320 48929 1348 49234
rect 1306 48920 1362 48929
rect 1306 48855 1362 48864
rect 1308 48204 1360 48210
rect 1308 48146 1360 48152
rect 1320 48113 1348 48146
rect 1306 48104 1362 48113
rect 1306 48039 1362 48048
rect 1308 47592 1360 47598
rect 1308 47534 1360 47540
rect 1320 47297 1348 47534
rect 1306 47288 1362 47297
rect 1306 47223 1362 47232
rect 1308 46504 1360 46510
rect 1306 46472 1308 46481
rect 1360 46472 1362 46481
rect 1306 46407 1362 46416
rect 1308 46028 1360 46034
rect 1308 45970 1360 45976
rect 1320 45665 1348 45970
rect 1306 45656 1362 45665
rect 1306 45591 1362 45600
rect 1308 44940 1360 44946
rect 1308 44882 1360 44888
rect 1320 44849 1348 44882
rect 1306 44840 1362 44849
rect 1306 44775 1362 44784
rect 1308 43240 1360 43246
rect 1306 43208 1308 43217
rect 1360 43208 1362 43217
rect 1306 43143 1362 43152
rect 1308 42764 1360 42770
rect 1308 42706 1360 42712
rect 1320 42401 1348 42706
rect 1306 42392 1362 42401
rect 1306 42327 1362 42336
rect 1308 41676 1360 41682
rect 1308 41618 1360 41624
rect 1320 41585 1348 41618
rect 1306 41576 1362 41585
rect 1306 41511 1362 41520
rect 1308 41064 1360 41070
rect 1308 41006 1360 41012
rect 1320 40769 1348 41006
rect 1306 40760 1362 40769
rect 1306 40695 1362 40704
rect 1688 39642 1716 52430
rect 2056 44538 2084 53518
rect 2240 53174 2268 56200
rect 2884 53650 2912 56200
rect 3422 54632 3478 54641
rect 3422 54567 3478 54576
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 3330 53680 3386 53689
rect 2872 53644 2924 53650
rect 3330 53615 3386 53624
rect 2872 53586 2924 53592
rect 2228 53168 2280 53174
rect 2228 53110 2280 53116
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2044 44532 2096 44538
rect 2044 44474 2096 44480
rect 2044 44328 2096 44334
rect 2044 44270 2096 44276
rect 2056 44033 2084 44270
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2042 44024 2098 44033
rect 2950 44027 3258 44036
rect 2042 43959 2098 43968
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2044 39976 2096 39982
rect 2042 39944 2044 39953
rect 2096 39944 2098 39953
rect 3344 39914 3372 53615
rect 3436 51074 3464 54567
rect 3528 54262 3556 56200
rect 3516 54256 3568 54262
rect 3516 54198 3568 54204
rect 3606 53000 3662 53009
rect 3606 52935 3662 52944
rect 3436 51046 3556 51074
rect 3528 44441 3556 51046
rect 3514 44432 3570 44441
rect 3424 44396 3476 44402
rect 3514 44367 3570 44376
rect 3424 44338 3476 44344
rect 2042 39879 2098 39888
rect 3332 39908 3384 39914
rect 3332 39850 3384 39856
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 1676 39636 1728 39642
rect 1676 39578 1728 39584
rect 1308 39364 1360 39370
rect 1308 39306 1360 39312
rect 1320 39137 1348 39306
rect 1306 39128 1362 39137
rect 1306 39063 1362 39072
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 1768 38480 1820 38486
rect 1768 38422 1820 38428
rect 1308 38412 1360 38418
rect 1308 38354 1360 38360
rect 1320 38321 1348 38354
rect 1306 38312 1362 38321
rect 1306 38247 1362 38256
rect 1780 37874 1808 38422
rect 1768 37868 1820 37874
rect 1768 37810 1820 37816
rect 1308 37800 1360 37806
rect 1308 37742 1360 37748
rect 1320 37505 1348 37742
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 1306 37496 1362 37505
rect 2950 37499 3258 37508
rect 1306 37431 1362 37440
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1308 36712 1360 36718
rect 1306 36680 1308 36689
rect 1360 36680 1362 36689
rect 1306 36615 1362 36624
rect 1780 36378 1808 36722
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 2780 36100 2832 36106
rect 2780 36042 2832 36048
rect 2792 35873 2820 36042
rect 2778 35864 2834 35873
rect 3436 35834 3464 44338
rect 3620 41478 3648 52935
rect 4172 52562 4200 56200
rect 4816 53038 4844 56200
rect 4896 54188 4948 54194
rect 4896 54130 4948 54136
rect 4804 53032 4856 53038
rect 4804 52974 4856 52980
rect 4160 52556 4212 52562
rect 4160 52498 4212 52504
rect 4712 52488 4764 52494
rect 4712 52430 4764 52436
rect 4068 47660 4120 47666
rect 4068 47602 4120 47608
rect 4080 43450 4108 47602
rect 4724 43926 4752 52430
rect 4908 51610 4936 54130
rect 5460 54126 5488 56200
rect 5540 54256 5592 54262
rect 5540 54198 5592 54204
rect 5448 54120 5500 54126
rect 5448 54062 5500 54068
rect 4896 51604 4948 51610
rect 4896 51546 4948 51552
rect 5552 44470 5580 54198
rect 6104 53650 6132 56200
rect 6092 53644 6144 53650
rect 6092 53586 6144 53592
rect 5816 53100 5868 53106
rect 5816 53042 5868 53048
rect 5828 52154 5856 53042
rect 6748 52562 6776 56200
rect 7392 53038 7420 56200
rect 8036 55214 8064 56200
rect 7852 55186 8064 55214
rect 7852 53650 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8680 54262 8708 56200
rect 8668 54256 8720 54262
rect 8668 54198 8720 54204
rect 7840 53644 7892 53650
rect 7840 53586 7892 53592
rect 8484 53576 8536 53582
rect 8484 53518 8536 53524
rect 8392 53508 8444 53514
rect 8392 53450 8444 53456
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7380 53032 7432 53038
rect 7380 52974 7432 52980
rect 6736 52556 6788 52562
rect 6736 52498 6788 52504
rect 8300 52488 8352 52494
rect 8300 52430 8352 52436
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 5816 52148 5868 52154
rect 5816 52090 5868 52096
rect 7564 51400 7616 51406
rect 7564 51342 7616 51348
rect 5632 50924 5684 50930
rect 5632 50866 5684 50872
rect 5644 45082 5672 50866
rect 5724 49836 5776 49842
rect 5724 49778 5776 49784
rect 5632 45076 5684 45082
rect 5632 45018 5684 45024
rect 5540 44464 5592 44470
rect 5540 44406 5592 44412
rect 5356 44396 5408 44402
rect 5356 44338 5408 44344
rect 4712 43920 4764 43926
rect 4712 43862 4764 43868
rect 4804 43716 4856 43722
rect 4804 43658 4856 43664
rect 4068 43444 4120 43450
rect 4068 43386 4120 43392
rect 3608 41472 3660 41478
rect 3608 41414 3660 41420
rect 4816 36038 4844 43658
rect 5368 37194 5396 44338
rect 5736 43926 5764 49778
rect 5816 49224 5868 49230
rect 5816 49166 5868 49172
rect 5828 43994 5856 49166
rect 7576 45558 7604 51342
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 8312 51066 8340 52430
rect 8300 51060 8352 51066
rect 8300 51002 8352 51008
rect 8404 50454 8432 53450
rect 8392 50448 8444 50454
rect 8392 50390 8444 50396
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 8496 49434 8524 53518
rect 9324 52562 9352 56200
rect 9680 53100 9732 53106
rect 9680 53042 9732 53048
rect 9312 52556 9364 52562
rect 9312 52498 9364 52504
rect 9692 51066 9720 53042
rect 9968 53038 9996 56200
rect 10612 54262 10640 56200
rect 10600 54256 10652 54262
rect 10600 54198 10652 54204
rect 10508 54188 10560 54194
rect 10508 54130 10560 54136
rect 9956 53032 10008 53038
rect 9956 52974 10008 52980
rect 9772 52488 9824 52494
rect 9772 52430 9824 52436
rect 9680 51060 9732 51066
rect 9680 51002 9732 51008
rect 9588 50244 9640 50250
rect 9588 50186 9640 50192
rect 8484 49428 8536 49434
rect 8484 49370 8536 49376
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 8668 46572 8720 46578
rect 8668 46514 8720 46520
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7564 45552 7616 45558
rect 7564 45494 7616 45500
rect 6828 45280 6880 45286
rect 6828 45222 6880 45228
rect 6840 44470 6868 45222
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 6828 44464 6880 44470
rect 6828 44406 6880 44412
rect 6920 44192 6972 44198
rect 6920 44134 6972 44140
rect 5816 43988 5868 43994
rect 5816 43930 5868 43936
rect 5724 43920 5776 43926
rect 5724 43862 5776 43868
rect 6932 43382 6960 44134
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8680 43450 8708 46514
rect 9600 44538 9628 50186
rect 9784 49366 9812 52430
rect 10520 51066 10548 54130
rect 11256 53650 11284 56200
rect 11244 53644 11296 53650
rect 11244 53586 11296 53592
rect 11900 52562 11928 56200
rect 12440 53100 12492 53106
rect 12440 53042 12492 53048
rect 11888 52556 11940 52562
rect 11888 52498 11940 52504
rect 10692 52012 10744 52018
rect 10692 51954 10744 51960
rect 10508 51060 10560 51066
rect 10508 51002 10560 51008
rect 9956 50924 10008 50930
rect 9956 50866 10008 50872
rect 9772 49360 9824 49366
rect 9772 49302 9824 49308
rect 9968 45354 9996 50866
rect 10704 47802 10732 51954
rect 10968 51332 11020 51338
rect 10968 51274 11020 51280
rect 10692 47796 10744 47802
rect 10692 47738 10744 47744
rect 10980 46714 11008 51274
rect 11612 50924 11664 50930
rect 11612 50866 11664 50872
rect 11060 48136 11112 48142
rect 11060 48078 11112 48084
rect 10968 46708 11020 46714
rect 10968 46650 11020 46656
rect 11072 46170 11100 48078
rect 11060 46164 11112 46170
rect 11060 46106 11112 46112
rect 9956 45348 10008 45354
rect 9956 45290 10008 45296
rect 11624 45082 11652 50866
rect 12452 50522 12480 53042
rect 12544 53038 12572 56200
rect 13188 55214 13216 56200
rect 13188 55186 13400 55214
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 13372 53650 13400 55186
rect 13832 54262 13860 56200
rect 13820 54256 13872 54262
rect 13820 54198 13872 54204
rect 13728 54188 13780 54194
rect 13728 54130 13780 54136
rect 13360 53644 13412 53650
rect 13360 53586 13412 53592
rect 13544 53508 13596 53514
rect 13544 53450 13596 53456
rect 12532 53032 12584 53038
rect 12532 52974 12584 52980
rect 12808 52964 12860 52970
rect 12808 52906 12860 52912
rect 12440 50516 12492 50522
rect 12440 50458 12492 50464
rect 12820 49978 12848 52906
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 13556 49978 13584 53450
rect 13740 50454 13768 54130
rect 14476 52562 14504 56200
rect 15016 54188 15068 54194
rect 15016 54130 15068 54136
rect 14464 52556 14516 52562
rect 14464 52498 14516 52504
rect 13820 52488 13872 52494
rect 13820 52430 13872 52436
rect 13728 50448 13780 50454
rect 13728 50390 13780 50396
rect 13832 50386 13860 52430
rect 14924 50924 14976 50930
rect 14924 50866 14976 50872
rect 13820 50380 13872 50386
rect 13820 50322 13872 50328
rect 14832 50244 14884 50250
rect 14832 50186 14884 50192
rect 12808 49972 12860 49978
rect 12808 49914 12860 49920
rect 13544 49972 13596 49978
rect 13544 49914 13596 49920
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 11980 49156 12032 49162
rect 11980 49098 12032 49104
rect 11612 45076 11664 45082
rect 11612 45018 11664 45024
rect 11060 44872 11112 44878
rect 11060 44814 11112 44820
rect 9588 44532 9640 44538
rect 9588 44474 9640 44480
rect 11072 43994 11100 44814
rect 11888 44260 11940 44266
rect 11888 44202 11940 44208
rect 11060 43988 11112 43994
rect 11060 43930 11112 43936
rect 9588 43784 9640 43790
rect 9588 43726 9640 43732
rect 8668 43444 8720 43450
rect 8668 43386 8720 43392
rect 6920 43376 6972 43382
rect 6920 43318 6972 43324
rect 9496 43240 9548 43246
rect 9496 43182 9548 43188
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 9508 41750 9536 43182
rect 9496 41744 9548 41750
rect 9496 41686 9548 41692
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 8392 40112 8444 40118
rect 8392 40054 8444 40060
rect 9312 40112 9364 40118
rect 9312 40054 9364 40060
rect 7564 39840 7616 39846
rect 7564 39782 7616 39788
rect 7576 39642 7604 39782
rect 7564 39636 7616 39642
rect 7564 39578 7616 39584
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 8404 38554 8432 40054
rect 8392 38548 8444 38554
rect 8392 38490 8444 38496
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 8576 37664 8628 37670
rect 8576 37606 8628 37612
rect 5356 37188 5408 37194
rect 5356 37130 5408 37136
rect 5368 36786 5396 37130
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 4896 36780 4948 36786
rect 4896 36722 4948 36728
rect 5356 36780 5408 36786
rect 5356 36722 5408 36728
rect 4804 36032 4856 36038
rect 4804 35974 4856 35980
rect 2778 35799 2834 35808
rect 3424 35828 3476 35834
rect 3424 35770 3476 35776
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 1308 35148 1360 35154
rect 1308 35090 1360 35096
rect 1320 35057 1348 35090
rect 1306 35048 1362 35057
rect 1306 34983 1362 34992
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 2056 34241 2084 34478
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2042 34232 2098 34241
rect 2950 34235 3258 34244
rect 2042 34167 2098 34176
rect 1308 33448 1360 33454
rect 1306 33416 1308 33425
rect 1360 33416 1362 33425
rect 1306 33351 1362 33360
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 1308 32972 1360 32978
rect 1308 32914 1360 32920
rect 1320 32609 1348 32914
rect 1306 32600 1362 32609
rect 1306 32535 1362 32544
rect 1860 32224 1912 32230
rect 1860 32166 1912 32172
rect 1308 31884 1360 31890
rect 1308 31826 1360 31832
rect 1320 31793 1348 31826
rect 1306 31784 1362 31793
rect 1306 31719 1362 31728
rect 1308 31272 1360 31278
rect 1308 31214 1360 31220
rect 1320 30977 1348 31214
rect 1306 30968 1362 30977
rect 1306 30903 1362 30912
rect 1308 30184 1360 30190
rect 1306 30152 1308 30161
rect 1360 30152 1362 30161
rect 1306 30087 1362 30096
rect 1308 29708 1360 29714
rect 1308 29650 1360 29656
rect 1320 29345 1348 29650
rect 1306 29336 1362 29345
rect 1306 29271 1362 29280
rect 1308 28620 1360 28626
rect 1308 28562 1360 28568
rect 1320 28529 1348 28562
rect 1306 28520 1362 28529
rect 1306 28455 1362 28464
rect 1308 28008 1360 28014
rect 1308 27950 1360 27956
rect 1320 27713 1348 27950
rect 1306 27704 1362 27713
rect 1306 27639 1362 27648
rect 940 26988 992 26994
rect 940 26930 992 26936
rect 952 26897 980 26930
rect 938 26888 994 26897
rect 938 26823 994 26832
rect 1676 26308 1728 26314
rect 1676 26250 1728 26256
rect 1688 26081 1716 26250
rect 1674 26072 1730 26081
rect 1674 26007 1730 26016
rect 940 25288 992 25294
rect 938 25256 940 25265
rect 992 25256 994 25265
rect 938 25191 994 25200
rect 940 24812 992 24818
rect 940 24754 992 24760
rect 952 24449 980 24754
rect 938 24440 994 24449
rect 938 24375 994 24384
rect 940 23724 992 23730
rect 940 23666 992 23672
rect 952 23633 980 23666
rect 938 23624 994 23633
rect 938 23559 994 23568
rect 940 23112 992 23118
rect 940 23054 992 23060
rect 952 22817 980 23054
rect 938 22808 994 22817
rect 938 22743 994 22752
rect 938 21992 994 22001
rect 938 21927 940 21936
rect 992 21927 994 21936
rect 940 21898 992 21904
rect 940 21548 992 21554
rect 940 21490 992 21496
rect 952 21185 980 21490
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 940 20460 992 20466
rect 940 20402 992 20408
rect 952 20369 980 20402
rect 938 20360 994 20369
rect 938 20295 994 20304
rect 940 19780 992 19786
rect 940 19722 992 19728
rect 952 19553 980 19722
rect 938 19544 994 19553
rect 938 19479 994 19488
rect 940 18760 992 18766
rect 938 18728 940 18737
rect 992 18728 994 18737
rect 938 18663 994 18672
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17921 1624 18226
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 17105 980 17138
rect 938 17096 994 17105
rect 938 17031 994 17040
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 952 16289 980 16458
rect 938 16280 994 16289
rect 938 16215 994 16224
rect 938 15464 994 15473
rect 938 15399 940 15408
rect 992 15399 994 15408
rect 940 15370 992 15376
rect 940 15020 992 15026
rect 940 14962 992 14968
rect 952 14657 980 14962
rect 938 14648 994 14657
rect 938 14583 994 14592
rect 940 13932 992 13938
rect 940 13874 992 13880
rect 952 13841 980 13874
rect 938 13832 994 13841
rect 938 13767 994 13776
rect 1872 13394 1900 32166
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 3436 25362 3464 35770
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 4816 23186 4844 35974
rect 4908 23798 4936 36722
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8588 33522 8616 37606
rect 9324 35766 9352 40054
rect 9508 36174 9536 41686
rect 9600 40662 9628 43726
rect 11900 42362 11928 44202
rect 11888 42356 11940 42362
rect 11888 42298 11940 42304
rect 11992 41818 12020 49098
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13728 46572 13780 46578
rect 13728 46514 13780 46520
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 12256 45960 12308 45966
rect 12256 45902 12308 45908
rect 13634 45928 13690 45937
rect 12268 43926 12296 45902
rect 12532 45892 12584 45898
rect 13634 45863 13636 45872
rect 12532 45834 12584 45840
rect 13688 45863 13690 45872
rect 13636 45834 13688 45840
rect 12440 44396 12492 44402
rect 12440 44338 12492 44344
rect 12256 43920 12308 43926
rect 12256 43862 12308 43868
rect 11980 41812 12032 41818
rect 11980 41754 12032 41760
rect 11060 41608 11112 41614
rect 11060 41550 11112 41556
rect 11072 41274 11100 41550
rect 11060 41268 11112 41274
rect 11060 41210 11112 41216
rect 12256 41132 12308 41138
rect 12256 41074 12308 41080
rect 12268 40730 12296 41074
rect 12256 40724 12308 40730
rect 12256 40666 12308 40672
rect 9588 40656 9640 40662
rect 9588 40598 9640 40604
rect 9600 40118 9628 40598
rect 9588 40112 9640 40118
rect 9588 40054 9640 40060
rect 12452 38554 12480 44338
rect 12440 38548 12492 38554
rect 12440 38490 12492 38496
rect 12544 37262 12572 45834
rect 12808 45484 12860 45490
rect 12808 45426 12860 45432
rect 12820 40186 12848 45426
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 13544 44804 13596 44810
rect 13544 44746 13596 44752
rect 13450 44160 13506 44169
rect 12950 44092 13258 44101
rect 13450 44095 13506 44104
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 13360 42832 13412 42838
rect 13360 42774 13412 42780
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 13372 41546 13400 42774
rect 13360 41540 13412 41546
rect 13360 41482 13412 41488
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12808 40180 12860 40186
rect 12808 40122 12860 40128
rect 12716 39840 12768 39846
rect 12716 39782 12768 39788
rect 12728 39438 12756 39782
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12716 39432 12768 39438
rect 12716 39374 12768 39380
rect 12624 39296 12676 39302
rect 12624 39238 12676 39244
rect 12532 37256 12584 37262
rect 12532 37198 12584 37204
rect 11978 36680 12034 36689
rect 11978 36615 12034 36624
rect 11796 36372 11848 36378
rect 11796 36314 11848 36320
rect 9588 36236 9640 36242
rect 9588 36178 9640 36184
rect 9496 36168 9548 36174
rect 9496 36110 9548 36116
rect 9312 35760 9364 35766
rect 9312 35702 9364 35708
rect 9600 35630 9628 36178
rect 11060 36100 11112 36106
rect 11060 36042 11112 36048
rect 11072 36009 11100 36042
rect 11058 36000 11114 36009
rect 11058 35935 11114 35944
rect 9588 35624 9640 35630
rect 9588 35566 9640 35572
rect 9600 34542 9628 35566
rect 10784 35488 10836 35494
rect 10784 35430 10836 35436
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 10796 34066 10824 35430
rect 10874 35184 10930 35193
rect 10874 35119 10930 35128
rect 10888 35086 10916 35119
rect 10876 35080 10928 35086
rect 10876 35022 10928 35028
rect 10968 34944 11020 34950
rect 10968 34886 11020 34892
rect 10980 34610 11008 34886
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 10784 34060 10836 34066
rect 10784 34002 10836 34008
rect 11808 33998 11836 36314
rect 11992 36174 12020 36615
rect 12440 36236 12492 36242
rect 12440 36178 12492 36184
rect 11980 36168 12032 36174
rect 11980 36110 12032 36116
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 8576 33516 8628 33522
rect 8576 33458 8628 33464
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7380 31816 7432 31822
rect 7380 31758 7432 31764
rect 7392 30258 7420 31758
rect 11060 31680 11112 31686
rect 11060 31622 11112 31628
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 11072 31414 11100 31622
rect 11060 31408 11112 31414
rect 11060 31350 11112 31356
rect 10692 31340 10744 31346
rect 10692 31282 10744 31288
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 8680 29646 8708 31078
rect 10704 30938 10732 31282
rect 10692 30932 10744 30938
rect 10692 30874 10744 30880
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 8668 29640 8720 29646
rect 8668 29582 8720 29588
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 11072 28558 11100 30534
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 11164 28082 11192 30670
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 12452 26790 12480 36178
rect 12636 35834 12664 39238
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12716 38548 12768 38554
rect 12716 38490 12768 38496
rect 12728 38350 12756 38490
rect 12716 38344 12768 38350
rect 12716 38286 12768 38292
rect 12808 38344 12860 38350
rect 12808 38286 12860 38292
rect 12716 36916 12768 36922
rect 12716 36858 12768 36864
rect 12624 35828 12676 35834
rect 12624 35770 12676 35776
rect 12636 35154 12664 35770
rect 12624 35148 12676 35154
rect 12624 35090 12676 35096
rect 12532 34060 12584 34066
rect 12532 34002 12584 34008
rect 12544 31278 12572 34002
rect 12728 32314 12756 36858
rect 12820 32570 12848 38286
rect 12900 38208 12952 38214
rect 12900 38150 12952 38156
rect 12912 37874 12940 38150
rect 12900 37868 12952 37874
rect 12900 37810 12952 37816
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12992 37324 13044 37330
rect 12992 37266 13044 37272
rect 13004 36718 13032 37266
rect 13464 36922 13492 44095
rect 13556 40934 13584 44746
rect 13636 43716 13688 43722
rect 13636 43658 13688 43664
rect 13544 40928 13596 40934
rect 13544 40870 13596 40876
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13556 36802 13584 40870
rect 13648 40497 13676 43658
rect 13740 41818 13768 46514
rect 13820 45416 13872 45422
rect 13820 45358 13872 45364
rect 13728 41812 13780 41818
rect 13728 41754 13780 41760
rect 13832 41002 13860 45358
rect 14844 44266 14872 50186
rect 14936 44538 14964 50866
rect 15028 49842 15056 54130
rect 15120 53038 15148 56200
rect 15764 54262 15792 56200
rect 15752 54256 15804 54262
rect 15752 54198 15804 54204
rect 15384 54120 15436 54126
rect 15384 54062 15436 54068
rect 15200 53576 15252 53582
rect 15200 53518 15252 53524
rect 15108 53032 15160 53038
rect 15108 52974 15160 52980
rect 15212 51066 15240 53518
rect 15292 53100 15344 53106
rect 15292 53042 15344 53048
rect 15200 51060 15252 51066
rect 15200 51002 15252 51008
rect 15108 50380 15160 50386
rect 15108 50322 15160 50328
rect 15120 49910 15148 50322
rect 15108 49904 15160 49910
rect 15108 49846 15160 49852
rect 15016 49836 15068 49842
rect 15016 49778 15068 49784
rect 15200 49632 15252 49638
rect 15200 49574 15252 49580
rect 15108 47660 15160 47666
rect 15108 47602 15160 47608
rect 15016 44872 15068 44878
rect 15016 44814 15068 44820
rect 14924 44532 14976 44538
rect 14924 44474 14976 44480
rect 14832 44260 14884 44266
rect 14832 44202 14884 44208
rect 14556 43648 14608 43654
rect 14556 43590 14608 43596
rect 14280 41676 14332 41682
rect 14280 41618 14332 41624
rect 13820 40996 13872 41002
rect 13820 40938 13872 40944
rect 13634 40488 13690 40497
rect 13634 40423 13690 40432
rect 13636 39432 13688 39438
rect 13636 39374 13688 39380
rect 13464 36786 13584 36802
rect 13452 36780 13584 36786
rect 13504 36774 13584 36780
rect 13452 36722 13504 36728
rect 12992 36712 13044 36718
rect 12992 36654 13044 36660
rect 13360 36712 13412 36718
rect 13360 36654 13412 36660
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12992 34944 13044 34950
rect 13372 34898 13400 36654
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13464 36242 13492 36314
rect 13452 36236 13504 36242
rect 13452 36178 13504 36184
rect 13544 35148 13596 35154
rect 13544 35090 13596 35096
rect 12992 34886 13044 34892
rect 13004 34678 13032 34886
rect 13280 34870 13400 34898
rect 13452 34944 13504 34950
rect 13452 34886 13504 34892
rect 12992 34672 13044 34678
rect 12992 34614 13044 34620
rect 13280 34490 13308 34870
rect 13464 34746 13492 34886
rect 13452 34740 13504 34746
rect 13452 34682 13504 34688
rect 13280 34462 13492 34490
rect 13360 34400 13412 34406
rect 13360 34342 13412 34348
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12808 32564 12860 32570
rect 12808 32506 12860 32512
rect 12636 32286 12756 32314
rect 12532 31272 12584 31278
rect 12532 31214 12584 31220
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12636 26382 12664 32286
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12728 31958 12756 32166
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 12716 31952 12768 31958
rect 12716 31894 12768 31900
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 12820 30394 12848 30602
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13372 24206 13400 34342
rect 13464 33402 13492 34462
rect 13556 33522 13584 35090
rect 13648 34542 13676 39374
rect 13820 37664 13872 37670
rect 13820 37606 13872 37612
rect 13832 36854 13860 37606
rect 13912 37256 13964 37262
rect 13912 37198 13964 37204
rect 13820 36848 13872 36854
rect 13820 36790 13872 36796
rect 13728 35624 13780 35630
rect 13728 35566 13780 35572
rect 13636 34536 13688 34542
rect 13636 34478 13688 34484
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13464 33374 13676 33402
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13556 31482 13584 32846
rect 13648 31890 13676 33374
rect 13740 32366 13768 35566
rect 13924 34678 13952 37198
rect 14188 36032 14240 36038
rect 14188 35974 14240 35980
rect 14096 35488 14148 35494
rect 14096 35430 14148 35436
rect 14108 35154 14136 35430
rect 14096 35148 14148 35154
rect 14096 35090 14148 35096
rect 13912 34672 13964 34678
rect 13912 34614 13964 34620
rect 14200 33590 14228 35974
rect 14292 34202 14320 41618
rect 14372 39840 14424 39846
rect 14372 39782 14424 39788
rect 14384 38554 14412 39782
rect 14464 39500 14516 39506
rect 14464 39442 14516 39448
rect 14372 38548 14424 38554
rect 14372 38490 14424 38496
rect 14476 38418 14504 39442
rect 14464 38412 14516 38418
rect 14464 38354 14516 38360
rect 14476 37874 14504 38354
rect 14568 38185 14596 43590
rect 14648 40044 14700 40050
rect 14648 39986 14700 39992
rect 14660 39642 14688 39986
rect 14924 39976 14976 39982
rect 14924 39918 14976 39924
rect 14648 39636 14700 39642
rect 14648 39578 14700 39584
rect 14648 39024 14700 39030
rect 14648 38966 14700 38972
rect 14554 38176 14610 38185
rect 14554 38111 14610 38120
rect 14464 37868 14516 37874
rect 14464 37810 14516 37816
rect 14372 37460 14424 37466
rect 14372 37402 14424 37408
rect 14384 36242 14412 37402
rect 14476 37262 14504 37810
rect 14464 37256 14516 37262
rect 14464 37198 14516 37204
rect 14476 36922 14504 37198
rect 14464 36916 14516 36922
rect 14464 36858 14516 36864
rect 14372 36236 14424 36242
rect 14372 36178 14424 36184
rect 14568 36122 14596 38111
rect 14660 37330 14688 38966
rect 14832 38276 14884 38282
rect 14832 38218 14884 38224
rect 14648 37324 14700 37330
rect 14648 37266 14700 37272
rect 14660 36378 14688 37266
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 14648 36372 14700 36378
rect 14648 36314 14700 36320
rect 14568 36106 14688 36122
rect 14568 36100 14700 36106
rect 14568 36094 14648 36100
rect 14648 36042 14700 36048
rect 14556 36032 14608 36038
rect 14556 35974 14608 35980
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 14476 35018 14504 35430
rect 14464 35012 14516 35018
rect 14464 34954 14516 34960
rect 14568 34746 14596 35974
rect 14648 35760 14700 35766
rect 14646 35728 14648 35737
rect 14700 35728 14702 35737
rect 14646 35663 14702 35672
rect 14646 35184 14702 35193
rect 14646 35119 14702 35128
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 14372 34604 14424 34610
rect 14372 34546 14424 34552
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 14384 33658 14412 34546
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 14464 33856 14516 33862
rect 14464 33798 14516 33804
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 14188 33584 14240 33590
rect 14188 33526 14240 33532
rect 13728 32360 13780 32366
rect 13728 32302 13780 32308
rect 13636 31884 13688 31890
rect 13636 31826 13688 31832
rect 13648 31482 13676 31826
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13740 30122 13768 31214
rect 14476 30802 14504 33798
rect 14568 32502 14596 34342
rect 14660 33946 14688 35119
rect 14752 34746 14780 37062
rect 14844 35834 14872 38218
rect 14936 37670 14964 39918
rect 15028 39098 15056 44814
rect 15120 43450 15148 47602
rect 15212 47258 15240 49574
rect 15304 49434 15332 53042
rect 15396 52630 15424 54062
rect 16408 53650 16436 56200
rect 16396 53644 16448 53650
rect 16396 53586 16448 53592
rect 16212 53168 16264 53174
rect 16212 53110 16264 53116
rect 15384 52624 15436 52630
rect 15384 52566 15436 52572
rect 16224 49978 16252 53110
rect 17052 52562 17080 56200
rect 17696 53038 17724 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18340 53650 18368 56200
rect 18984 54262 19012 56200
rect 18972 54256 19024 54262
rect 18972 54198 19024 54204
rect 18328 53644 18380 53650
rect 18328 53586 18380 53592
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 19340 53100 19392 53106
rect 19340 53042 19392 53048
rect 17684 53032 17736 53038
rect 17684 52974 17736 52980
rect 17040 52556 17092 52562
rect 17040 52498 17092 52504
rect 16856 52488 16908 52494
rect 16856 52430 16908 52436
rect 16868 50522 16896 52430
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 19352 51066 19380 53042
rect 19628 53038 19656 56200
rect 20272 54126 20300 56200
rect 20720 54256 20772 54262
rect 20720 54198 20772 54204
rect 20260 54120 20312 54126
rect 20260 54062 20312 54068
rect 20732 53242 20760 54198
rect 20916 53514 20944 56200
rect 20904 53508 20956 53514
rect 20904 53450 20956 53456
rect 20720 53236 20772 53242
rect 20720 53178 20772 53184
rect 21560 53106 21588 56200
rect 22100 53712 22152 53718
rect 22100 53654 22152 53660
rect 19892 53100 19944 53106
rect 19892 53042 19944 53048
rect 21548 53100 21600 53106
rect 21548 53042 21600 53048
rect 19616 53032 19668 53038
rect 19616 52974 19668 52980
rect 19904 52698 19932 53042
rect 19892 52692 19944 52698
rect 19892 52634 19944 52640
rect 19432 52488 19484 52494
rect 19432 52430 19484 52436
rect 19340 51060 19392 51066
rect 19340 51002 19392 51008
rect 19248 50924 19300 50930
rect 19248 50866 19300 50872
rect 16856 50516 16908 50522
rect 16856 50458 16908 50464
rect 18328 50312 18380 50318
rect 18328 50254 18380 50260
rect 17500 50244 17552 50250
rect 17500 50186 17552 50192
rect 16120 49972 16172 49978
rect 16120 49914 16172 49920
rect 16212 49972 16264 49978
rect 16212 49914 16264 49920
rect 15292 49428 15344 49434
rect 15292 49370 15344 49376
rect 15200 47252 15252 47258
rect 15200 47194 15252 47200
rect 16132 43994 16160 49914
rect 16672 49700 16724 49706
rect 16672 49642 16724 49648
rect 16396 49156 16448 49162
rect 16396 49098 16448 49104
rect 16304 44804 16356 44810
rect 16304 44746 16356 44752
rect 16316 44402 16344 44746
rect 16304 44396 16356 44402
rect 16304 44338 16356 44344
rect 16120 43988 16172 43994
rect 16120 43930 16172 43936
rect 15936 43784 15988 43790
rect 15936 43726 15988 43732
rect 15948 43450 15976 43726
rect 15108 43444 15160 43450
rect 15108 43386 15160 43392
rect 15936 43444 15988 43450
rect 15936 43386 15988 43392
rect 15108 42628 15160 42634
rect 15108 42570 15160 42576
rect 15120 42362 15148 42570
rect 16408 42566 16436 49098
rect 16580 48000 16632 48006
rect 16580 47942 16632 47948
rect 16592 45490 16620 47942
rect 16580 45484 16632 45490
rect 16580 45426 16632 45432
rect 16488 43784 16540 43790
rect 16488 43726 16540 43732
rect 16396 42560 16448 42566
rect 16396 42502 16448 42508
rect 15108 42356 15160 42362
rect 15108 42298 15160 42304
rect 16304 42220 16356 42226
rect 16304 42162 16356 42168
rect 15292 42016 15344 42022
rect 15292 41958 15344 41964
rect 15108 40996 15160 41002
rect 15108 40938 15160 40944
rect 15016 39092 15068 39098
rect 15016 39034 15068 39040
rect 15120 38842 15148 40938
rect 15028 38814 15148 38842
rect 14924 37664 14976 37670
rect 14924 37606 14976 37612
rect 15028 37126 15056 38814
rect 15108 38752 15160 38758
rect 15108 38694 15160 38700
rect 15120 38214 15148 38694
rect 15108 38208 15160 38214
rect 15108 38150 15160 38156
rect 15120 37890 15148 38150
rect 15200 38004 15252 38010
rect 15304 37992 15332 41958
rect 16316 41818 16344 42162
rect 16304 41812 16356 41818
rect 16304 41754 16356 41760
rect 16028 41676 16080 41682
rect 16028 41618 16080 41624
rect 15660 40520 15712 40526
rect 15660 40462 15712 40468
rect 15936 40520 15988 40526
rect 15936 40462 15988 40468
rect 15476 40044 15528 40050
rect 15476 39986 15528 39992
rect 15252 37964 15332 37992
rect 15200 37946 15252 37952
rect 15120 37862 15424 37890
rect 15108 37324 15160 37330
rect 15108 37266 15160 37272
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 14924 36780 14976 36786
rect 14924 36722 14976 36728
rect 14832 35828 14884 35834
rect 14832 35770 14884 35776
rect 14936 35737 14964 36722
rect 15028 36174 15056 37062
rect 15120 36417 15148 37266
rect 15200 36576 15252 36582
rect 15200 36518 15252 36524
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15106 36408 15162 36417
rect 15106 36343 15162 36352
rect 15120 36242 15148 36343
rect 15108 36236 15160 36242
rect 15108 36178 15160 36184
rect 15016 36168 15068 36174
rect 15016 36110 15068 36116
rect 15106 36136 15162 36145
rect 15106 36071 15162 36080
rect 15120 36038 15148 36071
rect 15108 36032 15160 36038
rect 15108 35974 15160 35980
rect 14922 35728 14978 35737
rect 14922 35663 14978 35672
rect 14832 35012 14884 35018
rect 14832 34954 14884 34960
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 14844 34542 14872 34954
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14660 33918 14780 33946
rect 14648 33448 14700 33454
rect 14648 33390 14700 33396
rect 14556 32496 14608 32502
rect 14556 32438 14608 32444
rect 14464 30796 14516 30802
rect 14464 30738 14516 30744
rect 14096 30184 14148 30190
rect 14096 30126 14148 30132
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 14108 29646 14136 30126
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 4896 23792 4948 23798
rect 4896 23734 4948 23740
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 17105 2084 17138
rect 2042 17096 2098 17105
rect 2042 17031 2098 17040
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 13025 980 13262
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 938 13016 994 13025
rect 7950 13019 8258 13028
rect 938 12951 994 12960
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 938 12200 994 12209
rect 938 12135 940 12144
rect 992 12135 994 12144
rect 940 12106 992 12112
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11393 980 11698
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 938 11384 994 11393
rect 2950 11387 3258 11396
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 938 11319 994 11328
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10577 980 10610
rect 938 10568 994 10577
rect 938 10503 994 10512
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 940 9988 992 9994
rect 940 9930 992 9936
rect 952 9761 980 9930
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 938 9752 994 9761
rect 7950 9755 8258 9764
rect 938 9687 994 9696
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8129 1624 8434
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 1582 8120 1638 8129
rect 2950 8123 3258 8132
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 1582 8055 1638 8064
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 952 7313 980 7346
rect 938 7304 994 7313
rect 938 7239 994 7248
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6497 980 6666
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 938 6488 994 6497
rect 7950 6491 8258 6500
rect 938 6423 994 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 14108 5778 14136 29582
rect 14660 29306 14688 33390
rect 14752 31482 14780 33918
rect 15120 31754 15148 35974
rect 15212 35834 15240 36518
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 15304 35630 15332 36518
rect 15292 35624 15344 35630
rect 15292 35566 15344 35572
rect 15292 35148 15344 35154
rect 15292 35090 15344 35096
rect 15304 34066 15332 35090
rect 15396 34746 15424 37862
rect 15488 36378 15516 39986
rect 15672 39098 15700 40462
rect 15948 39506 15976 40462
rect 16040 40458 16068 41618
rect 16120 41540 16172 41546
rect 16120 41482 16172 41488
rect 16028 40452 16080 40458
rect 16028 40394 16080 40400
rect 15936 39500 15988 39506
rect 15936 39442 15988 39448
rect 15844 39364 15896 39370
rect 15844 39306 15896 39312
rect 15660 39092 15712 39098
rect 15660 39034 15712 39040
rect 15856 38758 15884 39306
rect 16132 39137 16160 41482
rect 16304 40044 16356 40050
rect 16304 39986 16356 39992
rect 16316 39506 16344 39986
rect 16304 39500 16356 39506
rect 16304 39442 16356 39448
rect 16212 39364 16264 39370
rect 16212 39306 16264 39312
rect 16118 39128 16174 39137
rect 16118 39063 16174 39072
rect 16028 38888 16080 38894
rect 16028 38830 16080 38836
rect 16120 38888 16172 38894
rect 16120 38830 16172 38836
rect 15844 38752 15896 38758
rect 15844 38694 15896 38700
rect 15844 37256 15896 37262
rect 15844 37198 15896 37204
rect 15752 37188 15804 37194
rect 15752 37130 15804 37136
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 15476 36100 15528 36106
rect 15476 36042 15528 36048
rect 15384 34740 15436 34746
rect 15384 34682 15436 34688
rect 15292 34060 15344 34066
rect 15292 34002 15344 34008
rect 15304 32978 15332 34002
rect 15384 33856 15436 33862
rect 15384 33798 15436 33804
rect 15292 32972 15344 32978
rect 15292 32914 15344 32920
rect 15304 32366 15332 32914
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 14936 31726 15148 31754
rect 14740 31476 14792 31482
rect 14740 31418 14792 31424
rect 14740 31272 14792 31278
rect 14740 31214 14792 31220
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14752 29186 14780 31214
rect 14832 31136 14884 31142
rect 14832 31078 14884 31084
rect 14844 30734 14872 31078
rect 14832 30728 14884 30734
rect 14832 30670 14884 30676
rect 14936 30546 14964 31726
rect 15016 30796 15068 30802
rect 15016 30738 15068 30744
rect 14660 29158 14780 29186
rect 14844 30518 14964 30546
rect 14660 9926 14688 29158
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14752 27878 14780 28018
rect 14740 27872 14792 27878
rect 14740 27814 14792 27820
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 938 5672 994 5681
rect 938 5607 940 5616
rect 992 5607 994 5616
rect 9680 5636 9732 5642
rect 940 5578 992 5584
rect 9680 5578 9732 5584
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4865 980 5170
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 938 4856 994 4865
rect 2950 4859 3258 4868
rect 938 4791 994 4800
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 4049 980 4082
rect 938 4040 994 4049
rect 938 3975 994 3984
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 3233 980 3402
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 938 3224 994 3233
rect 7950 3227 8258 3236
rect 938 3159 994 3168
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2240 800 2268 2382
rect 5552 800 5580 2450
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8864 800 8892 2450
rect 9692 2310 9720 5578
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 2446 11100 4422
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 12176 800 12204 2450
rect 13648 2378 13676 4966
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14200 2446 14228 4626
rect 14752 3398 14780 27814
rect 14844 24614 14872 30518
rect 15028 30410 15056 30738
rect 15212 30734 15240 31826
rect 15396 31754 15424 33798
rect 15304 31726 15424 31754
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 14936 30382 15056 30410
rect 14936 29578 14964 30382
rect 15212 30274 15240 30670
rect 15028 30246 15240 30274
rect 15028 29714 15056 30246
rect 15016 29708 15068 29714
rect 15016 29650 15068 29656
rect 14924 29572 14976 29578
rect 14924 29514 14976 29520
rect 15304 28218 15332 31726
rect 15488 31346 15516 36042
rect 15764 35766 15792 37130
rect 15856 36718 15884 37198
rect 15844 36712 15896 36718
rect 15844 36654 15896 36660
rect 15934 36408 15990 36417
rect 15934 36343 15990 36352
rect 15660 35760 15712 35766
rect 15660 35702 15712 35708
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 15672 35222 15700 35702
rect 15660 35216 15712 35222
rect 15660 35158 15712 35164
rect 15844 35080 15896 35086
rect 15844 35022 15896 35028
rect 15856 34542 15884 35022
rect 15844 34536 15896 34542
rect 15844 34478 15896 34484
rect 15568 34468 15620 34474
rect 15568 34410 15620 34416
rect 15580 31754 15608 34410
rect 15948 32842 15976 36343
rect 16040 35834 16068 38830
rect 16132 37890 16160 38830
rect 16224 38826 16252 39306
rect 16212 38820 16264 38826
rect 16212 38762 16264 38768
rect 16224 38486 16252 38762
rect 16212 38480 16264 38486
rect 16212 38422 16264 38428
rect 16132 37862 16252 37890
rect 16120 37800 16172 37806
rect 16120 37742 16172 37748
rect 16132 37074 16160 37742
rect 16224 37330 16252 37862
rect 16302 37768 16358 37777
rect 16302 37703 16358 37712
rect 16212 37324 16264 37330
rect 16212 37266 16264 37272
rect 16212 37120 16264 37126
rect 16132 37068 16212 37074
rect 16132 37062 16264 37068
rect 16132 37046 16252 37062
rect 16132 36242 16160 37046
rect 16120 36236 16172 36242
rect 16120 36178 16172 36184
rect 16316 36106 16344 37703
rect 16500 37670 16528 43726
rect 16684 42634 16712 49642
rect 17512 44538 17540 50186
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18340 45354 18368 50254
rect 18972 49836 19024 49842
rect 18972 49778 19024 49784
rect 18880 48544 18932 48550
rect 18880 48486 18932 48492
rect 18512 48136 18564 48142
rect 18512 48078 18564 48084
rect 18328 45348 18380 45354
rect 18328 45290 18380 45296
rect 18524 44878 18552 48078
rect 18604 45824 18656 45830
rect 18604 45766 18656 45772
rect 18512 44872 18564 44878
rect 18512 44814 18564 44820
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17500 44532 17552 44538
rect 17500 44474 17552 44480
rect 17960 44260 18012 44266
rect 17960 44202 18012 44208
rect 17972 44146 18000 44202
rect 17880 44118 18000 44146
rect 18328 44192 18380 44198
rect 18328 44134 18380 44140
rect 17880 43858 17908 44118
rect 16856 43852 16908 43858
rect 16856 43794 16908 43800
rect 17868 43852 17920 43858
rect 18340 43840 18368 44134
rect 18420 43852 18472 43858
rect 18340 43812 18420 43840
rect 17868 43794 17920 43800
rect 18420 43794 18472 43800
rect 16672 42628 16724 42634
rect 16672 42570 16724 42576
rect 16868 42226 16896 43794
rect 18420 43716 18472 43722
rect 18420 43658 18472 43664
rect 18328 43648 18380 43654
rect 18328 43590 18380 43596
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17776 43308 17828 43314
rect 17776 43250 17828 43256
rect 17040 43172 17092 43178
rect 17040 43114 17092 43120
rect 16856 42220 16908 42226
rect 16856 42162 16908 42168
rect 16856 42084 16908 42090
rect 16856 42026 16908 42032
rect 16868 40712 16896 42026
rect 17052 41478 17080 43114
rect 17500 42696 17552 42702
rect 17500 42638 17552 42644
rect 17132 42152 17184 42158
rect 17132 42094 17184 42100
rect 17040 41472 17092 41478
rect 17040 41414 17092 41420
rect 17144 40730 17172 42094
rect 17132 40724 17184 40730
rect 16868 40684 17080 40712
rect 16948 40588 17000 40594
rect 16948 40530 17000 40536
rect 16672 40452 16724 40458
rect 16672 40394 16724 40400
rect 16856 40452 16908 40458
rect 16856 40394 16908 40400
rect 16684 39642 16712 40394
rect 16868 40118 16896 40394
rect 16856 40112 16908 40118
rect 16856 40054 16908 40060
rect 16672 39636 16724 39642
rect 16672 39578 16724 39584
rect 16868 39302 16896 40054
rect 16580 39296 16632 39302
rect 16580 39238 16632 39244
rect 16856 39296 16908 39302
rect 16856 39238 16908 39244
rect 16592 38264 16620 39238
rect 16960 39098 16988 40530
rect 16948 39092 17000 39098
rect 16948 39034 17000 39040
rect 17052 38486 17080 40684
rect 17132 40666 17184 40672
rect 17132 40588 17184 40594
rect 17132 40530 17184 40536
rect 17144 39030 17172 40530
rect 17316 40180 17368 40186
rect 17316 40122 17368 40128
rect 17328 39098 17356 40122
rect 17316 39092 17368 39098
rect 17316 39034 17368 39040
rect 17132 39024 17184 39030
rect 17132 38966 17184 38972
rect 17040 38480 17092 38486
rect 17040 38422 17092 38428
rect 16856 38344 16908 38350
rect 16856 38286 16908 38292
rect 16672 38276 16724 38282
rect 16592 38236 16672 38264
rect 16672 38218 16724 38224
rect 16684 37942 16712 38218
rect 16672 37936 16724 37942
rect 16672 37878 16724 37884
rect 16488 37664 16540 37670
rect 16488 37606 16540 37612
rect 16684 37194 16712 37878
rect 16672 37188 16724 37194
rect 16672 37130 16724 37136
rect 16684 36854 16712 37130
rect 16672 36848 16724 36854
rect 16672 36790 16724 36796
rect 16762 36816 16818 36825
rect 16762 36751 16764 36760
rect 16816 36751 16818 36760
rect 16764 36722 16816 36728
rect 16868 36718 16896 38286
rect 16856 36712 16908 36718
rect 16856 36654 16908 36660
rect 16488 36576 16540 36582
rect 16488 36518 16540 36524
rect 16304 36100 16356 36106
rect 16304 36042 16356 36048
rect 16396 36032 16448 36038
rect 16396 35974 16448 35980
rect 16028 35828 16080 35834
rect 16028 35770 16080 35776
rect 16026 35728 16082 35737
rect 16026 35663 16082 35672
rect 16040 35018 16068 35663
rect 16120 35488 16172 35494
rect 16120 35430 16172 35436
rect 16028 35012 16080 35018
rect 16028 34954 16080 34960
rect 16040 33930 16068 34954
rect 16028 33924 16080 33930
rect 16028 33866 16080 33872
rect 15936 32836 15988 32842
rect 15856 32796 15936 32824
rect 15580 31726 15700 31754
rect 15672 31482 15700 31726
rect 15660 31476 15712 31482
rect 15660 31418 15712 31424
rect 15752 31408 15804 31414
rect 15752 31350 15804 31356
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 15764 28558 15792 31350
rect 15856 31278 15884 32796
rect 15936 32778 15988 32784
rect 16040 32502 16068 33866
rect 16028 32496 16080 32502
rect 16028 32438 16080 32444
rect 16028 32224 16080 32230
rect 16028 32166 16080 32172
rect 16040 31754 16068 32166
rect 15948 31726 16068 31754
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15948 31142 15976 31726
rect 16132 31414 16160 35430
rect 16212 35216 16264 35222
rect 16212 35158 16264 35164
rect 16224 34678 16252 35158
rect 16408 35154 16436 35974
rect 16396 35148 16448 35154
rect 16396 35090 16448 35096
rect 16212 34672 16264 34678
rect 16212 34614 16264 34620
rect 16304 34604 16356 34610
rect 16304 34546 16356 34552
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 16224 32570 16252 32914
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 16120 31408 16172 31414
rect 16120 31350 16172 31356
rect 16212 31272 16264 31278
rect 16212 31214 16264 31220
rect 16028 31204 16080 31210
rect 16028 31146 16080 31152
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 15844 30592 15896 30598
rect 15844 30534 15896 30540
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15396 27470 15424 28358
rect 15856 27538 15884 30534
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15948 29510 15976 29990
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15948 28626 15976 29446
rect 16040 29306 16068 31146
rect 16224 31142 16252 31214
rect 16212 31136 16264 31142
rect 16212 31078 16264 31084
rect 16224 30190 16252 31078
rect 16212 30184 16264 30190
rect 16212 30126 16264 30132
rect 16028 29300 16080 29306
rect 16028 29242 16080 29248
rect 16120 29300 16172 29306
rect 16120 29242 16172 29248
rect 16026 29200 16082 29209
rect 16026 29135 16028 29144
rect 16080 29135 16082 29144
rect 16028 29106 16080 29112
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15384 27464 15436 27470
rect 15384 27406 15436 27412
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15672 13394 15700 24006
rect 16132 22094 16160 29242
rect 16224 28082 16252 30126
rect 16316 30054 16344 34546
rect 16396 34536 16448 34542
rect 16396 34478 16448 34484
rect 16408 33658 16436 34478
rect 16396 33652 16448 33658
rect 16396 33594 16448 33600
rect 16500 33522 16528 36518
rect 16946 36408 17002 36417
rect 16946 36343 17002 36352
rect 16854 36272 16910 36281
rect 16960 36242 16988 36343
rect 16854 36207 16856 36216
rect 16908 36207 16910 36216
rect 16948 36236 17000 36242
rect 16856 36178 16908 36184
rect 16948 36178 17000 36184
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16396 32768 16448 32774
rect 16396 32710 16448 32716
rect 16408 32502 16436 32710
rect 16396 32496 16448 32502
rect 16396 32438 16448 32444
rect 16408 31754 16436 32438
rect 16592 32026 16620 33798
rect 16684 33114 16712 34546
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 16396 31748 16448 31754
rect 16396 31690 16448 31696
rect 16488 31680 16540 31686
rect 16488 31622 16540 31628
rect 16396 30660 16448 30666
rect 16396 30602 16448 30608
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16316 29306 16344 29990
rect 16408 29510 16436 30602
rect 16396 29504 16448 29510
rect 16396 29446 16448 29452
rect 16304 29300 16356 29306
rect 16304 29242 16356 29248
rect 16302 29200 16358 29209
rect 16302 29135 16358 29144
rect 16212 28076 16264 28082
rect 16212 28018 16264 28024
rect 15856 22066 16160 22094
rect 16316 22094 16344 29135
rect 16408 27538 16436 29446
rect 16500 28014 16528 31622
rect 16672 30796 16724 30802
rect 16672 30738 16724 30744
rect 16684 30326 16712 30738
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16684 29578 16712 30262
rect 16672 29572 16724 29578
rect 16672 29514 16724 29520
rect 16488 28008 16540 28014
rect 16488 27950 16540 27956
rect 16396 27532 16448 27538
rect 16396 27474 16448 27480
rect 16316 22066 16436 22094
rect 15856 15366 15884 22066
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 16408 10538 16436 22066
rect 16776 20262 16804 36110
rect 16868 32042 16896 36178
rect 17052 36038 17080 38422
rect 17408 38208 17460 38214
rect 17406 38176 17408 38185
rect 17460 38176 17462 38185
rect 17406 38111 17462 38120
rect 17314 37224 17370 37233
rect 17314 37159 17370 37168
rect 17132 36712 17184 36718
rect 17132 36654 17184 36660
rect 17040 36032 17092 36038
rect 17040 35974 17092 35980
rect 17144 35766 17172 36654
rect 17224 36304 17276 36310
rect 17224 36246 17276 36252
rect 17132 35760 17184 35766
rect 17132 35702 17184 35708
rect 17144 34202 17172 35702
rect 17132 34196 17184 34202
rect 17132 34138 17184 34144
rect 17132 32768 17184 32774
rect 17132 32710 17184 32716
rect 16868 32014 17080 32042
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 16868 30802 16896 31690
rect 16856 30796 16908 30802
rect 16856 30738 16908 30744
rect 16856 29640 16908 29646
rect 16856 29582 16908 29588
rect 16868 29306 16896 29582
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 28218 16988 28358
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 16856 27600 16908 27606
rect 16856 27542 16908 27548
rect 16946 27568 17002 27577
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16868 19378 16896 27542
rect 16946 27503 17002 27512
rect 16960 27470 16988 27503
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 15856 5098 15884 10474
rect 16960 6662 16988 27406
rect 17052 19718 17080 32014
rect 17144 31362 17172 32710
rect 17236 31482 17264 36246
rect 17328 36009 17356 37159
rect 17420 36378 17448 38111
rect 17512 36553 17540 42638
rect 17684 42152 17736 42158
rect 17684 42094 17736 42100
rect 17592 41472 17644 41478
rect 17592 41414 17644 41420
rect 17604 37262 17632 41414
rect 17696 40118 17724 42094
rect 17684 40112 17736 40118
rect 17684 40054 17736 40060
rect 17684 39908 17736 39914
rect 17684 39850 17736 39856
rect 17696 38962 17724 39850
rect 17788 39642 17816 43250
rect 18340 43246 18368 43590
rect 18328 43240 18380 43246
rect 18328 43182 18380 43188
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 18340 42090 18368 43182
rect 18432 42294 18460 43658
rect 18512 43104 18564 43110
rect 18512 43046 18564 43052
rect 18420 42288 18472 42294
rect 18420 42230 18472 42236
rect 18328 42084 18380 42090
rect 18328 42026 18380 42032
rect 18524 41614 18552 43046
rect 18616 42770 18644 45766
rect 18696 45008 18748 45014
rect 18696 44950 18748 44956
rect 18708 44554 18736 44950
rect 18708 44526 18828 44554
rect 18696 43852 18748 43858
rect 18696 43794 18748 43800
rect 18604 42764 18656 42770
rect 18604 42706 18656 42712
rect 18512 41608 18564 41614
rect 18512 41550 18564 41556
rect 18708 41414 18736 43794
rect 18524 41386 18736 41414
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17868 40724 17920 40730
rect 17868 40666 17920 40672
rect 17776 39636 17828 39642
rect 17776 39578 17828 39584
rect 17880 39438 17908 40666
rect 18420 40384 18472 40390
rect 18420 40326 18472 40332
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 18432 39953 18460 40326
rect 18418 39944 18474 39953
rect 18418 39879 18474 39888
rect 17868 39432 17920 39438
rect 17868 39374 17920 39380
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17774 39128 17830 39137
rect 17950 39131 18258 39140
rect 17774 39063 17776 39072
rect 17828 39063 17830 39072
rect 18418 39128 18474 39137
rect 18418 39063 18420 39072
rect 17776 39034 17828 39040
rect 18472 39063 18474 39072
rect 18420 39034 18472 39040
rect 17684 38956 17736 38962
rect 17684 38898 17736 38904
rect 18328 38956 18380 38962
rect 18328 38898 18380 38904
rect 17868 38548 17920 38554
rect 17868 38490 17920 38496
rect 17592 37256 17644 37262
rect 17592 37198 17644 37204
rect 17684 37120 17736 37126
rect 17604 37080 17684 37108
rect 17498 36544 17554 36553
rect 17498 36479 17554 36488
rect 17408 36372 17460 36378
rect 17408 36314 17460 36320
rect 17314 36000 17370 36009
rect 17314 35935 17370 35944
rect 17328 32434 17356 35935
rect 17500 35148 17552 35154
rect 17500 35090 17552 35096
rect 17512 34610 17540 35090
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17408 33312 17460 33318
rect 17408 33254 17460 33260
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17316 32292 17368 32298
rect 17316 32234 17368 32240
rect 17328 32026 17356 32234
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 17420 31482 17448 33254
rect 17512 32774 17540 34546
rect 17604 34066 17632 37080
rect 17684 37062 17736 37068
rect 17776 35624 17828 35630
rect 17776 35566 17828 35572
rect 17684 34128 17736 34134
rect 17684 34070 17736 34076
rect 17592 34060 17644 34066
rect 17592 34002 17644 34008
rect 17696 33590 17724 34070
rect 17684 33584 17736 33590
rect 17684 33526 17736 33532
rect 17696 33454 17724 33526
rect 17788 33454 17816 35566
rect 17880 35086 17908 38490
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 17972 35698 18000 35770
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 18236 35692 18288 35698
rect 18236 35634 18288 35640
rect 17868 35080 17920 35086
rect 18248 35057 18276 35634
rect 18340 35154 18368 38898
rect 18524 38010 18552 41386
rect 18800 41206 18828 44526
rect 18892 43314 18920 48486
rect 18880 43308 18932 43314
rect 18880 43250 18932 43256
rect 18984 42566 19012 49778
rect 19156 47184 19208 47190
rect 19156 47126 19208 47132
rect 19064 44736 19116 44742
rect 19064 44678 19116 44684
rect 18972 42560 19024 42566
rect 18972 42502 19024 42508
rect 18880 41608 18932 41614
rect 18880 41550 18932 41556
rect 18788 41200 18840 41206
rect 18788 41142 18840 41148
rect 18788 41064 18840 41070
rect 18788 41006 18840 41012
rect 18696 40452 18748 40458
rect 18696 40394 18748 40400
rect 18708 39522 18736 40394
rect 18800 39982 18828 41006
rect 18892 40186 18920 41550
rect 18880 40180 18932 40186
rect 18880 40122 18932 40128
rect 18788 39976 18840 39982
rect 18788 39918 18840 39924
rect 18970 39944 19026 39953
rect 18970 39879 19026 39888
rect 18708 39494 18828 39522
rect 18696 39364 18748 39370
rect 18696 39306 18748 39312
rect 18604 39296 18656 39302
rect 18602 39264 18604 39273
rect 18656 39264 18658 39273
rect 18602 39199 18658 39208
rect 18604 38276 18656 38282
rect 18604 38218 18656 38224
rect 18512 38004 18564 38010
rect 18512 37946 18564 37952
rect 18420 37324 18472 37330
rect 18420 37266 18472 37272
rect 18432 36904 18460 37266
rect 18512 36916 18564 36922
rect 18432 36876 18512 36904
rect 18512 36858 18564 36864
rect 18512 36780 18564 36786
rect 18512 36722 18564 36728
rect 18524 36378 18552 36722
rect 18512 36372 18564 36378
rect 18512 36314 18564 36320
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 17868 35022 17920 35028
rect 18234 35048 18290 35057
rect 18234 34983 18290 34992
rect 17868 34944 17920 34950
rect 17868 34886 17920 34892
rect 17880 33658 17908 34886
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 18236 34604 18288 34610
rect 18236 34546 18288 34552
rect 18248 34241 18276 34546
rect 18234 34232 18290 34241
rect 18234 34167 18290 34176
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 17776 33448 17828 33454
rect 17776 33390 17828 33396
rect 17868 33312 17920 33318
rect 17868 33254 17920 33260
rect 17500 32768 17552 32774
rect 17500 32710 17552 32716
rect 17684 32496 17736 32502
rect 17684 32438 17736 32444
rect 17696 32366 17724 32438
rect 17500 32360 17552 32366
rect 17500 32302 17552 32308
rect 17684 32360 17736 32366
rect 17684 32302 17736 32308
rect 17512 32026 17540 32302
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17144 31334 17264 31362
rect 17132 30184 17184 30190
rect 17132 30126 17184 30132
rect 17144 29714 17172 30126
rect 17132 29708 17184 29714
rect 17132 29650 17184 29656
rect 17144 28626 17172 29650
rect 17236 29102 17264 31334
rect 17408 31272 17460 31278
rect 17408 31214 17460 31220
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 17420 28966 17448 31214
rect 17408 28960 17460 28966
rect 17408 28902 17460 28908
rect 17420 28626 17448 28902
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 17408 28620 17460 28626
rect 17408 28562 17460 28568
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17328 28082 17356 28358
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 17328 11354 17356 28018
rect 17512 12102 17540 31962
rect 17880 31210 17908 33254
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18064 32026 18092 32302
rect 18052 32020 18104 32026
rect 18052 31962 18104 31968
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17868 31204 17920 31210
rect 17868 31146 17920 31152
rect 17880 30802 17908 31146
rect 17868 30796 17920 30802
rect 17868 30738 17920 30744
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17592 29096 17644 29102
rect 17592 29038 17644 29044
rect 17684 29096 17736 29102
rect 17684 29038 17736 29044
rect 17604 28762 17632 29038
rect 17696 28966 17724 29038
rect 17684 28960 17736 28966
rect 17684 28902 17736 28908
rect 17592 28756 17644 28762
rect 17592 28698 17644 28704
rect 17604 27538 17632 28698
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17592 27532 17644 27538
rect 17592 27474 17644 27480
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 16658 18368 35090
rect 18420 34944 18472 34950
rect 18420 34886 18472 34892
rect 18432 33522 18460 34886
rect 18616 33590 18644 38218
rect 18708 36281 18736 39306
rect 18800 37233 18828 39494
rect 18984 38554 19012 39879
rect 19076 39545 19104 44678
rect 19168 41414 19196 47126
rect 19260 46170 19288 50866
rect 19444 50522 19472 52430
rect 19432 50516 19484 50522
rect 19432 50458 19484 50464
rect 22112 49978 22140 53654
rect 22204 53582 22232 56200
rect 22848 54194 22876 56200
rect 23492 54194 23520 56200
rect 24136 54194 24164 56200
rect 24780 54194 24808 56200
rect 25424 54194 25452 56200
rect 26068 54210 26096 56200
rect 26068 54194 26280 54210
rect 26712 54194 26740 56200
rect 27356 55214 27384 56200
rect 28000 56114 28028 56200
rect 28092 56114 28120 56222
rect 28000 56086 28120 56114
rect 27356 55186 27476 55214
rect 27448 54194 27476 55186
rect 27950 54428 28258 54437
rect 27950 54426 27956 54428
rect 28012 54426 28036 54428
rect 28092 54426 28116 54428
rect 28172 54426 28196 54428
rect 28252 54426 28258 54428
rect 28012 54374 28014 54426
rect 28194 54374 28196 54426
rect 27950 54372 27956 54374
rect 28012 54372 28036 54374
rect 28092 54372 28116 54374
rect 28172 54372 28196 54374
rect 28252 54372 28258 54374
rect 27950 54363 28258 54372
rect 28264 54256 28316 54262
rect 28264 54198 28316 54204
rect 22836 54188 22888 54194
rect 22836 54130 22888 54136
rect 23480 54188 23532 54194
rect 23480 54130 23532 54136
rect 24124 54188 24176 54194
rect 24124 54130 24176 54136
rect 24768 54188 24820 54194
rect 24768 54130 24820 54136
rect 25412 54188 25464 54194
rect 26068 54188 26292 54194
rect 26068 54182 26240 54188
rect 25412 54130 25464 54136
rect 26240 54130 26292 54136
rect 26700 54188 26752 54194
rect 26700 54130 26752 54136
rect 27436 54188 27488 54194
rect 27436 54130 27488 54136
rect 23572 54120 23624 54126
rect 23572 54062 23624 54068
rect 27712 54120 27764 54126
rect 27712 54062 27764 54068
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 22192 53576 22244 53582
rect 22192 53518 22244 53524
rect 22652 53440 22704 53446
rect 22652 53382 22704 53388
rect 23388 53440 23440 53446
rect 23388 53382 23440 53388
rect 22664 52698 22692 53382
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22652 52692 22704 52698
rect 22652 52634 22704 52640
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22468 50176 22520 50182
rect 22468 50118 22520 50124
rect 22100 49972 22152 49978
rect 22100 49914 22152 49920
rect 21916 49836 21968 49842
rect 21916 49778 21968 49784
rect 20996 48612 21048 48618
rect 20996 48554 21048 48560
rect 19800 48000 19852 48006
rect 19800 47942 19852 47948
rect 19524 47728 19576 47734
rect 19524 47670 19576 47676
rect 19248 46164 19300 46170
rect 19248 46106 19300 46112
rect 19536 44946 19564 47670
rect 19708 47592 19760 47598
rect 19708 47534 19760 47540
rect 19720 46510 19748 47534
rect 19708 46504 19760 46510
rect 19708 46446 19760 46452
rect 19720 45966 19748 46446
rect 19616 45960 19668 45966
rect 19616 45902 19668 45908
rect 19708 45960 19760 45966
rect 19708 45902 19760 45908
rect 19524 44940 19576 44946
rect 19524 44882 19576 44888
rect 19340 44328 19392 44334
rect 19340 44270 19392 44276
rect 19248 43920 19300 43926
rect 19248 43862 19300 43868
rect 19260 42226 19288 43862
rect 19352 43858 19380 44270
rect 19340 43852 19392 43858
rect 19340 43794 19392 43800
rect 19340 43716 19392 43722
rect 19340 43658 19392 43664
rect 19248 42220 19300 42226
rect 19248 42162 19300 42168
rect 19168 41386 19288 41414
rect 19260 40526 19288 41386
rect 19248 40520 19300 40526
rect 19154 40488 19210 40497
rect 19248 40462 19300 40468
rect 19154 40423 19210 40432
rect 19062 39536 19118 39545
rect 19062 39471 19118 39480
rect 18972 38548 19024 38554
rect 18972 38490 19024 38496
rect 18880 38412 18932 38418
rect 18880 38354 18932 38360
rect 18892 37398 18920 38354
rect 18880 37392 18932 37398
rect 18880 37334 18932 37340
rect 18786 37224 18842 37233
rect 18786 37159 18842 37168
rect 18788 37120 18840 37126
rect 18788 37062 18840 37068
rect 18694 36272 18750 36281
rect 18694 36207 18750 36216
rect 18800 35442 18828 37062
rect 19064 36916 19116 36922
rect 18892 36876 19064 36904
rect 18892 36825 18920 36876
rect 19064 36858 19116 36864
rect 18878 36816 18934 36825
rect 18878 36751 18934 36760
rect 19062 36816 19118 36825
rect 19062 36751 19118 36760
rect 18880 36236 18932 36242
rect 18880 36178 18932 36184
rect 18708 35414 18828 35442
rect 18708 34921 18736 35414
rect 18788 35284 18840 35290
rect 18788 35226 18840 35232
rect 18694 34912 18750 34921
rect 18694 34847 18750 34856
rect 18604 33584 18656 33590
rect 18604 33526 18656 33532
rect 18420 33516 18472 33522
rect 18420 33458 18472 33464
rect 18420 33108 18472 33114
rect 18420 33050 18472 33056
rect 18432 27606 18460 33050
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18420 27600 18472 27606
rect 18420 27542 18472 27548
rect 18524 27418 18552 31078
rect 18616 30258 18644 33526
rect 18708 33114 18736 34847
rect 18800 33998 18828 35226
rect 18892 34406 18920 36178
rect 19076 36174 19104 36751
rect 19064 36168 19116 36174
rect 19064 36110 19116 36116
rect 19168 36106 19196 40423
rect 19352 39030 19380 43658
rect 19524 43648 19576 43654
rect 19524 43590 19576 43596
rect 19432 42764 19484 42770
rect 19432 42706 19484 42712
rect 19444 41206 19472 42706
rect 19536 42702 19564 43590
rect 19524 42696 19576 42702
rect 19524 42638 19576 42644
rect 19628 41414 19656 45902
rect 19720 45490 19748 45902
rect 19708 45484 19760 45490
rect 19708 45426 19760 45432
rect 19812 45082 19840 47942
rect 20904 47116 20956 47122
rect 20904 47058 20956 47064
rect 20720 46980 20772 46986
rect 20720 46922 20772 46928
rect 20732 45422 20760 46922
rect 20812 45620 20864 45626
rect 20812 45562 20864 45568
rect 19984 45416 20036 45422
rect 19984 45358 20036 45364
rect 20720 45416 20772 45422
rect 20720 45358 20772 45364
rect 19800 45076 19852 45082
rect 19800 45018 19852 45024
rect 19996 44962 20024 45358
rect 20444 45280 20496 45286
rect 20444 45222 20496 45228
rect 19996 44946 20208 44962
rect 19996 44940 20220 44946
rect 19996 44934 20168 44940
rect 19708 44872 19760 44878
rect 19708 44814 19760 44820
rect 19720 44198 19748 44814
rect 19892 44736 19944 44742
rect 19892 44678 19944 44684
rect 19708 44192 19760 44198
rect 19708 44134 19760 44140
rect 19720 43314 19748 44134
rect 19904 43738 19932 44678
rect 19996 43994 20024 44934
rect 20168 44882 20220 44888
rect 20168 44804 20220 44810
rect 20168 44746 20220 44752
rect 20076 44532 20128 44538
rect 20076 44474 20128 44480
rect 20088 44266 20116 44474
rect 20076 44260 20128 44266
rect 20076 44202 20128 44208
rect 20180 44198 20208 44746
rect 20456 44470 20484 45222
rect 20444 44464 20496 44470
rect 20444 44406 20496 44412
rect 20168 44192 20220 44198
rect 20168 44134 20220 44140
rect 20260 44192 20312 44198
rect 20260 44134 20312 44140
rect 19984 43988 20036 43994
rect 19984 43930 20036 43936
rect 20076 43988 20128 43994
rect 20076 43930 20128 43936
rect 19812 43710 19932 43738
rect 19708 43308 19760 43314
rect 19708 43250 19760 43256
rect 19720 42770 19748 43250
rect 19708 42764 19760 42770
rect 19708 42706 19760 42712
rect 19628 41386 19748 41414
rect 19432 41200 19484 41206
rect 19432 41142 19484 41148
rect 19524 40112 19576 40118
rect 19524 40054 19576 40060
rect 19432 40044 19484 40050
rect 19432 39986 19484 39992
rect 19340 39024 19392 39030
rect 19340 38966 19392 38972
rect 19444 38350 19472 39986
rect 19536 38962 19564 40054
rect 19616 39976 19668 39982
rect 19616 39918 19668 39924
rect 19628 38962 19656 39918
rect 19524 38956 19576 38962
rect 19524 38898 19576 38904
rect 19616 38956 19668 38962
rect 19616 38898 19668 38904
rect 19720 38593 19748 41386
rect 19706 38584 19762 38593
rect 19706 38519 19762 38528
rect 19432 38344 19484 38350
rect 19432 38286 19484 38292
rect 19444 38185 19472 38286
rect 19430 38176 19486 38185
rect 19430 38111 19486 38120
rect 19340 37800 19392 37806
rect 19340 37742 19392 37748
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19524 37800 19576 37806
rect 19524 37742 19576 37748
rect 19248 37324 19300 37330
rect 19248 37266 19300 37272
rect 19260 36718 19288 37266
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 19248 36576 19300 36582
rect 19246 36544 19248 36553
rect 19300 36544 19302 36553
rect 19246 36479 19302 36488
rect 19352 36378 19380 37742
rect 19340 36372 19392 36378
rect 19340 36314 19392 36320
rect 19156 36100 19208 36106
rect 19156 36042 19208 36048
rect 19156 35828 19208 35834
rect 19156 35770 19208 35776
rect 19064 35624 19116 35630
rect 19064 35566 19116 35572
rect 19076 34610 19104 35566
rect 19064 34604 19116 34610
rect 19064 34546 19116 34552
rect 18880 34400 18932 34406
rect 18880 34342 18932 34348
rect 18788 33992 18840 33998
rect 18788 33934 18840 33940
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18800 33590 18828 33798
rect 18788 33584 18840 33590
rect 18788 33526 18840 33532
rect 18788 33448 18840 33454
rect 18788 33390 18840 33396
rect 18696 33108 18748 33114
rect 18696 33050 18748 33056
rect 18800 32026 18828 33390
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18800 30734 18828 31962
rect 18788 30728 18840 30734
rect 18788 30670 18840 30676
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18800 29730 18828 30670
rect 18708 29702 18828 29730
rect 18892 29714 18920 34342
rect 18970 34232 19026 34241
rect 19076 34202 19104 34546
rect 18970 34167 19026 34176
rect 19064 34196 19116 34202
rect 18984 33114 19012 34167
rect 19064 34138 19116 34144
rect 19064 33584 19116 33590
rect 19064 33526 19116 33532
rect 18972 33108 19024 33114
rect 18972 33050 19024 33056
rect 19076 32434 19104 33526
rect 19064 32428 19116 32434
rect 19064 32370 19116 32376
rect 19064 32292 19116 32298
rect 19064 32234 19116 32240
rect 19076 31958 19104 32234
rect 19064 31952 19116 31958
rect 19064 31894 19116 31900
rect 19064 31748 19116 31754
rect 19064 31690 19116 31696
rect 19076 31414 19104 31690
rect 19064 31408 19116 31414
rect 19064 31350 19116 31356
rect 19076 30870 19104 31350
rect 19064 30864 19116 30870
rect 19064 30806 19116 30812
rect 18972 30592 19024 30598
rect 18972 30534 19024 30540
rect 18880 29708 18932 29714
rect 18604 29096 18656 29102
rect 18604 29038 18656 29044
rect 18616 27538 18644 29038
rect 18708 28762 18736 29702
rect 18880 29650 18932 29656
rect 18788 29504 18840 29510
rect 18788 29446 18840 29452
rect 18800 28762 18828 29446
rect 18696 28756 18748 28762
rect 18696 28698 18748 28704
rect 18788 28756 18840 28762
rect 18788 28698 18840 28704
rect 18604 27532 18656 27538
rect 18604 27474 18656 27480
rect 18524 27390 18644 27418
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18432 26382 18460 27270
rect 18616 26450 18644 27390
rect 18800 26450 18828 28698
rect 18892 28082 18920 29650
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18880 27940 18932 27946
rect 18880 27882 18932 27888
rect 18604 26444 18656 26450
rect 18604 26386 18656 26392
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18892 22094 18920 27882
rect 18984 27470 19012 30534
rect 19076 29578 19104 30806
rect 19064 29572 19116 29578
rect 19064 29514 19116 29520
rect 19076 29238 19104 29514
rect 19064 29232 19116 29238
rect 19064 29174 19116 29180
rect 19076 28490 19104 29174
rect 19064 28484 19116 28490
rect 19064 28426 19116 28432
rect 19168 28218 19196 35770
rect 19352 35766 19380 36314
rect 19340 35760 19392 35766
rect 19340 35702 19392 35708
rect 19340 34536 19392 34542
rect 19340 34478 19392 34484
rect 19248 34196 19300 34202
rect 19248 34138 19300 34144
rect 19260 33590 19288 34138
rect 19248 33584 19300 33590
rect 19248 33526 19300 33532
rect 19248 33380 19300 33386
rect 19248 33322 19300 33328
rect 19260 31890 19288 33322
rect 19352 32774 19380 34478
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19248 31884 19300 31890
rect 19248 31826 19300 31832
rect 19352 30870 19380 32710
rect 19444 32026 19472 37742
rect 19536 34406 19564 37742
rect 19812 37126 19840 43710
rect 19892 43648 19944 43654
rect 19892 43590 19944 43596
rect 19904 40730 19932 43590
rect 20088 43382 20116 43930
rect 20076 43376 20128 43382
rect 20076 43318 20128 43324
rect 19984 42696 20036 42702
rect 19984 42638 20036 42644
rect 19892 40724 19944 40730
rect 19892 40666 19944 40672
rect 19996 39284 20024 42638
rect 20088 40633 20116 43318
rect 20180 42838 20208 44134
rect 20272 43450 20300 44134
rect 20720 43648 20772 43654
rect 20720 43590 20772 43596
rect 20260 43444 20312 43450
rect 20260 43386 20312 43392
rect 20628 43240 20680 43246
rect 20628 43182 20680 43188
rect 20168 42832 20220 42838
rect 20168 42774 20220 42780
rect 20536 42764 20588 42770
rect 20536 42706 20588 42712
rect 20548 42226 20576 42706
rect 20640 42634 20668 43182
rect 20628 42628 20680 42634
rect 20628 42570 20680 42576
rect 20352 42220 20404 42226
rect 20352 42162 20404 42168
rect 20536 42220 20588 42226
rect 20536 42162 20588 42168
rect 20364 41585 20392 42162
rect 20444 42084 20496 42090
rect 20444 42026 20496 42032
rect 20350 41576 20406 41585
rect 20350 41511 20406 41520
rect 20074 40624 20130 40633
rect 20074 40559 20076 40568
rect 20128 40559 20130 40568
rect 20076 40530 20128 40536
rect 19904 39256 20024 39284
rect 20168 39296 20220 39302
rect 19904 37194 19932 39256
rect 20168 39238 20220 39244
rect 20180 38554 20208 39238
rect 20168 38548 20220 38554
rect 20168 38490 20220 38496
rect 20076 38480 20128 38486
rect 19982 38448 20038 38457
rect 20076 38422 20128 38428
rect 19982 38383 20038 38392
rect 19996 38350 20024 38383
rect 19984 38344 20036 38350
rect 20088 38321 20116 38422
rect 19984 38286 20036 38292
rect 20074 38312 20130 38321
rect 20074 38247 20130 38256
rect 20076 37732 20128 37738
rect 20076 37674 20128 37680
rect 19892 37188 19944 37194
rect 19892 37130 19944 37136
rect 19800 37120 19852 37126
rect 19800 37062 19852 37068
rect 19616 36916 19668 36922
rect 19616 36858 19668 36864
rect 19628 36145 19656 36858
rect 19800 36712 19852 36718
rect 19800 36654 19852 36660
rect 19614 36136 19670 36145
rect 19614 36071 19670 36080
rect 19708 36100 19760 36106
rect 19708 36042 19760 36048
rect 19616 35148 19668 35154
rect 19616 35090 19668 35096
rect 19524 34400 19576 34406
rect 19524 34342 19576 34348
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19628 31822 19656 35090
rect 19720 34542 19748 36042
rect 19812 35601 19840 36654
rect 19798 35592 19854 35601
rect 19798 35527 19854 35536
rect 19708 34536 19760 34542
rect 19708 34478 19760 34484
rect 19812 32502 19840 35527
rect 19892 34944 19944 34950
rect 19892 34886 19944 34892
rect 19800 32496 19852 32502
rect 19800 32438 19852 32444
rect 19708 32224 19760 32230
rect 19708 32166 19760 32172
rect 19616 31816 19668 31822
rect 19616 31758 19668 31764
rect 19524 31680 19576 31686
rect 19524 31622 19576 31628
rect 19536 31210 19564 31622
rect 19524 31204 19576 31210
rect 19524 31146 19576 31152
rect 19340 30864 19392 30870
rect 19340 30806 19392 30812
rect 19524 30252 19576 30258
rect 19524 30194 19576 30200
rect 19536 29850 19564 30194
rect 19524 29844 19576 29850
rect 19524 29786 19576 29792
rect 19248 28688 19300 28694
rect 19248 28630 19300 28636
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 19260 27946 19288 28630
rect 19536 28558 19564 29786
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19720 28014 19748 32166
rect 19904 31754 19932 34886
rect 20088 33046 20116 37674
rect 20258 36952 20314 36961
rect 20258 36887 20314 36896
rect 20168 33924 20220 33930
rect 20168 33866 20220 33872
rect 20076 33040 20128 33046
rect 20076 32982 20128 32988
rect 20076 32836 20128 32842
rect 20076 32778 20128 32784
rect 20088 32502 20116 32778
rect 20076 32496 20128 32502
rect 20076 32438 20128 32444
rect 20088 31754 20116 32438
rect 20180 31754 20208 33866
rect 20272 32570 20300 36887
rect 20364 35086 20392 41511
rect 20456 41206 20484 42026
rect 20444 41200 20496 41206
rect 20444 41142 20496 41148
rect 20442 40624 20498 40633
rect 20548 40594 20576 42162
rect 20640 41682 20668 42570
rect 20628 41676 20680 41682
rect 20628 41618 20680 41624
rect 20628 40928 20680 40934
rect 20628 40870 20680 40876
rect 20442 40559 20498 40568
rect 20536 40588 20588 40594
rect 20456 37806 20484 40559
rect 20536 40530 20588 40536
rect 20640 40186 20668 40870
rect 20628 40180 20680 40186
rect 20628 40122 20680 40128
rect 20732 38010 20760 43590
rect 20824 42106 20852 45562
rect 20916 45370 20944 47058
rect 21008 46034 21036 48554
rect 21456 48204 21508 48210
rect 21456 48146 21508 48152
rect 21468 47802 21496 48146
rect 21456 47796 21508 47802
rect 21456 47738 21508 47744
rect 21088 47660 21140 47666
rect 21088 47602 21140 47608
rect 21100 46578 21128 47602
rect 21272 47456 21324 47462
rect 21272 47398 21324 47404
rect 21284 47054 21312 47398
rect 21468 47122 21496 47738
rect 21456 47116 21508 47122
rect 21456 47058 21508 47064
rect 21272 47048 21324 47054
rect 21272 46990 21324 46996
rect 21180 46912 21232 46918
rect 21180 46854 21232 46860
rect 21088 46572 21140 46578
rect 21088 46514 21140 46520
rect 20996 46028 21048 46034
rect 20996 45970 21048 45976
rect 21100 45490 21128 46514
rect 21192 46510 21220 46854
rect 21640 46640 21692 46646
rect 21640 46582 21692 46588
rect 21180 46504 21232 46510
rect 21180 46446 21232 46452
rect 21088 45484 21140 45490
rect 21088 45426 21140 45432
rect 20916 45354 21036 45370
rect 20916 45348 21048 45354
rect 20916 45342 20996 45348
rect 20996 45290 21048 45296
rect 21100 44792 21128 45426
rect 21192 45370 21220 46446
rect 21652 46374 21680 46582
rect 21640 46368 21692 46374
rect 21640 46310 21692 46316
rect 21364 46028 21416 46034
rect 21364 45970 21416 45976
rect 21192 45342 21312 45370
rect 21180 44804 21232 44810
rect 21100 44764 21180 44792
rect 21100 44402 21128 44764
rect 21180 44746 21232 44752
rect 21088 44396 21140 44402
rect 21088 44338 21140 44344
rect 21100 43314 21128 44338
rect 21284 44334 21312 45342
rect 21272 44328 21324 44334
rect 21272 44270 21324 44276
rect 21376 43858 21404 45970
rect 21548 45348 21600 45354
rect 21548 45290 21600 45296
rect 21456 44872 21508 44878
rect 21456 44814 21508 44820
rect 21468 44538 21496 44814
rect 21456 44532 21508 44538
rect 21456 44474 21508 44480
rect 21560 44266 21588 45290
rect 21548 44260 21600 44266
rect 21548 44202 21600 44208
rect 21364 43852 21416 43858
rect 21364 43794 21416 43800
rect 21272 43648 21324 43654
rect 21272 43590 21324 43596
rect 21088 43308 21140 43314
rect 21088 43250 21140 43256
rect 21100 42634 21128 43250
rect 21088 42628 21140 42634
rect 21088 42570 21140 42576
rect 20824 42078 20944 42106
rect 21100 42090 21128 42570
rect 20812 42016 20864 42022
rect 20812 41958 20864 41964
rect 20824 40458 20852 41958
rect 20916 41449 20944 42078
rect 21088 42084 21140 42090
rect 21088 42026 21140 42032
rect 21180 41744 21232 41750
rect 21180 41686 21232 41692
rect 21088 41608 21140 41614
rect 21088 41550 21140 41556
rect 20996 41472 21048 41478
rect 20902 41440 20958 41449
rect 20996 41414 21048 41420
rect 20902 41375 20958 41384
rect 21008 41002 21036 41414
rect 21100 41138 21128 41550
rect 21192 41528 21220 41686
rect 21284 41682 21312 43590
rect 21376 43450 21404 43794
rect 21364 43444 21416 43450
rect 21364 43386 21416 43392
rect 21652 43110 21680 46310
rect 21732 46164 21784 46170
rect 21732 46106 21784 46112
rect 21744 44742 21772 46106
rect 21824 45076 21876 45082
rect 21824 45018 21876 45024
rect 21836 44810 21864 45018
rect 21824 44804 21876 44810
rect 21824 44746 21876 44752
rect 21732 44736 21784 44742
rect 21732 44678 21784 44684
rect 21640 43104 21692 43110
rect 21640 43046 21692 43052
rect 21640 42900 21692 42906
rect 21640 42842 21692 42848
rect 21548 42560 21600 42566
rect 21548 42502 21600 42508
rect 21560 42090 21588 42502
rect 21548 42084 21600 42090
rect 21548 42026 21600 42032
rect 21652 41818 21680 42842
rect 21640 41812 21692 41818
rect 21640 41754 21692 41760
rect 21272 41676 21324 41682
rect 21272 41618 21324 41624
rect 21192 41500 21496 41528
rect 21178 41440 21234 41449
rect 21178 41375 21234 41384
rect 21192 41290 21220 41375
rect 21192 41262 21312 41290
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 20996 40996 21048 41002
rect 20996 40938 21048 40944
rect 20904 40928 20956 40934
rect 20904 40870 20956 40876
rect 20916 40730 20944 40870
rect 20904 40724 20956 40730
rect 20904 40666 20956 40672
rect 20996 40724 21048 40730
rect 20996 40666 21048 40672
rect 20812 40452 20864 40458
rect 20812 40394 20864 40400
rect 20904 40452 20956 40458
rect 20904 40394 20956 40400
rect 20812 40180 20864 40186
rect 20812 40122 20864 40128
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 20444 37800 20496 37806
rect 20444 37742 20496 37748
rect 20824 36854 20852 40122
rect 20916 39506 20944 40394
rect 21008 40390 21036 40666
rect 20996 40384 21048 40390
rect 20996 40326 21048 40332
rect 20996 40044 21048 40050
rect 20996 39986 21048 39992
rect 20904 39500 20956 39506
rect 20904 39442 20956 39448
rect 20904 39296 20956 39302
rect 20904 39238 20956 39244
rect 20916 38214 20944 39238
rect 21008 39030 21036 39986
rect 20996 39024 21048 39030
rect 20996 38966 21048 38972
rect 21088 38752 21140 38758
rect 21088 38694 21140 38700
rect 20904 38208 20956 38214
rect 20904 38150 20956 38156
rect 20996 37868 21048 37874
rect 20996 37810 21048 37816
rect 21008 37466 21036 37810
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 20812 36848 20864 36854
rect 20812 36790 20864 36796
rect 20902 36680 20958 36689
rect 20902 36615 20958 36624
rect 20720 36304 20772 36310
rect 20720 36246 20772 36252
rect 20444 36236 20496 36242
rect 20444 36178 20496 36184
rect 20456 35154 20484 36178
rect 20732 35834 20760 36246
rect 20812 36168 20864 36174
rect 20812 36110 20864 36116
rect 20720 35828 20772 35834
rect 20720 35770 20772 35776
rect 20824 35766 20852 36110
rect 20812 35760 20864 35766
rect 20812 35702 20864 35708
rect 20444 35148 20496 35154
rect 20444 35090 20496 35096
rect 20352 35080 20404 35086
rect 20352 35022 20404 35028
rect 20824 35018 20852 35702
rect 20536 35012 20588 35018
rect 20812 35012 20864 35018
rect 20536 34954 20588 34960
rect 20732 34972 20812 35000
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20456 32774 20484 34886
rect 20548 33658 20576 34954
rect 20732 34678 20760 34972
rect 20812 34954 20864 34960
rect 20720 34672 20772 34678
rect 20720 34614 20772 34620
rect 20628 34536 20680 34542
rect 20628 34478 20680 34484
rect 20536 33652 20588 33658
rect 20536 33594 20588 33600
rect 20640 32978 20668 34478
rect 20732 33930 20760 34614
rect 20720 33924 20772 33930
rect 20720 33866 20772 33872
rect 20628 32972 20680 32978
rect 20628 32914 20680 32920
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20444 32768 20496 32774
rect 20444 32710 20496 32716
rect 20260 32564 20312 32570
rect 20260 32506 20312 32512
rect 19904 31726 20024 31754
rect 19800 31680 19852 31686
rect 19800 31622 19852 31628
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 19248 27940 19300 27946
rect 19248 27882 19300 27888
rect 19156 27600 19208 27606
rect 19156 27542 19208 27548
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18892 22066 19012 22094
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18984 15910 19012 22066
rect 19168 21894 19196 27542
rect 19812 27062 19840 31622
rect 19892 30320 19944 30326
rect 19892 30262 19944 30268
rect 19904 29646 19932 30262
rect 19892 29640 19944 29646
rect 19892 29582 19944 29588
rect 19904 29238 19932 29582
rect 19892 29232 19944 29238
rect 19892 29174 19944 29180
rect 19996 29050 20024 31726
rect 20076 31748 20128 31754
rect 20076 31690 20128 31696
rect 20168 31748 20220 31754
rect 20168 31690 20220 31696
rect 20548 31226 20576 32846
rect 20732 32842 20760 33866
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20628 32768 20680 32774
rect 20628 32710 20680 32716
rect 20180 31198 20576 31226
rect 20180 30870 20208 31198
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20168 30864 20220 30870
rect 20168 30806 20220 30812
rect 19904 29022 20024 29050
rect 19904 28762 19932 29022
rect 19892 28756 19944 28762
rect 19892 28698 19944 28704
rect 19800 27056 19852 27062
rect 19800 26998 19852 27004
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19904 21350 19932 28698
rect 20180 28422 20208 30806
rect 20352 30184 20404 30190
rect 20352 30126 20404 30132
rect 20260 29232 20312 29238
rect 20260 29174 20312 29180
rect 20272 28490 20300 29174
rect 20260 28484 20312 28490
rect 20260 28426 20312 28432
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18432 12850 18460 13262
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17328 6914 17356 11290
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18420 7268 18472 7274
rect 18420 7210 18472 7216
rect 17236 6886 17356 6914
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 17236 5574 17264 6886
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18432 5302 18460 7210
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 18616 4622 18644 11630
rect 18984 10470 19012 15846
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 19536 6798 19564 13126
rect 19996 11762 20024 19450
rect 20088 12782 20116 28018
rect 20168 26512 20220 26518
rect 20168 26454 20220 26460
rect 20180 18766 20208 26454
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20088 7206 20116 12718
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20180 11694 20208 12174
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20272 9586 20300 28426
rect 20364 28014 20392 30126
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20456 27606 20484 31078
rect 20640 30648 20668 32710
rect 20720 32224 20772 32230
rect 20720 32166 20772 32172
rect 20732 31958 20760 32166
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 20732 31793 20760 31894
rect 20812 31816 20864 31822
rect 20718 31784 20774 31793
rect 20812 31758 20864 31764
rect 20718 31719 20774 31728
rect 20732 30802 20760 31719
rect 20824 31482 20852 31758
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 20916 31414 20944 36615
rect 21100 33658 21128 38694
rect 21284 38554 21312 41262
rect 21364 41200 21416 41206
rect 21364 41142 21416 41148
rect 21376 40458 21404 41142
rect 21364 40452 21416 40458
rect 21364 40394 21416 40400
rect 21376 40050 21404 40394
rect 21364 40044 21416 40050
rect 21364 39986 21416 39992
rect 21376 39030 21404 39986
rect 21468 39658 21496 41500
rect 21744 40050 21772 44678
rect 21928 43217 21956 49778
rect 22100 48136 22152 48142
rect 22100 48078 22152 48084
rect 22008 48000 22060 48006
rect 22008 47942 22060 47948
rect 22020 47802 22048 47942
rect 22008 47796 22060 47802
rect 22008 47738 22060 47744
rect 22112 47530 22140 48078
rect 22192 47796 22244 47802
rect 22192 47738 22244 47744
rect 22100 47524 22152 47530
rect 22100 47466 22152 47472
rect 22112 47054 22140 47466
rect 22204 47190 22232 47738
rect 22480 47734 22508 50118
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22744 49156 22796 49162
rect 22744 49098 22796 49104
rect 22560 48068 22612 48074
rect 22560 48010 22612 48016
rect 22468 47728 22520 47734
rect 22468 47670 22520 47676
rect 22192 47184 22244 47190
rect 22192 47126 22244 47132
rect 22100 47048 22152 47054
rect 22100 46990 22152 46996
rect 22008 46980 22060 46986
rect 22008 46922 22060 46928
rect 22020 44538 22048 46922
rect 22112 46374 22140 46990
rect 22572 46714 22600 48010
rect 22652 48000 22704 48006
rect 22652 47942 22704 47948
rect 22664 47598 22692 47942
rect 22652 47592 22704 47598
rect 22652 47534 22704 47540
rect 22560 46708 22612 46714
rect 22560 46650 22612 46656
rect 22100 46368 22152 46374
rect 22100 46310 22152 46316
rect 22112 46034 22140 46310
rect 22100 46028 22152 46034
rect 22100 45970 22152 45976
rect 22192 45280 22244 45286
rect 22192 45222 22244 45228
rect 22008 44532 22060 44538
rect 22008 44474 22060 44480
rect 21914 43208 21970 43217
rect 21914 43143 21970 43152
rect 21824 42696 21876 42702
rect 21824 42638 21876 42644
rect 21836 42294 21864 42638
rect 21916 42560 21968 42566
rect 21916 42502 21968 42508
rect 21824 42288 21876 42294
rect 21824 42230 21876 42236
rect 21928 42158 21956 42502
rect 21916 42152 21968 42158
rect 21916 42094 21968 42100
rect 21824 42084 21876 42090
rect 21824 42026 21876 42032
rect 21836 41414 21864 42026
rect 21928 41818 21956 42094
rect 21916 41812 21968 41818
rect 21916 41754 21968 41760
rect 22008 41540 22060 41546
rect 22008 41482 22060 41488
rect 21836 41386 21956 41414
rect 21824 40180 21876 40186
rect 21824 40122 21876 40128
rect 21732 40044 21784 40050
rect 21732 39986 21784 39992
rect 21468 39642 21772 39658
rect 21468 39636 21784 39642
rect 21468 39630 21732 39636
rect 21548 39568 21600 39574
rect 21548 39510 21600 39516
rect 21456 39500 21508 39506
rect 21456 39442 21508 39448
rect 21468 39098 21496 39442
rect 21560 39098 21588 39510
rect 21456 39092 21508 39098
rect 21456 39034 21508 39040
rect 21548 39092 21600 39098
rect 21548 39034 21600 39040
rect 21364 39024 21416 39030
rect 21364 38966 21416 38972
rect 21456 38956 21508 38962
rect 21456 38898 21508 38904
rect 21272 38548 21324 38554
rect 21272 38490 21324 38496
rect 21468 38282 21496 38898
rect 21560 38894 21588 39034
rect 21548 38888 21600 38894
rect 21548 38830 21600 38836
rect 21456 38276 21508 38282
rect 21456 38218 21508 38224
rect 21468 37874 21496 38218
rect 21652 38010 21680 39630
rect 21732 39578 21784 39584
rect 21836 38826 21864 40122
rect 21824 38820 21876 38826
rect 21824 38762 21876 38768
rect 21730 38584 21786 38593
rect 21730 38519 21786 38528
rect 21744 38350 21772 38519
rect 21836 38486 21864 38762
rect 21824 38480 21876 38486
rect 21824 38422 21876 38428
rect 21732 38344 21784 38350
rect 21732 38286 21784 38292
rect 21640 38004 21692 38010
rect 21640 37946 21692 37952
rect 21548 37936 21600 37942
rect 21548 37878 21600 37884
rect 21456 37868 21508 37874
rect 21456 37810 21508 37816
rect 21180 36712 21232 36718
rect 21180 36654 21232 36660
rect 21364 36712 21416 36718
rect 21364 36654 21416 36660
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21008 32570 21036 33458
rect 20996 32564 21048 32570
rect 20996 32506 21048 32512
rect 20904 31408 20956 31414
rect 20904 31350 20956 31356
rect 20904 31272 20956 31278
rect 20904 31214 20956 31220
rect 20916 31142 20944 31214
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20720 30796 20772 30802
rect 20720 30738 20772 30744
rect 20548 30620 20668 30648
rect 20548 29510 20576 30620
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20640 29578 20668 30262
rect 21008 30190 21036 32506
rect 21088 31748 21140 31754
rect 21088 31690 21140 31696
rect 21100 31278 21128 31690
rect 21088 31272 21140 31278
rect 21088 31214 21140 31220
rect 21192 30598 21220 36654
rect 21272 35488 21324 35494
rect 21272 35430 21324 35436
rect 21284 35154 21312 35430
rect 21272 35148 21324 35154
rect 21272 35090 21324 35096
rect 21376 33590 21404 36654
rect 21456 35488 21508 35494
rect 21456 35430 21508 35436
rect 21468 35290 21496 35430
rect 21456 35284 21508 35290
rect 21456 35226 21508 35232
rect 21456 34196 21508 34202
rect 21456 34138 21508 34144
rect 21272 33584 21324 33590
rect 21272 33526 21324 33532
rect 21364 33584 21416 33590
rect 21364 33526 21416 33532
rect 21284 31346 21312 33526
rect 21364 33448 21416 33454
rect 21364 33390 21416 33396
rect 21376 32910 21404 33390
rect 21468 33318 21496 34138
rect 21456 33312 21508 33318
rect 21456 33254 21508 33260
rect 21364 32904 21416 32910
rect 21364 32846 21416 32852
rect 21376 31890 21404 32846
rect 21560 32230 21588 37878
rect 21732 37120 21784 37126
rect 21732 37062 21784 37068
rect 21640 34400 21692 34406
rect 21640 34342 21692 34348
rect 21652 34202 21680 34342
rect 21640 34196 21692 34202
rect 21640 34138 21692 34144
rect 21640 33312 21692 33318
rect 21640 33254 21692 33260
rect 21548 32224 21600 32230
rect 21548 32166 21600 32172
rect 21456 31952 21508 31958
rect 21456 31894 21508 31900
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 21362 31784 21418 31793
rect 21362 31719 21418 31728
rect 21376 31686 21404 31719
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 21180 30592 21232 30598
rect 21180 30534 21232 30540
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 20628 29572 20680 29578
rect 20628 29514 20680 29520
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20640 29238 20668 29514
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20444 27600 20496 27606
rect 20444 27542 20496 27548
rect 20916 27130 20944 28358
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 21284 22094 21312 31282
rect 21468 30190 21496 31894
rect 21652 31890 21680 33254
rect 21744 32570 21772 37062
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 21732 32564 21784 32570
rect 21732 32506 21784 32512
rect 21640 31884 21692 31890
rect 21640 31826 21692 31832
rect 21640 31680 21692 31686
rect 21640 31622 21692 31628
rect 21652 31414 21680 31622
rect 21640 31408 21692 31414
rect 21640 31350 21692 31356
rect 21456 30184 21508 30190
rect 21456 30126 21508 30132
rect 21468 29866 21496 30126
rect 21468 29838 21588 29866
rect 21456 29708 21508 29714
rect 21456 29650 21508 29656
rect 21468 29306 21496 29650
rect 21456 29300 21508 29306
rect 21456 29242 21508 29248
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21376 28218 21404 28358
rect 21364 28212 21416 28218
rect 21364 28154 21416 28160
rect 21468 26926 21496 29242
rect 21560 28966 21588 29838
rect 21548 28960 21600 28966
rect 21548 28902 21600 28908
rect 21560 28626 21588 28902
rect 21548 28620 21600 28626
rect 21548 28562 21600 28568
rect 21652 28082 21680 31350
rect 21732 31136 21784 31142
rect 21732 31078 21784 31084
rect 21640 28076 21692 28082
rect 21640 28018 21692 28024
rect 21456 26920 21508 26926
rect 21456 26862 21508 26868
rect 21744 22094 21772 31078
rect 21836 29306 21864 36722
rect 21928 36582 21956 41386
rect 22020 41206 22048 41482
rect 22100 41268 22152 41274
rect 22100 41210 22152 41216
rect 22008 41200 22060 41206
rect 22008 41142 22060 41148
rect 22112 40662 22140 41210
rect 22100 40656 22152 40662
rect 22100 40598 22152 40604
rect 22008 37868 22060 37874
rect 22008 37810 22060 37816
rect 22020 36854 22048 37810
rect 22008 36848 22060 36854
rect 22008 36790 22060 36796
rect 21916 36576 21968 36582
rect 21916 36518 21968 36524
rect 22020 36242 22048 36790
rect 22008 36236 22060 36242
rect 22008 36178 22060 36184
rect 22112 35766 22140 40598
rect 22204 39982 22232 45222
rect 22374 44432 22430 44441
rect 22284 44396 22336 44402
rect 22374 44367 22430 44376
rect 22284 44338 22336 44344
rect 22296 40186 22324 44338
rect 22388 44334 22416 44367
rect 22376 44328 22428 44334
rect 22376 44270 22428 44276
rect 22388 41070 22416 44270
rect 22468 43852 22520 43858
rect 22468 43794 22520 43800
rect 22480 43382 22508 43794
rect 22468 43376 22520 43382
rect 22468 43318 22520 43324
rect 22468 43240 22520 43246
rect 22468 43182 22520 43188
rect 22480 41682 22508 43182
rect 22572 42922 22600 46650
rect 22652 46368 22704 46374
rect 22652 46310 22704 46316
rect 22664 43790 22692 46310
rect 22652 43784 22704 43790
rect 22652 43726 22704 43732
rect 22572 42894 22692 42922
rect 22560 42764 22612 42770
rect 22560 42706 22612 42712
rect 22572 42294 22600 42706
rect 22560 42288 22612 42294
rect 22560 42230 22612 42236
rect 22468 41676 22520 41682
rect 22468 41618 22520 41624
rect 22572 41546 22600 42230
rect 22560 41540 22612 41546
rect 22560 41482 22612 41488
rect 22376 41064 22428 41070
rect 22376 41006 22428 41012
rect 22388 40934 22416 41006
rect 22376 40928 22428 40934
rect 22376 40870 22428 40876
rect 22284 40180 22336 40186
rect 22284 40122 22336 40128
rect 22388 40066 22416 40870
rect 22558 40624 22614 40633
rect 22558 40559 22560 40568
rect 22612 40559 22614 40568
rect 22560 40530 22612 40536
rect 22468 40384 22520 40390
rect 22468 40326 22520 40332
rect 22480 40118 22508 40326
rect 22296 40038 22416 40066
rect 22468 40112 22520 40118
rect 22468 40054 22520 40060
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 22192 36916 22244 36922
rect 22192 36858 22244 36864
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 22204 35698 22232 36858
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22296 35578 22324 40038
rect 22560 39976 22612 39982
rect 22560 39918 22612 39924
rect 22468 39636 22520 39642
rect 22468 39578 22520 39584
rect 22480 39302 22508 39578
rect 22468 39296 22520 39302
rect 22468 39238 22520 39244
rect 22572 38298 22600 39918
rect 22664 39506 22692 42894
rect 22756 41478 22784 49098
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22836 47660 22888 47666
rect 22836 47602 22888 47608
rect 22848 47258 22876 47602
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22836 47252 22888 47258
rect 22836 47194 22888 47200
rect 22836 46504 22888 46510
rect 22836 46446 22888 46452
rect 22848 45422 22876 46446
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 23296 46028 23348 46034
rect 23296 45970 23348 45976
rect 22836 45416 22888 45422
rect 22836 45358 22888 45364
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 23308 44334 23336 45970
rect 23400 45914 23428 53382
rect 23584 53242 23612 54062
rect 25412 53984 25464 53990
rect 25412 53926 25464 53932
rect 26056 53984 26108 53990
rect 26056 53926 26108 53932
rect 27436 53984 27488 53990
rect 27436 53926 27488 53932
rect 23572 53236 23624 53242
rect 23572 53178 23624 53184
rect 24860 53168 24912 53174
rect 24860 53110 24912 53116
rect 24768 52556 24820 52562
rect 24768 52498 24820 52504
rect 23940 51264 23992 51270
rect 23940 51206 23992 51212
rect 23480 48680 23532 48686
rect 23480 48622 23532 48628
rect 23492 46918 23520 48622
rect 23572 47592 23624 47598
rect 23572 47534 23624 47540
rect 23480 46912 23532 46918
rect 23480 46854 23532 46860
rect 23492 46170 23520 46854
rect 23480 46164 23532 46170
rect 23480 46106 23532 46112
rect 23400 45886 23520 45914
rect 23492 45830 23520 45886
rect 23388 45824 23440 45830
rect 23388 45766 23440 45772
rect 23480 45824 23532 45830
rect 23480 45766 23532 45772
rect 23400 45286 23428 45766
rect 23388 45280 23440 45286
rect 23388 45222 23440 45228
rect 23584 44470 23612 47534
rect 23848 46980 23900 46986
rect 23848 46922 23900 46928
rect 23860 46646 23888 46922
rect 23848 46640 23900 46646
rect 23848 46582 23900 46588
rect 23860 45898 23888 46582
rect 23848 45892 23900 45898
rect 23848 45834 23900 45840
rect 23952 45558 23980 51206
rect 24492 50924 24544 50930
rect 24492 50866 24544 50872
rect 24308 46096 24360 46102
rect 24308 46038 24360 46044
rect 23756 45552 23808 45558
rect 23756 45494 23808 45500
rect 23940 45552 23992 45558
rect 23940 45494 23992 45500
rect 23664 44736 23716 44742
rect 23664 44678 23716 44684
rect 23572 44464 23624 44470
rect 23572 44406 23624 44412
rect 23296 44328 23348 44334
rect 23296 44270 23348 44276
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22836 43376 22888 43382
rect 22836 43318 22888 43324
rect 22848 42770 22876 43318
rect 23308 43246 23336 44270
rect 23388 44192 23440 44198
rect 23440 44140 23520 44146
rect 23388 44134 23520 44140
rect 23400 44118 23520 44134
rect 23388 43852 23440 43858
rect 23388 43794 23440 43800
rect 23296 43240 23348 43246
rect 23296 43182 23348 43188
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 23308 42770 23336 43182
rect 22836 42764 22888 42770
rect 22836 42706 22888 42712
rect 23296 42764 23348 42770
rect 23296 42706 23348 42712
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 23296 41676 23348 41682
rect 23400 41664 23428 43794
rect 23348 41636 23428 41664
rect 23296 41618 23348 41624
rect 22744 41472 22796 41478
rect 22744 41414 22796 41420
rect 23308 41002 23336 41618
rect 23296 40996 23348 41002
rect 23296 40938 23348 40944
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22834 40216 22890 40225
rect 22834 40151 22890 40160
rect 22848 40118 22876 40151
rect 22836 40112 22888 40118
rect 22836 40054 22888 40060
rect 22744 39840 22796 39846
rect 22744 39782 22796 39788
rect 22652 39500 22704 39506
rect 22652 39442 22704 39448
rect 22756 39370 22784 39782
rect 22848 39624 22876 40054
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22848 39596 22968 39624
rect 22744 39364 22796 39370
rect 22744 39306 22796 39312
rect 22652 39296 22704 39302
rect 22652 39238 22704 39244
rect 22480 38270 22600 38298
rect 22376 37324 22428 37330
rect 22376 37266 22428 37272
rect 22204 35550 22324 35578
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 22020 33998 22048 34478
rect 22100 34400 22152 34406
rect 22100 34342 22152 34348
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 22020 33454 22048 33934
rect 22112 33658 22140 34342
rect 22100 33652 22152 33658
rect 22100 33594 22152 33600
rect 22008 33448 22060 33454
rect 22008 33390 22060 33396
rect 22112 32842 22140 33594
rect 22204 33300 22232 35550
rect 22388 35290 22416 37266
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22388 34678 22416 35226
rect 22480 34950 22508 38270
rect 22560 38208 22612 38214
rect 22560 38150 22612 38156
rect 22572 38010 22600 38150
rect 22560 38004 22612 38010
rect 22560 37946 22612 37952
rect 22664 37890 22692 39238
rect 22744 39024 22796 39030
rect 22742 38992 22744 39001
rect 22796 38992 22798 39001
rect 22742 38927 22798 38936
rect 22940 38865 22968 39596
rect 23020 39568 23072 39574
rect 23018 39536 23020 39545
rect 23072 39536 23074 39545
rect 23018 39471 23074 39480
rect 23296 39364 23348 39370
rect 23296 39306 23348 39312
rect 22926 38856 22982 38865
rect 22926 38791 22982 38800
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22744 38412 22796 38418
rect 23308 38400 23336 39306
rect 23386 38992 23442 39001
rect 23386 38927 23442 38936
rect 22744 38354 22796 38360
rect 22848 38372 23336 38400
rect 22572 37862 22692 37890
rect 22572 36582 22600 37862
rect 22756 36718 22784 38354
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22744 36712 22796 36718
rect 22744 36654 22796 36660
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22376 34672 22428 34678
rect 22376 34614 22428 34620
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22296 33454 22324 33526
rect 22284 33448 22336 33454
rect 22284 33390 22336 33396
rect 22204 33272 22324 33300
rect 22100 32836 22152 32842
rect 22100 32778 22152 32784
rect 22008 31748 22060 31754
rect 22112 31736 22140 32778
rect 22296 32502 22324 33272
rect 22374 33008 22430 33017
rect 22374 32943 22430 32952
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22060 31708 22140 31736
rect 22008 31690 22060 31696
rect 22204 31686 22232 32370
rect 22284 32292 22336 32298
rect 22284 32234 22336 32240
rect 22296 31890 22324 32234
rect 22284 31884 22336 31890
rect 22284 31826 22336 31832
rect 22192 31680 22244 31686
rect 22112 31640 22192 31668
rect 21916 31272 21968 31278
rect 21916 31214 21968 31220
rect 21928 29714 21956 31214
rect 22008 30048 22060 30054
rect 22008 29990 22060 29996
rect 21916 29708 21968 29714
rect 21916 29650 21968 29656
rect 22020 29510 22048 29990
rect 22008 29504 22060 29510
rect 22008 29446 22060 29452
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 22112 29209 22140 31640
rect 22192 31622 22244 31628
rect 22388 31210 22416 32943
rect 22572 32366 22600 35090
rect 22664 33153 22692 36654
rect 22744 36576 22796 36582
rect 22744 36518 22796 36524
rect 22650 33144 22706 33153
rect 22650 33079 22706 33088
rect 22756 32994 22784 36518
rect 22664 32966 22784 32994
rect 22560 32360 22612 32366
rect 22560 32302 22612 32308
rect 22664 32212 22692 32966
rect 22848 32570 22876 38372
rect 23296 38276 23348 38282
rect 23296 38218 23348 38224
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23308 37262 23336 38218
rect 23400 37913 23428 38927
rect 23386 37904 23442 37913
rect 23386 37839 23388 37848
rect 23440 37839 23442 37848
rect 23388 37810 23440 37816
rect 23492 37738 23520 44118
rect 23572 42696 23624 42702
rect 23572 42638 23624 42644
rect 23584 42294 23612 42638
rect 23572 42288 23624 42294
rect 23572 42230 23624 42236
rect 23676 41274 23704 44678
rect 23768 42566 23796 45494
rect 23848 45484 23900 45490
rect 23848 45426 23900 45432
rect 23860 44305 23888 45426
rect 24032 45416 24084 45422
rect 24032 45358 24084 45364
rect 24124 45416 24176 45422
rect 24124 45358 24176 45364
rect 23940 44940 23992 44946
rect 23940 44882 23992 44888
rect 23952 44334 23980 44882
rect 24044 44878 24072 45358
rect 24032 44872 24084 44878
rect 24032 44814 24084 44820
rect 23940 44328 23992 44334
rect 23846 44296 23902 44305
rect 23940 44270 23992 44276
rect 23846 44231 23902 44240
rect 24136 43994 24164 45358
rect 24124 43988 24176 43994
rect 24124 43930 24176 43936
rect 23756 42560 23808 42566
rect 23756 42502 23808 42508
rect 23756 42016 23808 42022
rect 23756 41958 23808 41964
rect 24216 42016 24268 42022
rect 24216 41958 24268 41964
rect 23768 41750 23796 41958
rect 23756 41744 23808 41750
rect 23756 41686 23808 41692
rect 23768 41546 23796 41686
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 23756 41540 23808 41546
rect 23756 41482 23808 41488
rect 23664 41268 23716 41274
rect 23664 41210 23716 41216
rect 23572 41132 23624 41138
rect 23572 41074 23624 41080
rect 23584 40730 23612 41074
rect 23940 41064 23992 41070
rect 23940 41006 23992 41012
rect 24032 41064 24084 41070
rect 24032 41006 24084 41012
rect 23572 40724 23624 40730
rect 23572 40666 23624 40672
rect 23848 40588 23900 40594
rect 23848 40530 23900 40536
rect 23756 40180 23808 40186
rect 23860 40168 23888 40530
rect 23808 40140 23888 40168
rect 23756 40122 23808 40128
rect 23756 39908 23808 39914
rect 23756 39850 23808 39856
rect 23768 39098 23796 39850
rect 23756 39092 23808 39098
rect 23756 39034 23808 39040
rect 23572 38208 23624 38214
rect 23572 38150 23624 38156
rect 23664 38208 23716 38214
rect 23664 38150 23716 38156
rect 23388 37732 23440 37738
rect 23388 37674 23440 37680
rect 23480 37732 23532 37738
rect 23480 37674 23532 37680
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23296 37120 23348 37126
rect 23296 37062 23348 37068
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23204 34740 23256 34746
rect 23204 34682 23256 34688
rect 22928 34672 22980 34678
rect 23216 34649 23244 34682
rect 22928 34614 22980 34620
rect 23202 34640 23258 34649
rect 22940 34406 22968 34614
rect 23202 34575 23258 34584
rect 22928 34400 22980 34406
rect 22928 34342 22980 34348
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 22940 33017 22968 33050
rect 22926 33008 22982 33017
rect 22926 32943 22982 32952
rect 22836 32564 22888 32570
rect 22480 32184 22692 32212
rect 22756 32524 22836 32552
rect 22376 31204 22428 31210
rect 22376 31146 22428 31152
rect 22192 30660 22244 30666
rect 22192 30602 22244 30608
rect 22204 30258 22232 30602
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22098 29200 22154 29209
rect 22098 29135 22154 29144
rect 22296 28558 22324 29990
rect 22376 29640 22428 29646
rect 22376 29582 22428 29588
rect 22388 29306 22416 29582
rect 22376 29300 22428 29306
rect 22376 29242 22428 29248
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 21284 22066 21588 22094
rect 21744 22066 21864 22094
rect 21560 14822 21588 22066
rect 21836 16522 21864 22066
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21836 11626 21864 16458
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 13636 2372 13688 2378
rect 13636 2314 13688 2320
rect 15488 800 15516 2450
rect 17880 2446 17908 4422
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18800 800 18828 2450
rect 19628 2446 19656 6598
rect 21376 5710 21404 11494
rect 21928 11218 21956 18566
rect 22204 11218 22232 19450
rect 22296 19378 22324 26726
rect 22480 22094 22508 32184
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22572 30938 22600 31214
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22664 29102 22692 31962
rect 22756 30394 22784 32524
rect 22836 32506 22888 32512
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22652 29096 22704 29102
rect 22652 29038 22704 29044
rect 22480 22066 22692 22094
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22664 15162 22692 22066
rect 22848 15978 22876 32370
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 23308 30938 23336 37062
rect 23400 35630 23428 37674
rect 23388 35624 23440 35630
rect 23386 35592 23388 35601
rect 23440 35592 23442 35601
rect 23386 35527 23442 35536
rect 23388 35488 23440 35494
rect 23386 35456 23388 35465
rect 23440 35456 23442 35465
rect 23386 35391 23442 35400
rect 23400 34785 23428 35391
rect 23386 34776 23442 34785
rect 23386 34711 23442 34720
rect 23584 34202 23612 38150
rect 23676 35290 23704 38150
rect 23756 37868 23808 37874
rect 23756 37810 23808 37816
rect 23768 36378 23796 37810
rect 23860 37670 23888 40140
rect 23952 39846 23980 41006
rect 23940 39840 23992 39846
rect 23940 39782 23992 39788
rect 24044 39098 24072 41006
rect 24032 39092 24084 39098
rect 24032 39034 24084 39040
rect 23848 37664 23900 37670
rect 23848 37606 23900 37612
rect 23940 37324 23992 37330
rect 23940 37266 23992 37272
rect 24032 37324 24084 37330
rect 24032 37266 24084 37272
rect 23848 36712 23900 36718
rect 23848 36654 23900 36660
rect 23860 36378 23888 36654
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23848 36372 23900 36378
rect 23848 36314 23900 36320
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 23860 36009 23888 36042
rect 23846 36000 23902 36009
rect 23846 35935 23902 35944
rect 23860 35766 23888 35935
rect 23848 35760 23900 35766
rect 23848 35702 23900 35708
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23756 35148 23808 35154
rect 23756 35090 23808 35096
rect 23664 34740 23716 34746
rect 23664 34682 23716 34688
rect 23572 34196 23624 34202
rect 23572 34138 23624 34144
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 23584 32842 23612 32982
rect 23676 32978 23704 34682
rect 23664 32972 23716 32978
rect 23664 32914 23716 32920
rect 23572 32836 23624 32842
rect 23572 32778 23624 32784
rect 23388 31136 23440 31142
rect 23388 31078 23440 31084
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 23400 30394 23428 31078
rect 23584 30802 23612 32778
rect 23676 32026 23704 32914
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23572 30796 23624 30802
rect 23572 30738 23624 30744
rect 23388 30388 23440 30394
rect 23388 30330 23440 30336
rect 23584 30326 23612 30738
rect 23664 30592 23716 30598
rect 23664 30534 23716 30540
rect 23676 30394 23704 30534
rect 23664 30388 23716 30394
rect 23664 30330 23716 30336
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23768 28694 23796 35090
rect 23860 34406 23888 35702
rect 23848 34400 23900 34406
rect 23848 34342 23900 34348
rect 23952 33658 23980 37266
rect 24044 34746 24072 37266
rect 24032 34740 24084 34746
rect 24032 34682 24084 34688
rect 24136 34134 24164 41550
rect 24228 41070 24256 41958
rect 24216 41064 24268 41070
rect 24216 41006 24268 41012
rect 24320 40526 24348 46038
rect 24400 44736 24452 44742
rect 24400 44678 24452 44684
rect 24412 43110 24440 44678
rect 24504 44538 24532 50866
rect 24780 48890 24808 52498
rect 24872 50794 24900 53110
rect 25320 52896 25372 52902
rect 25320 52838 25372 52844
rect 24952 52352 25004 52358
rect 24952 52294 25004 52300
rect 24860 50788 24912 50794
rect 24860 50730 24912 50736
rect 24964 49434 24992 52294
rect 24952 49428 25004 49434
rect 24952 49370 25004 49376
rect 24768 48884 24820 48890
rect 24768 48826 24820 48832
rect 25044 48748 25096 48754
rect 25044 48690 25096 48696
rect 24676 48136 24728 48142
rect 24676 48078 24728 48084
rect 24584 48068 24636 48074
rect 24584 48010 24636 48016
rect 24596 47666 24624 48010
rect 24584 47660 24636 47666
rect 24584 47602 24636 47608
rect 24596 46986 24624 47602
rect 24584 46980 24636 46986
rect 24584 46922 24636 46928
rect 24688 46646 24716 48078
rect 24768 48000 24820 48006
rect 24768 47942 24820 47948
rect 24780 47598 24808 47942
rect 24768 47592 24820 47598
rect 24768 47534 24820 47540
rect 24860 47116 24912 47122
rect 24860 47058 24912 47064
rect 24872 46730 24900 47058
rect 24952 47048 25004 47054
rect 24952 46990 25004 46996
rect 24780 46714 24900 46730
rect 24768 46708 24900 46714
rect 24820 46702 24900 46708
rect 24768 46650 24820 46656
rect 24676 46640 24728 46646
rect 24676 46582 24728 46588
rect 24860 46572 24912 46578
rect 24860 46514 24912 46520
rect 24768 45280 24820 45286
rect 24768 45222 24820 45228
rect 24780 45064 24808 45222
rect 24596 45036 24808 45064
rect 24492 44532 24544 44538
rect 24492 44474 24544 44480
rect 24596 43790 24624 45036
rect 24768 44804 24820 44810
rect 24872 44792 24900 46514
rect 24820 44764 24900 44792
rect 24768 44746 24820 44752
rect 24584 43784 24636 43790
rect 24584 43726 24636 43732
rect 24492 43716 24544 43722
rect 24492 43658 24544 43664
rect 24676 43716 24728 43722
rect 24676 43658 24728 43664
rect 24400 43104 24452 43110
rect 24400 43046 24452 43052
rect 24412 42362 24440 43046
rect 24400 42356 24452 42362
rect 24400 42298 24452 42304
rect 24504 41818 24532 43658
rect 24492 41812 24544 41818
rect 24492 41754 24544 41760
rect 24584 41676 24636 41682
rect 24584 41618 24636 41624
rect 24308 40520 24360 40526
rect 24308 40462 24360 40468
rect 24596 40050 24624 41618
rect 24688 41414 24716 43658
rect 24780 42158 24808 44746
rect 24964 44418 24992 46990
rect 25056 46170 25084 48690
rect 25228 48340 25280 48346
rect 25228 48282 25280 48288
rect 25136 48068 25188 48074
rect 25136 48010 25188 48016
rect 25148 47734 25176 48010
rect 25136 47728 25188 47734
rect 25136 47670 25188 47676
rect 25136 47456 25188 47462
rect 25136 47398 25188 47404
rect 25044 46164 25096 46170
rect 25044 46106 25096 46112
rect 25044 45484 25096 45490
rect 25044 45426 25096 45432
rect 25056 44742 25084 45426
rect 25044 44736 25096 44742
rect 25044 44678 25096 44684
rect 24964 44390 25084 44418
rect 24952 44328 25004 44334
rect 24952 44270 25004 44276
rect 24860 43648 24912 43654
rect 24860 43590 24912 43596
rect 24872 42242 24900 43590
rect 24964 43382 24992 44270
rect 25056 43722 25084 44390
rect 25044 43716 25096 43722
rect 25044 43658 25096 43664
rect 24952 43376 25004 43382
rect 24952 43318 25004 43324
rect 24964 42362 24992 43318
rect 25044 42900 25096 42906
rect 25044 42842 25096 42848
rect 25056 42702 25084 42842
rect 25148 42838 25176 47398
rect 25240 46374 25268 48282
rect 25332 47138 25360 52838
rect 25424 51074 25452 53926
rect 26068 51074 26096 53926
rect 26240 53576 26292 53582
rect 26240 53518 26292 53524
rect 25424 51046 25820 51074
rect 25596 50244 25648 50250
rect 25596 50186 25648 50192
rect 25412 49224 25464 49230
rect 25412 49166 25464 49172
rect 25424 48210 25452 49166
rect 25412 48204 25464 48210
rect 25412 48146 25464 48152
rect 25504 48068 25556 48074
rect 25504 48010 25556 48016
rect 25516 47666 25544 48010
rect 25504 47660 25556 47666
rect 25504 47602 25556 47608
rect 25504 47456 25556 47462
rect 25504 47398 25556 47404
rect 25516 47190 25544 47398
rect 25504 47184 25556 47190
rect 25332 47110 25452 47138
rect 25504 47126 25556 47132
rect 25320 47048 25372 47054
rect 25318 47016 25320 47025
rect 25372 47016 25374 47025
rect 25318 46951 25374 46960
rect 25228 46368 25280 46374
rect 25228 46310 25280 46316
rect 25320 46368 25372 46374
rect 25320 46310 25372 46316
rect 25228 43716 25280 43722
rect 25228 43658 25280 43664
rect 25136 42832 25188 42838
rect 25136 42774 25188 42780
rect 25044 42696 25096 42702
rect 25044 42638 25096 42644
rect 25044 42560 25096 42566
rect 25044 42502 25096 42508
rect 24952 42356 25004 42362
rect 24952 42298 25004 42304
rect 24872 42214 24992 42242
rect 24768 42152 24820 42158
rect 24768 42094 24820 42100
rect 24858 41440 24914 41449
rect 24688 41386 24808 41414
rect 24780 41274 24808 41386
rect 24858 41375 24914 41384
rect 24768 41268 24820 41274
rect 24768 41210 24820 41216
rect 24872 41002 24900 41375
rect 24860 40996 24912 41002
rect 24860 40938 24912 40944
rect 24872 40066 24900 40938
rect 24964 40730 24992 42214
rect 24952 40724 25004 40730
rect 24952 40666 25004 40672
rect 24584 40044 24636 40050
rect 24584 39986 24636 39992
rect 24780 40038 24900 40066
rect 24952 40112 25004 40118
rect 24952 40054 25004 40060
rect 24492 39840 24544 39846
rect 24492 39782 24544 39788
rect 24400 39636 24452 39642
rect 24400 39578 24452 39584
rect 24412 39545 24440 39578
rect 24398 39536 24454 39545
rect 24398 39471 24454 39480
rect 24504 38826 24532 39782
rect 24676 39092 24728 39098
rect 24676 39034 24728 39040
rect 24584 38956 24636 38962
rect 24584 38898 24636 38904
rect 24596 38865 24624 38898
rect 24582 38856 24638 38865
rect 24492 38820 24544 38826
rect 24582 38791 24638 38800
rect 24492 38762 24544 38768
rect 24584 38752 24636 38758
rect 24584 38694 24636 38700
rect 24398 37904 24454 37913
rect 24398 37839 24454 37848
rect 24412 36854 24440 37839
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24412 36009 24440 36790
rect 24596 36718 24624 38694
rect 24688 38536 24716 39034
rect 24780 38894 24808 40038
rect 24768 38888 24820 38894
rect 24768 38830 24820 38836
rect 24780 38758 24808 38830
rect 24768 38752 24820 38758
rect 24768 38694 24820 38700
rect 24964 38554 24992 40054
rect 25056 39642 25084 42502
rect 25136 42152 25188 42158
rect 25136 42094 25188 42100
rect 25148 41682 25176 42094
rect 25136 41676 25188 41682
rect 25136 41618 25188 41624
rect 25240 41414 25268 43658
rect 25332 41562 25360 46310
rect 25424 46170 25452 47110
rect 25412 46164 25464 46170
rect 25412 46106 25464 46112
rect 25424 45626 25452 46106
rect 25504 45960 25556 45966
rect 25504 45902 25556 45908
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 25332 41546 25452 41562
rect 25332 41540 25464 41546
rect 25332 41534 25412 41540
rect 25332 41449 25360 41534
rect 25412 41482 25464 41488
rect 25148 41386 25268 41414
rect 25318 41440 25374 41449
rect 25044 39636 25096 39642
rect 25044 39578 25096 39584
rect 25148 39506 25176 41386
rect 25318 41375 25374 41384
rect 25226 41304 25282 41313
rect 25226 41239 25228 41248
rect 25280 41239 25282 41248
rect 25228 41210 25280 41216
rect 25516 41002 25544 45902
rect 25608 44946 25636 50186
rect 25688 49156 25740 49162
rect 25688 49098 25740 49104
rect 25700 47802 25728 49098
rect 25688 47796 25740 47802
rect 25688 47738 25740 47744
rect 25688 47660 25740 47666
rect 25688 47602 25740 47608
rect 25700 47258 25728 47602
rect 25688 47252 25740 47258
rect 25688 47194 25740 47200
rect 25700 46646 25728 47194
rect 25792 46986 25820 51046
rect 25976 51046 26096 51074
rect 26252 51066 26280 53518
rect 27344 53100 27396 53106
rect 27344 53042 27396 53048
rect 27356 51066 27384 53042
rect 26240 51060 26292 51066
rect 25872 50380 25924 50386
rect 25872 50322 25924 50328
rect 25884 47122 25912 50322
rect 25872 47116 25924 47122
rect 25872 47058 25924 47064
rect 25780 46980 25832 46986
rect 25780 46922 25832 46928
rect 25688 46640 25740 46646
rect 25688 46582 25740 46588
rect 25596 44940 25648 44946
rect 25596 44882 25648 44888
rect 25596 44804 25648 44810
rect 25700 44792 25728 46582
rect 25872 46504 25924 46510
rect 25872 46446 25924 46452
rect 25884 45014 25912 46446
rect 25976 45966 26004 51046
rect 26240 51002 26292 51008
rect 27344 51060 27396 51066
rect 27344 51002 27396 51008
rect 26700 50720 26752 50726
rect 26700 50662 26752 50668
rect 26332 49972 26384 49978
rect 26332 49914 26384 49920
rect 26056 48204 26108 48210
rect 26056 48146 26108 48152
rect 26068 47122 26096 48146
rect 26240 47660 26292 47666
rect 26240 47602 26292 47608
rect 26056 47116 26108 47122
rect 26056 47058 26108 47064
rect 26068 46714 26096 47058
rect 26148 46980 26200 46986
rect 26148 46922 26200 46928
rect 26056 46708 26108 46714
rect 26056 46650 26108 46656
rect 26160 46510 26188 46922
rect 26252 46753 26280 47602
rect 26238 46744 26294 46753
rect 26238 46679 26294 46688
rect 26148 46504 26200 46510
rect 26148 46446 26200 46452
rect 25964 45960 26016 45966
rect 25964 45902 26016 45908
rect 26344 45558 26372 49914
rect 26608 49836 26660 49842
rect 26608 49778 26660 49784
rect 26424 48680 26476 48686
rect 26424 48622 26476 48628
rect 26516 48680 26568 48686
rect 26516 48622 26568 48628
rect 26436 45626 26464 48622
rect 26424 45620 26476 45626
rect 26424 45562 26476 45568
rect 26332 45552 26384 45558
rect 26332 45494 26384 45500
rect 25872 45008 25924 45014
rect 25872 44950 25924 44956
rect 25648 44764 25728 44792
rect 25596 44746 25648 44752
rect 25608 44402 25636 44746
rect 25596 44396 25648 44402
rect 25596 44338 25648 44344
rect 26332 44396 26384 44402
rect 26332 44338 26384 44344
rect 25608 43722 25636 44338
rect 26148 44328 26200 44334
rect 26148 44270 26200 44276
rect 25872 44260 25924 44266
rect 25872 44202 25924 44208
rect 25596 43716 25648 43722
rect 25596 43658 25648 43664
rect 25608 43382 25636 43658
rect 25596 43376 25648 43382
rect 25596 43318 25648 43324
rect 25608 42770 25636 43318
rect 25596 42764 25648 42770
rect 25596 42706 25648 42712
rect 25608 41546 25636 42706
rect 25596 41540 25648 41546
rect 25596 41482 25648 41488
rect 25504 40996 25556 41002
rect 25504 40938 25556 40944
rect 25516 40662 25544 40938
rect 25504 40656 25556 40662
rect 25504 40598 25556 40604
rect 25504 40112 25556 40118
rect 25608 40100 25636 41482
rect 25884 41414 25912 44202
rect 25556 40072 25636 40100
rect 25792 41386 25912 41414
rect 25504 40054 25556 40060
rect 25136 39500 25188 39506
rect 25136 39442 25188 39448
rect 25412 39432 25464 39438
rect 25412 39374 25464 39380
rect 24952 38548 25004 38554
rect 24688 38508 24808 38536
rect 24676 38412 24728 38418
rect 24676 38354 24728 38360
rect 24584 36712 24636 36718
rect 24584 36654 24636 36660
rect 24688 36378 24716 38354
rect 24780 37913 24808 38508
rect 24952 38490 25004 38496
rect 25320 38208 25372 38214
rect 25424 38185 25452 39374
rect 25320 38150 25372 38156
rect 25410 38176 25466 38185
rect 24766 37904 24822 37913
rect 24766 37839 24768 37848
rect 24820 37839 24822 37848
rect 24860 37868 24912 37874
rect 24768 37810 24820 37816
rect 24860 37810 24912 37816
rect 24676 36372 24728 36378
rect 24676 36314 24728 36320
rect 24584 36236 24636 36242
rect 24584 36178 24636 36184
rect 24492 36100 24544 36106
rect 24492 36042 24544 36048
rect 24398 36000 24454 36009
rect 24398 35935 24454 35944
rect 24504 35154 24532 36042
rect 24596 35494 24624 36178
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24596 35154 24624 35430
rect 24492 35148 24544 35154
rect 24492 35090 24544 35096
rect 24584 35148 24636 35154
rect 24584 35090 24636 35096
rect 24400 34740 24452 34746
rect 24400 34682 24452 34688
rect 24412 34406 24440 34682
rect 24400 34400 24452 34406
rect 24400 34342 24452 34348
rect 24124 34128 24176 34134
rect 24124 34070 24176 34076
rect 23940 33652 23992 33658
rect 23940 33594 23992 33600
rect 23848 32768 23900 32774
rect 23848 32710 23900 32716
rect 23860 32502 23888 32710
rect 23952 32502 23980 33594
rect 24032 33448 24084 33454
rect 24032 33390 24084 33396
rect 24412 33436 24440 34342
rect 24596 33590 24624 35090
rect 24688 34678 24716 36314
rect 24676 34672 24728 34678
rect 24676 34614 24728 34620
rect 24584 33584 24636 33590
rect 24584 33526 24636 33532
rect 24676 33584 24728 33590
rect 24676 33526 24728 33532
rect 24688 33436 24716 33526
rect 24412 33408 24716 33436
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23940 32496 23992 32502
rect 23940 32438 23992 32444
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23952 31890 23980 32166
rect 24044 32026 24072 33390
rect 24412 32502 24440 33408
rect 24872 33114 24900 37810
rect 25044 37800 25096 37806
rect 25044 37742 25096 37748
rect 25228 37800 25280 37806
rect 25228 37742 25280 37748
rect 25056 36122 25084 37742
rect 25240 36961 25268 37742
rect 25226 36952 25282 36961
rect 25226 36887 25282 36896
rect 25228 36780 25280 36786
rect 25228 36722 25280 36728
rect 25136 36712 25188 36718
rect 25136 36654 25188 36660
rect 24964 36094 25084 36122
rect 25148 36106 25176 36654
rect 25136 36100 25188 36106
rect 24964 35630 24992 36094
rect 25136 36042 25188 36048
rect 24952 35624 25004 35630
rect 24952 35566 25004 35572
rect 24964 35290 24992 35566
rect 25044 35488 25096 35494
rect 25044 35430 25096 35436
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 25056 35018 25084 35430
rect 25044 35012 25096 35018
rect 25044 34954 25096 34960
rect 25240 33998 25268 36722
rect 25332 34898 25360 38150
rect 25410 38111 25466 38120
rect 25424 35578 25452 38111
rect 25516 36106 25544 40054
rect 25792 39030 25820 41386
rect 25872 40384 25924 40390
rect 25872 40326 25924 40332
rect 25884 39642 25912 40326
rect 25964 39840 26016 39846
rect 25964 39782 26016 39788
rect 25872 39636 25924 39642
rect 25872 39578 25924 39584
rect 25780 39024 25832 39030
rect 25780 38966 25832 38972
rect 25688 38548 25740 38554
rect 25688 38490 25740 38496
rect 25596 38480 25648 38486
rect 25596 38422 25648 38428
rect 25504 36100 25556 36106
rect 25504 36042 25556 36048
rect 25516 36009 25544 36042
rect 25502 36000 25558 36009
rect 25502 35935 25558 35944
rect 25424 35550 25544 35578
rect 25332 34870 25452 34898
rect 25228 33992 25280 33998
rect 25148 33952 25228 33980
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24400 32496 24452 32502
rect 24400 32438 24452 32444
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 23940 31884 23992 31890
rect 23940 31826 23992 31832
rect 23952 30802 23980 31826
rect 25148 31210 25176 33952
rect 25228 33934 25280 33940
rect 25228 33448 25280 33454
rect 25228 33390 25280 33396
rect 25136 31204 25188 31210
rect 25136 31146 25188 31152
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 23940 30796 23992 30802
rect 23940 30738 23992 30744
rect 24964 30734 24992 31078
rect 25240 30802 25268 33390
rect 25424 32910 25452 34870
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25320 32836 25372 32842
rect 25320 32778 25372 32784
rect 25228 30796 25280 30802
rect 25228 30738 25280 30744
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24492 29504 24544 29510
rect 24492 29446 24544 29452
rect 24504 29238 24532 29446
rect 25332 29306 25360 32778
rect 25516 31754 25544 35550
rect 25608 34746 25636 38422
rect 25700 38321 25728 38490
rect 25792 38418 25820 38966
rect 25780 38412 25832 38418
rect 25780 38354 25832 38360
rect 25686 38312 25742 38321
rect 25686 38247 25742 38256
rect 25700 38214 25728 38247
rect 25688 38208 25740 38214
rect 25688 38150 25740 38156
rect 25870 37904 25926 37913
rect 25870 37839 25872 37848
rect 25924 37839 25926 37848
rect 25872 37810 25924 37816
rect 25872 37732 25924 37738
rect 25872 37674 25924 37680
rect 25884 36038 25912 37674
rect 25976 36718 26004 39782
rect 26056 39296 26108 39302
rect 26056 39238 26108 39244
rect 26068 37194 26096 39238
rect 26056 37188 26108 37194
rect 26056 37130 26108 37136
rect 25964 36712 26016 36718
rect 25964 36654 26016 36660
rect 26056 36712 26108 36718
rect 26056 36654 26108 36660
rect 26068 36145 26096 36654
rect 26160 36650 26188 44270
rect 26238 40488 26294 40497
rect 26238 40423 26240 40432
rect 26292 40423 26294 40432
rect 26240 40394 26292 40400
rect 26344 39817 26372 44338
rect 26528 44282 26556 48622
rect 26620 45506 26648 49778
rect 26712 46034 26740 50662
rect 27344 49700 27396 49706
rect 27344 49642 27396 49648
rect 27160 49632 27212 49638
rect 27160 49574 27212 49580
rect 27172 49366 27200 49574
rect 27160 49360 27212 49366
rect 27160 49302 27212 49308
rect 26792 49224 26844 49230
rect 26976 49224 27028 49230
rect 26844 49184 26924 49212
rect 26792 49166 26844 49172
rect 26792 47796 26844 47802
rect 26792 47738 26844 47744
rect 26804 47122 26832 47738
rect 26896 47258 26924 49184
rect 26976 49166 27028 49172
rect 26884 47252 26936 47258
rect 26884 47194 26936 47200
rect 26896 47161 26924 47194
rect 26882 47152 26938 47161
rect 26792 47116 26844 47122
rect 26882 47087 26938 47096
rect 26792 47058 26844 47064
rect 26804 46714 26832 47058
rect 26896 46986 26924 47087
rect 26884 46980 26936 46986
rect 26884 46922 26936 46928
rect 26792 46708 26844 46714
rect 26792 46650 26844 46656
rect 26988 46102 27016 49166
rect 27252 49088 27304 49094
rect 27252 49030 27304 49036
rect 27264 48822 27292 49030
rect 27252 48816 27304 48822
rect 27252 48758 27304 48764
rect 27068 48544 27120 48550
rect 27068 48486 27120 48492
rect 27160 48544 27212 48550
rect 27160 48486 27212 48492
rect 26976 46096 27028 46102
rect 26976 46038 27028 46044
rect 26700 46028 26752 46034
rect 26700 45970 26752 45976
rect 26792 46028 26844 46034
rect 26792 45970 26844 45976
rect 26804 45830 26832 45970
rect 26700 45824 26752 45830
rect 26700 45766 26752 45772
rect 26792 45824 26844 45830
rect 26792 45766 26844 45772
rect 26712 45626 26740 45766
rect 26700 45620 26752 45626
rect 26700 45562 26752 45568
rect 26620 45478 26740 45506
rect 26608 45416 26660 45422
rect 26608 45358 26660 45364
rect 26620 44742 26648 45358
rect 26608 44736 26660 44742
rect 26608 44678 26660 44684
rect 26436 44254 26556 44282
rect 26436 43450 26464 44254
rect 26516 44192 26568 44198
rect 26516 44134 26568 44140
rect 26424 43444 26476 43450
rect 26424 43386 26476 43392
rect 26436 41682 26464 43386
rect 26424 41676 26476 41682
rect 26424 41618 26476 41624
rect 26424 40384 26476 40390
rect 26424 40326 26476 40332
rect 26330 39808 26386 39817
rect 26330 39743 26386 39752
rect 26332 39296 26384 39302
rect 26332 39238 26384 39244
rect 26344 39098 26372 39238
rect 26332 39092 26384 39098
rect 26332 39034 26384 39040
rect 26344 39001 26372 39034
rect 26330 38992 26386 39001
rect 26330 38927 26386 38936
rect 26240 38752 26292 38758
rect 26240 38694 26292 38700
rect 26252 37942 26280 38694
rect 26436 38282 26464 40326
rect 26528 39914 26556 44134
rect 26620 43994 26648 44678
rect 26608 43988 26660 43994
rect 26608 43930 26660 43936
rect 26620 42838 26648 43930
rect 26712 43450 26740 45478
rect 26700 43444 26752 43450
rect 26700 43386 26752 43392
rect 26698 43208 26754 43217
rect 26698 43143 26754 43152
rect 26712 42906 26740 43143
rect 26700 42900 26752 42906
rect 26700 42842 26752 42848
rect 26608 42832 26660 42838
rect 26608 42774 26660 42780
rect 26608 42016 26660 42022
rect 26608 41958 26660 41964
rect 26620 41750 26648 41958
rect 26608 41744 26660 41750
rect 26608 41686 26660 41692
rect 26606 41576 26662 41585
rect 26606 41511 26662 41520
rect 26620 41478 26648 41511
rect 26608 41472 26660 41478
rect 26608 41414 26660 41420
rect 26804 41414 26832 45766
rect 26976 45416 27028 45422
rect 26976 45358 27028 45364
rect 26884 42696 26936 42702
rect 26884 42638 26936 42644
rect 26896 42226 26924 42638
rect 26884 42220 26936 42226
rect 26884 42162 26936 42168
rect 26988 41614 27016 45358
rect 27080 45082 27108 48486
rect 27172 48346 27200 48486
rect 27160 48340 27212 48346
rect 27160 48282 27212 48288
rect 27252 48000 27304 48006
rect 27252 47942 27304 47948
rect 27264 47530 27292 47942
rect 27252 47524 27304 47530
rect 27252 47466 27304 47472
rect 27356 47138 27384 49642
rect 27448 48754 27476 53926
rect 27528 50924 27580 50930
rect 27528 50866 27580 50872
rect 27540 50522 27568 50866
rect 27528 50516 27580 50522
rect 27528 50458 27580 50464
rect 27620 50448 27672 50454
rect 27540 50396 27620 50402
rect 27540 50390 27672 50396
rect 27540 50374 27660 50390
rect 27436 48748 27488 48754
rect 27436 48690 27488 48696
rect 27436 48068 27488 48074
rect 27436 48010 27488 48016
rect 27448 47598 27476 48010
rect 27540 47716 27568 50374
rect 27620 49768 27672 49774
rect 27620 49710 27672 49716
rect 27632 48192 27660 49710
rect 27724 48346 27752 54062
rect 27896 54052 27948 54058
rect 27896 53994 27948 54000
rect 27908 53530 27936 53994
rect 28276 53802 28304 54198
rect 28368 54194 28396 56222
rect 28630 56200 28686 57000
rect 29274 56200 29330 57000
rect 29918 56200 29974 57000
rect 30024 56222 30328 56250
rect 28356 54188 28408 54194
rect 28356 54130 28408 54136
rect 28356 53984 28408 53990
rect 28408 53944 28488 53972
rect 28356 53926 28408 53932
rect 28276 53774 28396 53802
rect 27816 53502 27936 53530
rect 27712 48340 27764 48346
rect 27712 48282 27764 48288
rect 27712 48204 27764 48210
rect 27632 48164 27712 48192
rect 27712 48146 27764 48152
rect 27712 48000 27764 48006
rect 27712 47942 27764 47948
rect 27620 47728 27672 47734
rect 27540 47688 27620 47716
rect 27620 47670 27672 47676
rect 27436 47592 27488 47598
rect 27436 47534 27488 47540
rect 27448 47240 27476 47534
rect 27528 47252 27580 47258
rect 27448 47212 27528 47240
rect 27528 47194 27580 47200
rect 27620 47184 27672 47190
rect 27264 47110 27384 47138
rect 27618 47152 27620 47161
rect 27672 47152 27674 47161
rect 27068 45076 27120 45082
rect 27068 45018 27120 45024
rect 27264 44946 27292 47110
rect 27618 47087 27674 47096
rect 27618 46744 27674 46753
rect 27618 46679 27674 46688
rect 27528 46436 27580 46442
rect 27528 46378 27580 46384
rect 27342 46064 27398 46073
rect 27342 45999 27398 46008
rect 27356 45966 27384 45999
rect 27344 45960 27396 45966
rect 27344 45902 27396 45908
rect 27252 44940 27304 44946
rect 27252 44882 27304 44888
rect 27344 44940 27396 44946
rect 27344 44882 27396 44888
rect 27252 43308 27304 43314
rect 27252 43250 27304 43256
rect 27160 42560 27212 42566
rect 27160 42502 27212 42508
rect 27172 42294 27200 42502
rect 27160 42288 27212 42294
rect 27160 42230 27212 42236
rect 27068 42152 27120 42158
rect 27068 42094 27120 42100
rect 26976 41608 27028 41614
rect 26976 41550 27028 41556
rect 26804 41386 26924 41414
rect 26700 40180 26752 40186
rect 26700 40122 26752 40128
rect 26516 39908 26568 39914
rect 26516 39850 26568 39856
rect 26424 38276 26476 38282
rect 26424 38218 26476 38224
rect 26240 37936 26292 37942
rect 26240 37878 26292 37884
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 26516 37120 26568 37126
rect 26516 37062 26568 37068
rect 26252 36922 26280 37062
rect 26240 36916 26292 36922
rect 26240 36858 26292 36864
rect 26148 36644 26200 36650
rect 26148 36586 26200 36592
rect 26054 36136 26110 36145
rect 26054 36071 26110 36080
rect 25872 36032 25924 36038
rect 25686 36000 25742 36009
rect 25872 35974 25924 35980
rect 25686 35935 25742 35944
rect 25700 35018 25728 35935
rect 25884 35630 25912 35974
rect 25872 35624 25924 35630
rect 25872 35566 25924 35572
rect 25688 35012 25740 35018
rect 25688 34954 25740 34960
rect 25596 34740 25648 34746
rect 25596 34682 25648 34688
rect 25608 33454 25636 34682
rect 25700 34610 25728 34954
rect 25688 34604 25740 34610
rect 25688 34546 25740 34552
rect 25884 34066 25912 35566
rect 26330 35456 26386 35465
rect 26330 35391 26386 35400
rect 25964 34944 26016 34950
rect 25964 34886 26016 34892
rect 25976 34202 26004 34886
rect 26344 34542 26372 35391
rect 26332 34536 26384 34542
rect 26332 34478 26384 34484
rect 25964 34196 26016 34202
rect 25964 34138 26016 34144
rect 25872 34060 25924 34066
rect 25872 34002 25924 34008
rect 25596 33448 25648 33454
rect 25596 33390 25648 33396
rect 26344 31890 26372 34478
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 25516 31726 25636 31754
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 23756 28688 23808 28694
rect 23756 28630 23808 28636
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 25332 16574 25360 29106
rect 25240 16546 25360 16574
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23584 12986 23612 16118
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 24688 12442 24716 15370
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22388 9654 22416 9862
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22296 8090 22324 9454
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22296 5846 22324 8026
rect 22284 5840 22336 5846
rect 22284 5782 22336 5788
rect 22388 5710 22416 9590
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23400 8090 23428 11086
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 22112 800 22140 2450
rect 22204 2446 22232 5578
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23400 4622 23428 8026
rect 24596 6914 24624 11018
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24688 7886 24716 8434
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24596 6886 24716 6914
rect 24688 5710 24716 6886
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 24780 2310 24808 15982
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24872 7274 24900 12786
rect 25240 9586 25268 16546
rect 25608 15570 25636 31726
rect 26528 31278 26556 37062
rect 26712 35193 26740 40122
rect 26896 39982 26924 41386
rect 26884 39976 26936 39982
rect 26884 39918 26936 39924
rect 26896 39506 26924 39918
rect 27080 39506 27108 42094
rect 27160 39840 27212 39846
rect 27160 39782 27212 39788
rect 26884 39500 26936 39506
rect 26884 39442 26936 39448
rect 27068 39500 27120 39506
rect 27068 39442 27120 39448
rect 26976 39364 27028 39370
rect 26976 39306 27028 39312
rect 26884 38412 26936 38418
rect 26884 38354 26936 38360
rect 26698 35184 26754 35193
rect 26698 35119 26754 35128
rect 26516 31272 26568 31278
rect 26516 31214 26568 31220
rect 25872 29572 25924 29578
rect 25872 29514 25924 29520
rect 25596 15564 25648 15570
rect 25596 15506 25648 15512
rect 25504 15088 25556 15094
rect 25504 15030 25556 15036
rect 25516 12442 25544 15030
rect 25504 12436 25556 12442
rect 25504 12378 25556 12384
rect 25320 12232 25372 12238
rect 25320 12174 25372 12180
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25332 11286 25360 12174
rect 25320 11280 25372 11286
rect 25320 11222 25372 11228
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 25240 6914 25268 9522
rect 25332 8634 25360 11222
rect 25516 11218 25544 12174
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25424 9382 25452 9930
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25424 8294 25452 9318
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25240 6886 25360 6914
rect 25228 5636 25280 5642
rect 25228 5578 25280 5584
rect 25240 2446 25268 5578
rect 25332 3942 25360 6886
rect 25608 4554 25636 8570
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25884 3466 25912 29514
rect 26528 28490 26556 31214
rect 26896 30802 26924 38354
rect 26988 31890 27016 39306
rect 27172 38350 27200 39782
rect 27264 39302 27292 43250
rect 27356 41750 27384 44882
rect 27540 44878 27568 46378
rect 27528 44872 27580 44878
rect 27528 44814 27580 44820
rect 27632 44538 27660 46679
rect 27724 45898 27752 47942
rect 27712 45892 27764 45898
rect 27712 45834 27764 45840
rect 27712 45552 27764 45558
rect 27712 45494 27764 45500
rect 27620 44532 27672 44538
rect 27620 44474 27672 44480
rect 27436 44464 27488 44470
rect 27436 44406 27488 44412
rect 27448 44180 27476 44406
rect 27528 44328 27580 44334
rect 27580 44276 27660 44282
rect 27528 44270 27660 44276
rect 27540 44254 27660 44270
rect 27448 44152 27568 44180
rect 27436 43852 27488 43858
rect 27436 43794 27488 43800
rect 27448 42770 27476 43794
rect 27540 43450 27568 44152
rect 27528 43444 27580 43450
rect 27528 43386 27580 43392
rect 27632 42922 27660 44254
rect 27724 43840 27752 45494
rect 27816 44470 27844 53502
rect 27950 53340 28258 53349
rect 27950 53338 27956 53340
rect 28012 53338 28036 53340
rect 28092 53338 28116 53340
rect 28172 53338 28196 53340
rect 28252 53338 28258 53340
rect 28012 53286 28014 53338
rect 28194 53286 28196 53338
rect 27950 53284 27956 53286
rect 28012 53284 28036 53286
rect 28092 53284 28116 53286
rect 28172 53284 28196 53286
rect 28252 53284 28258 53286
rect 27950 53275 28258 53284
rect 27950 52252 28258 52261
rect 27950 52250 27956 52252
rect 28012 52250 28036 52252
rect 28092 52250 28116 52252
rect 28172 52250 28196 52252
rect 28252 52250 28258 52252
rect 28012 52198 28014 52250
rect 28194 52198 28196 52250
rect 27950 52196 27956 52198
rect 28012 52196 28036 52198
rect 28092 52196 28116 52198
rect 28172 52196 28196 52198
rect 28252 52196 28258 52198
rect 27950 52187 28258 52196
rect 27950 51164 28258 51173
rect 27950 51162 27956 51164
rect 28012 51162 28036 51164
rect 28092 51162 28116 51164
rect 28172 51162 28196 51164
rect 28252 51162 28258 51164
rect 28012 51110 28014 51162
rect 28194 51110 28196 51162
rect 27950 51108 27956 51110
rect 28012 51108 28036 51110
rect 28092 51108 28116 51110
rect 28172 51108 28196 51110
rect 28252 51108 28258 51110
rect 27950 51099 28258 51108
rect 27950 50076 28258 50085
rect 27950 50074 27956 50076
rect 28012 50074 28036 50076
rect 28092 50074 28116 50076
rect 28172 50074 28196 50076
rect 28252 50074 28258 50076
rect 28012 50022 28014 50074
rect 28194 50022 28196 50074
rect 27950 50020 27956 50022
rect 28012 50020 28036 50022
rect 28092 50020 28116 50022
rect 28172 50020 28196 50022
rect 28252 50020 28258 50022
rect 27950 50011 28258 50020
rect 27950 48988 28258 48997
rect 27950 48986 27956 48988
rect 28012 48986 28036 48988
rect 28092 48986 28116 48988
rect 28172 48986 28196 48988
rect 28252 48986 28258 48988
rect 28012 48934 28014 48986
rect 28194 48934 28196 48986
rect 27950 48932 27956 48934
rect 28012 48932 28036 48934
rect 28092 48932 28116 48934
rect 28172 48932 28196 48934
rect 28252 48932 28258 48934
rect 27950 48923 28258 48932
rect 28368 48210 28396 53774
rect 28356 48204 28408 48210
rect 28356 48146 28408 48152
rect 27950 47900 28258 47909
rect 27950 47898 27956 47900
rect 28012 47898 28036 47900
rect 28092 47898 28116 47900
rect 28172 47898 28196 47900
rect 28252 47898 28258 47900
rect 28012 47846 28014 47898
rect 28194 47846 28196 47898
rect 27950 47844 27956 47846
rect 28012 47844 28036 47846
rect 28092 47844 28116 47846
rect 28172 47844 28196 47846
rect 28252 47844 28258 47846
rect 27950 47835 28258 47844
rect 28264 47796 28316 47802
rect 28264 47738 28316 47744
rect 28276 46968 28304 47738
rect 28356 47660 28408 47666
rect 28356 47602 28408 47608
rect 28368 47258 28396 47602
rect 28356 47252 28408 47258
rect 28356 47194 28408 47200
rect 28356 46980 28408 46986
rect 28276 46940 28356 46968
rect 28356 46922 28408 46928
rect 27950 46812 28258 46821
rect 27950 46810 27956 46812
rect 28012 46810 28036 46812
rect 28092 46810 28116 46812
rect 28172 46810 28196 46812
rect 28252 46810 28258 46812
rect 28012 46758 28014 46810
rect 28194 46758 28196 46810
rect 27950 46756 27956 46758
rect 28012 46756 28036 46758
rect 28092 46756 28116 46758
rect 28172 46756 28196 46758
rect 28252 46756 28258 46758
rect 27950 46747 28258 46756
rect 27896 46640 27948 46646
rect 27896 46582 27948 46588
rect 27908 45937 27936 46582
rect 27894 45928 27950 45937
rect 27894 45863 27950 45872
rect 27950 45724 28258 45733
rect 27950 45722 27956 45724
rect 28012 45722 28036 45724
rect 28092 45722 28116 45724
rect 28172 45722 28196 45724
rect 28252 45722 28258 45724
rect 28012 45670 28014 45722
rect 28194 45670 28196 45722
rect 27950 45668 27956 45670
rect 28012 45668 28036 45670
rect 28092 45668 28116 45670
rect 28172 45668 28196 45670
rect 28252 45668 28258 45670
rect 27950 45659 28258 45668
rect 28172 45620 28224 45626
rect 28172 45562 28224 45568
rect 28264 45620 28316 45626
rect 28264 45562 28316 45568
rect 28184 45286 28212 45562
rect 28172 45280 28224 45286
rect 28172 45222 28224 45228
rect 28276 44724 28304 45562
rect 28368 45404 28396 46922
rect 28460 45558 28488 53944
rect 28644 53582 28672 56200
rect 29288 54194 29316 56200
rect 29932 56114 29960 56200
rect 30024 56114 30052 56222
rect 29932 56086 30052 56114
rect 30104 54324 30156 54330
rect 30104 54266 30156 54272
rect 29276 54188 29328 54194
rect 29276 54130 29328 54136
rect 28816 54120 28868 54126
rect 28816 54062 28868 54068
rect 29736 54120 29788 54126
rect 29736 54062 29788 54068
rect 28632 53576 28684 53582
rect 28632 53518 28684 53524
rect 28632 53440 28684 53446
rect 28632 53382 28684 53388
rect 28644 51074 28672 53382
rect 28552 51046 28672 51074
rect 28552 48618 28580 51046
rect 28540 48612 28592 48618
rect 28540 48554 28592 48560
rect 28552 46986 28580 48554
rect 28632 48272 28684 48278
rect 28632 48214 28684 48220
rect 28644 47258 28672 48214
rect 28724 48204 28776 48210
rect 28724 48146 28776 48152
rect 28632 47252 28684 47258
rect 28632 47194 28684 47200
rect 28540 46980 28592 46986
rect 28540 46922 28592 46928
rect 28644 46918 28672 47194
rect 28632 46912 28684 46918
rect 28538 46880 28594 46889
rect 28632 46854 28684 46860
rect 28538 46815 28594 46824
rect 28552 46646 28580 46815
rect 28540 46640 28592 46646
rect 28540 46582 28592 46588
rect 28632 46640 28684 46646
rect 28632 46582 28684 46588
rect 28644 45626 28672 46582
rect 28632 45620 28684 45626
rect 28632 45562 28684 45568
rect 28448 45552 28500 45558
rect 28448 45494 28500 45500
rect 28632 45484 28684 45490
rect 28632 45426 28684 45432
rect 28368 45376 28580 45404
rect 28448 44872 28500 44878
rect 28448 44814 28500 44820
rect 28276 44696 28396 44724
rect 27950 44636 28258 44645
rect 27950 44634 27956 44636
rect 28012 44634 28036 44636
rect 28092 44634 28116 44636
rect 28172 44634 28196 44636
rect 28252 44634 28258 44636
rect 28012 44582 28014 44634
rect 28194 44582 28196 44634
rect 27950 44580 27956 44582
rect 28012 44580 28036 44582
rect 28092 44580 28116 44582
rect 28172 44580 28196 44582
rect 28252 44580 28258 44582
rect 27950 44571 28258 44580
rect 27804 44464 27856 44470
rect 27804 44406 27856 44412
rect 27724 43812 27844 43840
rect 27712 43716 27764 43722
rect 27712 43658 27764 43664
rect 27540 42906 27660 42922
rect 27528 42900 27660 42906
rect 27580 42894 27660 42900
rect 27528 42842 27580 42848
rect 27436 42764 27488 42770
rect 27436 42706 27488 42712
rect 27344 41744 27396 41750
rect 27344 41686 27396 41692
rect 27344 41608 27396 41614
rect 27344 41550 27396 41556
rect 27356 40594 27384 41550
rect 27344 40588 27396 40594
rect 27344 40530 27396 40536
rect 27448 40118 27476 42706
rect 27528 42560 27580 42566
rect 27528 42502 27580 42508
rect 27436 40112 27488 40118
rect 27436 40054 27488 40060
rect 27344 39976 27396 39982
rect 27342 39944 27344 39953
rect 27396 39944 27398 39953
rect 27342 39879 27398 39888
rect 27252 39296 27304 39302
rect 27252 39238 27304 39244
rect 27356 39137 27384 39879
rect 27434 39264 27490 39273
rect 27434 39199 27490 39208
rect 27342 39128 27398 39137
rect 27342 39063 27398 39072
rect 27252 38956 27304 38962
rect 27252 38898 27304 38904
rect 27160 38344 27212 38350
rect 27160 38286 27212 38292
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 27068 37800 27120 37806
rect 27068 37742 27120 37748
rect 27080 37330 27108 37742
rect 27068 37324 27120 37330
rect 27068 37266 27120 37272
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 26884 30796 26936 30802
rect 26884 30738 26936 30744
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26516 28484 26568 28490
rect 26516 28426 26568 28432
rect 26712 21554 26740 30534
rect 27080 29102 27108 37266
rect 27172 36786 27200 37810
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 27264 35494 27292 38898
rect 27344 38888 27396 38894
rect 27448 38865 27476 39199
rect 27344 38830 27396 38836
rect 27434 38856 27490 38865
rect 27356 38758 27384 38830
rect 27434 38791 27490 38800
rect 27344 38752 27396 38758
rect 27344 38694 27396 38700
rect 27356 37777 27384 38694
rect 27448 38418 27476 38791
rect 27436 38412 27488 38418
rect 27436 38354 27488 38360
rect 27540 38298 27568 42502
rect 27724 41274 27752 43658
rect 27816 42362 27844 43812
rect 27950 43548 28258 43557
rect 27950 43546 27956 43548
rect 28012 43546 28036 43548
rect 28092 43546 28116 43548
rect 28172 43546 28196 43548
rect 28252 43546 28258 43548
rect 28012 43494 28014 43546
rect 28194 43494 28196 43546
rect 27950 43492 27956 43494
rect 28012 43492 28036 43494
rect 28092 43492 28116 43494
rect 28172 43492 28196 43494
rect 28252 43492 28258 43494
rect 27950 43483 28258 43492
rect 28264 43444 28316 43450
rect 28264 43386 28316 43392
rect 28276 42820 28304 43386
rect 28368 42888 28396 44696
rect 28460 43058 28488 44814
rect 28552 44470 28580 45376
rect 28540 44464 28592 44470
rect 28540 44406 28592 44412
rect 28540 44328 28592 44334
rect 28538 44296 28540 44305
rect 28592 44296 28594 44305
rect 28538 44231 28594 44240
rect 28460 43030 28580 43058
rect 28368 42860 28488 42888
rect 28276 42792 28396 42820
rect 27950 42460 28258 42469
rect 27950 42458 27956 42460
rect 28012 42458 28036 42460
rect 28092 42458 28116 42460
rect 28172 42458 28196 42460
rect 28252 42458 28258 42460
rect 28012 42406 28014 42458
rect 28194 42406 28196 42458
rect 27950 42404 27956 42406
rect 28012 42404 28036 42406
rect 28092 42404 28116 42406
rect 28172 42404 28196 42406
rect 28252 42404 28258 42406
rect 27950 42395 28258 42404
rect 27804 42356 27856 42362
rect 27804 42298 27856 42304
rect 27804 41472 27856 41478
rect 27804 41414 27856 41420
rect 27712 41268 27764 41274
rect 27712 41210 27764 41216
rect 27712 41064 27764 41070
rect 27712 41006 27764 41012
rect 27620 39364 27672 39370
rect 27620 39306 27672 39312
rect 27632 39098 27660 39306
rect 27620 39092 27672 39098
rect 27620 39034 27672 39040
rect 27540 38282 27660 38298
rect 27540 38276 27672 38282
rect 27540 38270 27620 38276
rect 27620 38218 27672 38224
rect 27436 38208 27488 38214
rect 27436 38150 27488 38156
rect 27342 37768 27398 37777
rect 27342 37703 27398 37712
rect 27448 36530 27476 38150
rect 27632 37262 27660 38218
rect 27620 37256 27672 37262
rect 27620 37198 27672 37204
rect 27528 37188 27580 37194
rect 27528 37130 27580 37136
rect 27356 36502 27476 36530
rect 27252 35488 27304 35494
rect 27252 35430 27304 35436
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 27172 33522 27200 34546
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 27068 29096 27120 29102
rect 27068 29038 27120 29044
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 26712 18086 26740 21490
rect 26700 18080 26752 18086
rect 26700 18022 26752 18028
rect 27172 16574 27200 33458
rect 27264 33318 27292 35430
rect 27356 34649 27384 36502
rect 27436 36236 27488 36242
rect 27540 36224 27568 37130
rect 27488 36196 27568 36224
rect 27632 36394 27660 37198
rect 27724 36854 27752 41006
rect 27816 40186 27844 41414
rect 27950 41372 28258 41381
rect 27950 41370 27956 41372
rect 28012 41370 28036 41372
rect 28092 41370 28116 41372
rect 28172 41370 28196 41372
rect 28252 41370 28258 41372
rect 28012 41318 28014 41370
rect 28194 41318 28196 41370
rect 27950 41316 27956 41318
rect 28012 41316 28036 41318
rect 28092 41316 28116 41318
rect 28172 41316 28196 41318
rect 28252 41316 28258 41318
rect 27950 41307 28258 41316
rect 28368 41138 28396 42792
rect 28356 41132 28408 41138
rect 28356 41074 28408 41080
rect 28460 41070 28488 42860
rect 28448 41064 28500 41070
rect 28448 41006 28500 41012
rect 28356 40928 28408 40934
rect 28356 40870 28408 40876
rect 27950 40284 28258 40293
rect 27950 40282 27956 40284
rect 28012 40282 28036 40284
rect 28092 40282 28116 40284
rect 28172 40282 28196 40284
rect 28252 40282 28258 40284
rect 28012 40230 28014 40282
rect 28194 40230 28196 40282
rect 27950 40228 27956 40230
rect 28012 40228 28036 40230
rect 28092 40228 28116 40230
rect 28172 40228 28196 40230
rect 28252 40228 28258 40230
rect 27950 40219 28258 40228
rect 27804 40180 27856 40186
rect 27804 40122 27856 40128
rect 27804 39840 27856 39846
rect 27804 39782 27856 39788
rect 27816 39030 27844 39782
rect 27950 39196 28258 39205
rect 27950 39194 27956 39196
rect 28012 39194 28036 39196
rect 28092 39194 28116 39196
rect 28172 39194 28196 39196
rect 28252 39194 28258 39196
rect 28012 39142 28014 39194
rect 28194 39142 28196 39194
rect 27950 39140 27956 39142
rect 28012 39140 28036 39142
rect 28092 39140 28116 39142
rect 28172 39140 28196 39142
rect 28252 39140 28258 39142
rect 27950 39131 28258 39140
rect 27804 39024 27856 39030
rect 27804 38966 27856 38972
rect 27950 38108 28258 38117
rect 27950 38106 27956 38108
rect 28012 38106 28036 38108
rect 28092 38106 28116 38108
rect 28172 38106 28196 38108
rect 28252 38106 28258 38108
rect 28012 38054 28014 38106
rect 28194 38054 28196 38106
rect 27950 38052 27956 38054
rect 28012 38052 28036 38054
rect 28092 38052 28116 38054
rect 28172 38052 28196 38054
rect 28252 38052 28258 38054
rect 27950 38043 28258 38052
rect 28172 37936 28224 37942
rect 28172 37878 28224 37884
rect 28184 37806 28212 37878
rect 28172 37800 28224 37806
rect 28172 37742 28224 37748
rect 28262 37768 28318 37777
rect 28184 37108 28212 37742
rect 28262 37703 28318 37712
rect 28276 37466 28304 37703
rect 28264 37460 28316 37466
rect 28264 37402 28316 37408
rect 28368 37330 28396 40870
rect 28552 40769 28580 43030
rect 28644 40905 28672 45426
rect 28736 45354 28764 48146
rect 28828 47138 28856 54062
rect 29092 53984 29144 53990
rect 29092 53926 29144 53932
rect 29104 51074 29132 53926
rect 29460 53712 29512 53718
rect 29460 53654 29512 53660
rect 29104 51046 29224 51074
rect 28908 50856 28960 50862
rect 28908 50798 28960 50804
rect 29092 50856 29144 50862
rect 29092 50798 29144 50804
rect 28920 48618 28948 50798
rect 29000 49836 29052 49842
rect 29000 49778 29052 49784
rect 29012 49178 29040 49778
rect 29104 49638 29132 50798
rect 29092 49632 29144 49638
rect 29092 49574 29144 49580
rect 29012 49150 29132 49178
rect 29196 49162 29224 51046
rect 29368 49632 29420 49638
rect 29368 49574 29420 49580
rect 29380 49298 29408 49574
rect 29472 49366 29500 53654
rect 29644 53508 29696 53514
rect 29644 53450 29696 53456
rect 29460 49360 29512 49366
rect 29460 49302 29512 49308
rect 29368 49292 29420 49298
rect 29368 49234 29420 49240
rect 29000 49088 29052 49094
rect 29000 49030 29052 49036
rect 28908 48612 28960 48618
rect 28908 48554 28960 48560
rect 29012 47734 29040 49030
rect 29104 48074 29132 49150
rect 29184 49156 29236 49162
rect 29184 49098 29236 49104
rect 29092 48068 29144 48074
rect 29092 48010 29144 48016
rect 29000 47728 29052 47734
rect 29000 47670 29052 47676
rect 29104 47190 29132 48010
rect 29092 47184 29144 47190
rect 28828 47110 28948 47138
rect 29092 47126 29144 47132
rect 28816 47048 28868 47054
rect 28814 47016 28816 47025
rect 28868 47016 28870 47025
rect 28814 46951 28870 46960
rect 28920 46714 28948 47110
rect 29092 46912 29144 46918
rect 29092 46854 29144 46860
rect 28908 46708 28960 46714
rect 28908 46650 28960 46656
rect 28920 46458 28948 46650
rect 29104 46510 29132 46854
rect 29196 46714 29224 49098
rect 29276 48816 29328 48822
rect 29276 48758 29328 48764
rect 29288 48618 29316 48758
rect 29276 48612 29328 48618
rect 29276 48554 29328 48560
rect 29380 47802 29408 49234
rect 29368 47796 29420 47802
rect 29368 47738 29420 47744
rect 29368 47592 29420 47598
rect 29368 47534 29420 47540
rect 29276 47184 29328 47190
rect 29276 47126 29328 47132
rect 29184 46708 29236 46714
rect 29184 46650 29236 46656
rect 29092 46504 29144 46510
rect 28920 46430 29040 46458
rect 29092 46446 29144 46452
rect 28908 46368 28960 46374
rect 28908 46310 28960 46316
rect 28724 45348 28776 45354
rect 28724 45290 28776 45296
rect 28736 45014 28764 45290
rect 28724 45008 28776 45014
rect 28724 44950 28776 44956
rect 28724 44872 28776 44878
rect 28724 44814 28776 44820
rect 28736 44538 28764 44814
rect 28724 44532 28776 44538
rect 28724 44474 28776 44480
rect 28724 44192 28776 44198
rect 28724 44134 28776 44140
rect 28736 41414 28764 44134
rect 28736 41386 28856 41414
rect 28828 41154 28856 41386
rect 28920 41206 28948 46310
rect 29012 46102 29040 46430
rect 29288 46152 29316 47126
rect 29196 46124 29316 46152
rect 29000 46096 29052 46102
rect 29000 46038 29052 46044
rect 29196 45966 29224 46124
rect 29274 46064 29330 46073
rect 29274 45999 29330 46008
rect 29184 45960 29236 45966
rect 29184 45902 29236 45908
rect 29288 45830 29316 45999
rect 29276 45824 29328 45830
rect 29276 45766 29328 45772
rect 29000 45484 29052 45490
rect 29000 45426 29052 45432
rect 29012 44266 29040 45426
rect 29276 45416 29328 45422
rect 29276 45358 29328 45364
rect 29288 45286 29316 45358
rect 29276 45280 29328 45286
rect 29276 45222 29328 45228
rect 29276 45008 29328 45014
rect 29276 44950 29328 44956
rect 29092 44804 29144 44810
rect 29092 44746 29144 44752
rect 29000 44260 29052 44266
rect 29000 44202 29052 44208
rect 29000 41608 29052 41614
rect 29000 41550 29052 41556
rect 29012 41274 29040 41550
rect 29000 41268 29052 41274
rect 29000 41210 29052 41216
rect 28736 41126 28856 41154
rect 28908 41200 28960 41206
rect 28908 41142 28960 41148
rect 28736 40934 28764 41126
rect 28816 41064 28868 41070
rect 28816 41006 28868 41012
rect 28724 40928 28776 40934
rect 28630 40896 28686 40905
rect 28724 40870 28776 40876
rect 28630 40831 28686 40840
rect 28538 40760 28594 40769
rect 28538 40695 28594 40704
rect 28632 40520 28684 40526
rect 28538 40488 28594 40497
rect 28632 40462 28684 40468
rect 28538 40423 28594 40432
rect 28448 38888 28500 38894
rect 28448 38830 28500 38836
rect 28460 38350 28488 38830
rect 28552 38554 28580 40423
rect 28644 39642 28672 40462
rect 28724 40384 28776 40390
rect 28724 40326 28776 40332
rect 28632 39636 28684 39642
rect 28632 39578 28684 39584
rect 28632 39500 28684 39506
rect 28632 39442 28684 39448
rect 28644 39370 28672 39442
rect 28632 39364 28684 39370
rect 28632 39306 28684 39312
rect 28540 38548 28592 38554
rect 28540 38490 28592 38496
rect 28448 38344 28500 38350
rect 28448 38286 28500 38292
rect 28460 38010 28488 38286
rect 28448 38004 28500 38010
rect 28448 37946 28500 37952
rect 28356 37324 28408 37330
rect 28356 37266 28408 37272
rect 28184 37080 28396 37108
rect 27950 37020 28258 37029
rect 27950 37018 27956 37020
rect 28012 37018 28036 37020
rect 28092 37018 28116 37020
rect 28172 37018 28196 37020
rect 28252 37018 28258 37020
rect 28012 36966 28014 37018
rect 28194 36966 28196 37018
rect 27950 36964 27956 36966
rect 28012 36964 28036 36966
rect 28092 36964 28116 36966
rect 28172 36964 28196 36966
rect 28252 36964 28258 36966
rect 27950 36955 28258 36964
rect 27712 36848 27764 36854
rect 28172 36848 28224 36854
rect 27764 36808 27936 36836
rect 27712 36790 27764 36796
rect 27804 36712 27856 36718
rect 27804 36654 27856 36660
rect 27632 36378 27752 36394
rect 27632 36372 27764 36378
rect 27632 36366 27712 36372
rect 27436 36178 27488 36184
rect 27448 34678 27476 36178
rect 27632 36122 27660 36366
rect 27712 36314 27764 36320
rect 27540 36094 27660 36122
rect 27712 36100 27764 36106
rect 27436 34672 27488 34678
rect 27342 34640 27398 34649
rect 27436 34614 27488 34620
rect 27342 34575 27398 34584
rect 27252 33312 27304 33318
rect 27252 33254 27304 33260
rect 27264 32978 27292 33254
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27540 29850 27568 36094
rect 27712 36042 27764 36048
rect 27724 34746 27752 36042
rect 27816 34746 27844 36654
rect 27908 36038 27936 36808
rect 28368 36836 28396 37080
rect 28224 36808 28396 36836
rect 28172 36790 28224 36796
rect 28184 36145 28212 36790
rect 28356 36236 28408 36242
rect 28356 36178 28408 36184
rect 28170 36136 28226 36145
rect 28170 36071 28172 36080
rect 28224 36071 28226 36080
rect 28172 36042 28224 36048
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 27950 35932 28258 35941
rect 27950 35930 27956 35932
rect 28012 35930 28036 35932
rect 28092 35930 28116 35932
rect 28172 35930 28196 35932
rect 28252 35930 28258 35932
rect 28012 35878 28014 35930
rect 28194 35878 28196 35930
rect 27950 35876 27956 35878
rect 28012 35876 28036 35878
rect 28092 35876 28116 35878
rect 28172 35876 28196 35878
rect 28252 35876 28258 35878
rect 27950 35867 28258 35876
rect 27986 35320 28042 35329
rect 27986 35255 28042 35264
rect 28000 35154 28028 35255
rect 27988 35148 28040 35154
rect 27988 35090 28040 35096
rect 28000 35057 28028 35090
rect 27986 35048 28042 35057
rect 27986 34983 28042 34992
rect 27950 34844 28258 34853
rect 27950 34842 27956 34844
rect 28012 34842 28036 34844
rect 28092 34842 28116 34844
rect 28172 34842 28196 34844
rect 28252 34842 28258 34844
rect 28012 34790 28014 34842
rect 28194 34790 28196 34842
rect 27950 34788 27956 34790
rect 28012 34788 28036 34790
rect 28092 34788 28116 34790
rect 28172 34788 28196 34790
rect 28252 34788 28258 34790
rect 27950 34779 28258 34788
rect 27712 34740 27764 34746
rect 27712 34682 27764 34688
rect 27804 34740 27856 34746
rect 27804 34682 27856 34688
rect 27896 34672 27948 34678
rect 27896 34614 27948 34620
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27632 32910 27660 33934
rect 27620 32904 27672 32910
rect 27620 32846 27672 32852
rect 27620 32768 27672 32774
rect 27620 32710 27672 32716
rect 27632 31278 27660 32710
rect 27620 31272 27672 31278
rect 27620 31214 27672 31220
rect 27528 29844 27580 29850
rect 27528 29786 27580 29792
rect 27632 22094 27660 31214
rect 27724 30598 27752 33934
rect 27908 33912 27936 34614
rect 27816 33884 27936 33912
rect 27816 33572 27844 33884
rect 27950 33756 28258 33765
rect 27950 33754 27956 33756
rect 28012 33754 28036 33756
rect 28092 33754 28116 33756
rect 28172 33754 28196 33756
rect 28252 33754 28258 33756
rect 28012 33702 28014 33754
rect 28194 33702 28196 33754
rect 27950 33700 27956 33702
rect 28012 33700 28036 33702
rect 28092 33700 28116 33702
rect 28172 33700 28196 33702
rect 28252 33700 28258 33702
rect 27950 33691 28258 33700
rect 27896 33584 27948 33590
rect 27816 33544 27896 33572
rect 27896 33526 27948 33532
rect 28368 32978 28396 36178
rect 28460 35766 28488 37946
rect 28644 37806 28672 39306
rect 28632 37800 28684 37806
rect 28632 37742 28684 37748
rect 28630 36136 28686 36145
rect 28630 36071 28686 36080
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28448 35760 28500 35766
rect 28448 35702 28500 35708
rect 28552 34762 28580 35974
rect 28644 35766 28672 36071
rect 28632 35760 28684 35766
rect 28632 35702 28684 35708
rect 28460 34734 28580 34762
rect 28356 32972 28408 32978
rect 28356 32914 28408 32920
rect 28460 32858 28488 34734
rect 28632 32972 28684 32978
rect 28632 32914 28684 32920
rect 28368 32830 28488 32858
rect 27950 32668 28258 32677
rect 27950 32666 27956 32668
rect 28012 32666 28036 32668
rect 28092 32666 28116 32668
rect 28172 32666 28196 32668
rect 28252 32666 28258 32668
rect 28012 32614 28014 32666
rect 28194 32614 28196 32666
rect 27950 32612 27956 32614
rect 28012 32612 28036 32614
rect 28092 32612 28116 32614
rect 28172 32612 28196 32614
rect 28252 32612 28258 32614
rect 27950 32603 28258 32612
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 27816 31482 27844 31758
rect 27950 31580 28258 31589
rect 27950 31578 27956 31580
rect 28012 31578 28036 31580
rect 28092 31578 28116 31580
rect 28172 31578 28196 31580
rect 28252 31578 28258 31580
rect 28012 31526 28014 31578
rect 28194 31526 28196 31578
rect 27950 31524 27956 31526
rect 28012 31524 28036 31526
rect 28092 31524 28116 31526
rect 28172 31524 28196 31526
rect 28252 31524 28258 31526
rect 27950 31515 28258 31524
rect 27804 31476 27856 31482
rect 27804 31418 27856 31424
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 27950 30492 28258 30501
rect 27950 30490 27956 30492
rect 28012 30490 28036 30492
rect 28092 30490 28116 30492
rect 28172 30490 28196 30492
rect 28252 30490 28258 30492
rect 28012 30438 28014 30490
rect 28194 30438 28196 30490
rect 27950 30436 27956 30438
rect 28012 30436 28036 30438
rect 28092 30436 28116 30438
rect 28172 30436 28196 30438
rect 28252 30436 28258 30438
rect 27950 30427 28258 30436
rect 27950 29404 28258 29413
rect 27950 29402 27956 29404
rect 28012 29402 28036 29404
rect 28092 29402 28116 29404
rect 28172 29402 28196 29404
rect 28252 29402 28258 29404
rect 28012 29350 28014 29402
rect 28194 29350 28196 29402
rect 27950 29348 27956 29350
rect 28012 29348 28036 29350
rect 28092 29348 28116 29350
rect 28172 29348 28196 29350
rect 28252 29348 28258 29350
rect 27950 29339 28258 29348
rect 27950 28316 28258 28325
rect 27950 28314 27956 28316
rect 28012 28314 28036 28316
rect 28092 28314 28116 28316
rect 28172 28314 28196 28316
rect 28252 28314 28258 28316
rect 28012 28262 28014 28314
rect 28194 28262 28196 28314
rect 27950 28260 27956 28262
rect 28012 28260 28036 28262
rect 28092 28260 28116 28262
rect 28172 28260 28196 28262
rect 28252 28260 28258 28262
rect 27950 28251 28258 28260
rect 28368 27402 28396 32830
rect 28540 32768 28592 32774
rect 28540 32710 28592 32716
rect 28552 32502 28580 32710
rect 28540 32496 28592 32502
rect 28540 32438 28592 32444
rect 28540 32224 28592 32230
rect 28460 32184 28540 32212
rect 28460 28762 28488 32184
rect 28540 32166 28592 32172
rect 28644 29714 28672 32914
rect 28736 32230 28764 40326
rect 28828 38010 28856 41006
rect 29000 40996 29052 41002
rect 29000 40938 29052 40944
rect 28906 40896 28962 40905
rect 28906 40831 28962 40840
rect 28920 39846 28948 40831
rect 29012 40633 29040 40938
rect 29104 40730 29132 44746
rect 29184 44260 29236 44266
rect 29184 44202 29236 44208
rect 29196 42566 29224 44202
rect 29288 42906 29316 44950
rect 29380 43858 29408 47534
rect 29472 46714 29500 49302
rect 29552 48748 29604 48754
rect 29552 48690 29604 48696
rect 29460 46708 29512 46714
rect 29460 46650 29512 46656
rect 29460 46028 29512 46034
rect 29460 45970 29512 45976
rect 29368 43852 29420 43858
rect 29368 43794 29420 43800
rect 29472 43314 29500 45970
rect 29564 43994 29592 48690
rect 29656 45558 29684 53450
rect 29644 45552 29696 45558
rect 29644 45494 29696 45500
rect 29552 43988 29604 43994
rect 29552 43930 29604 43936
rect 29460 43308 29512 43314
rect 29460 43250 29512 43256
rect 29368 43240 29420 43246
rect 29368 43182 29420 43188
rect 29276 42900 29328 42906
rect 29276 42842 29328 42848
rect 29184 42560 29236 42566
rect 29184 42502 29236 42508
rect 29196 41750 29224 42502
rect 29276 42152 29328 42158
rect 29276 42094 29328 42100
rect 29184 41744 29236 41750
rect 29184 41686 29236 41692
rect 29184 40996 29236 41002
rect 29184 40938 29236 40944
rect 29092 40724 29144 40730
rect 29092 40666 29144 40672
rect 28998 40624 29054 40633
rect 28998 40559 29054 40568
rect 28908 39840 28960 39846
rect 29196 39817 29224 40938
rect 28908 39782 28960 39788
rect 29182 39808 29238 39817
rect 29182 39743 29238 39752
rect 28906 39672 28962 39681
rect 28906 39607 28962 39616
rect 29092 39636 29144 39642
rect 28920 39522 28948 39607
rect 29092 39578 29144 39584
rect 28920 39506 28994 39522
rect 28920 39500 29006 39506
rect 28920 39494 28954 39500
rect 28954 39442 29006 39448
rect 28908 39364 28960 39370
rect 28908 39306 28960 39312
rect 28816 38004 28868 38010
rect 28816 37946 28868 37952
rect 28828 36310 28856 37946
rect 28816 36304 28868 36310
rect 28816 36246 28868 36252
rect 28814 34640 28870 34649
rect 28814 34575 28870 34584
rect 28828 34542 28856 34575
rect 28816 34536 28868 34542
rect 28816 34478 28868 34484
rect 28920 34202 28948 39306
rect 29104 35630 29132 39578
rect 29288 38978 29316 42094
rect 29380 40594 29408 43182
rect 29472 42770 29500 43250
rect 29460 42764 29512 42770
rect 29460 42706 29512 42712
rect 29472 41682 29500 42706
rect 29656 42362 29684 45494
rect 29748 45490 29776 54062
rect 30012 50448 30064 50454
rect 30012 50390 30064 50396
rect 30024 48226 30052 50390
rect 30116 49434 30144 54266
rect 30196 54256 30248 54262
rect 30196 54198 30248 54204
rect 30208 49858 30236 54198
rect 30300 54194 30328 56222
rect 30562 56200 30618 57000
rect 31206 56200 31262 57000
rect 31850 56200 31906 57000
rect 32494 56200 32550 57000
rect 33138 56200 33194 57000
rect 33782 56200 33838 57000
rect 34426 56200 34482 57000
rect 35070 56200 35126 57000
rect 35714 56200 35770 57000
rect 36358 56200 36414 57000
rect 37002 56200 37058 57000
rect 37646 56200 37702 57000
rect 38290 56200 38346 57000
rect 38934 56200 38990 57000
rect 39578 56200 39634 57000
rect 40222 56200 40278 57000
rect 42154 56200 42210 57000
rect 42798 56200 42854 57000
rect 43442 56200 43498 57000
rect 44086 56200 44142 57000
rect 44730 56200 44786 57000
rect 45374 56200 45430 57000
rect 46018 56200 46074 57000
rect 46662 56200 46718 57000
rect 47306 56200 47362 57000
rect 47950 56200 48006 57000
rect 48594 56200 48650 57000
rect 49238 56200 49294 57000
rect 30576 55214 30604 56200
rect 30576 55186 30696 55214
rect 30564 54664 30616 54670
rect 30564 54606 30616 54612
rect 30288 54188 30340 54194
rect 30288 54130 30340 54136
rect 30380 53984 30432 53990
rect 30380 53926 30432 53932
rect 30392 50726 30420 53926
rect 30472 53440 30524 53446
rect 30472 53382 30524 53388
rect 30380 50720 30432 50726
rect 30380 50662 30432 50668
rect 30288 50176 30340 50182
rect 30484 50130 30512 53382
rect 30576 51074 30604 54606
rect 30668 54194 30696 55186
rect 30656 54188 30708 54194
rect 30656 54130 30708 54136
rect 30748 53984 30800 53990
rect 30748 53926 30800 53932
rect 30576 51046 30696 51074
rect 30564 50720 30616 50726
rect 30564 50662 30616 50668
rect 30576 50318 30604 50662
rect 30564 50312 30616 50318
rect 30564 50254 30616 50260
rect 30340 50124 30512 50130
rect 30288 50118 30512 50124
rect 30300 50102 30512 50118
rect 30208 49830 30328 49858
rect 30196 49768 30248 49774
rect 30196 49710 30248 49716
rect 30104 49428 30156 49434
rect 30104 49370 30156 49376
rect 30116 49162 30144 49370
rect 30104 49156 30156 49162
rect 30104 49098 30156 49104
rect 29932 48198 30052 48226
rect 29828 47184 29880 47190
rect 29828 47126 29880 47132
rect 29736 45484 29788 45490
rect 29736 45426 29788 45432
rect 29736 45280 29788 45286
rect 29736 45222 29788 45228
rect 29644 42356 29696 42362
rect 29644 42298 29696 42304
rect 29552 42220 29604 42226
rect 29552 42162 29604 42168
rect 29460 41676 29512 41682
rect 29460 41618 29512 41624
rect 29564 41478 29592 42162
rect 29644 42084 29696 42090
rect 29644 42026 29696 42032
rect 29552 41472 29604 41478
rect 29552 41414 29604 41420
rect 29656 40594 29684 42026
rect 29748 41274 29776 45222
rect 29736 41268 29788 41274
rect 29736 41210 29788 41216
rect 29736 40928 29788 40934
rect 29736 40870 29788 40876
rect 29368 40588 29420 40594
rect 29368 40530 29420 40536
rect 29644 40588 29696 40594
rect 29644 40530 29696 40536
rect 29748 40338 29776 40870
rect 29840 40662 29868 47126
rect 29932 47122 29960 48198
rect 30012 48136 30064 48142
rect 30012 48078 30064 48084
rect 29920 47116 29972 47122
rect 29920 47058 29972 47064
rect 30024 46578 30052 48078
rect 30208 47462 30236 49710
rect 30300 48618 30328 49830
rect 30392 49094 30420 50102
rect 30472 49904 30524 49910
rect 30472 49846 30524 49852
rect 30380 49088 30432 49094
rect 30380 49030 30432 49036
rect 30288 48612 30340 48618
rect 30288 48554 30340 48560
rect 30196 47456 30248 47462
rect 30116 47416 30196 47444
rect 30012 46572 30064 46578
rect 30012 46514 30064 46520
rect 29920 46164 29972 46170
rect 29920 46106 29972 46112
rect 29932 45966 29960 46106
rect 30024 46034 30052 46514
rect 30012 46028 30064 46034
rect 30012 45970 30064 45976
rect 29920 45960 29972 45966
rect 29920 45902 29972 45908
rect 30116 45354 30144 47416
rect 30196 47398 30248 47404
rect 30196 47116 30248 47122
rect 30196 47058 30248 47064
rect 30208 46034 30236 47058
rect 30300 46986 30328 48554
rect 30484 47054 30512 49846
rect 30472 47048 30524 47054
rect 30472 46990 30524 46996
rect 30576 46986 30604 50254
rect 30668 50250 30696 51046
rect 30656 50244 30708 50250
rect 30656 50186 30708 50192
rect 30668 49722 30696 50186
rect 30760 49910 30788 53926
rect 31220 53582 31248 56200
rect 31864 54194 31892 56200
rect 32508 55214 32536 56200
rect 33152 55214 33180 56200
rect 32508 55186 32628 55214
rect 33152 55186 33272 55214
rect 32496 54596 32548 54602
rect 32496 54538 32548 54544
rect 32220 54324 32272 54330
rect 32220 54266 32272 54272
rect 31852 54188 31904 54194
rect 31852 54130 31904 54136
rect 31944 54052 31996 54058
rect 31944 53994 31996 54000
rect 31208 53576 31260 53582
rect 31208 53518 31260 53524
rect 31760 53440 31812 53446
rect 31760 53382 31812 53388
rect 31772 51074 31800 53382
rect 31772 51046 31892 51074
rect 31300 50924 31352 50930
rect 31300 50866 31352 50872
rect 31024 50720 31076 50726
rect 31024 50662 31076 50668
rect 30748 49904 30800 49910
rect 30748 49846 30800 49852
rect 30668 49694 30880 49722
rect 30656 48680 30708 48686
rect 30656 48622 30708 48628
rect 30668 48210 30696 48622
rect 30748 48544 30800 48550
rect 30748 48486 30800 48492
rect 30656 48204 30708 48210
rect 30656 48146 30708 48152
rect 30288 46980 30340 46986
rect 30288 46922 30340 46928
rect 30564 46980 30616 46986
rect 30564 46922 30616 46928
rect 30288 46368 30340 46374
rect 30288 46310 30340 46316
rect 30472 46368 30524 46374
rect 30472 46310 30524 46316
rect 30196 46028 30248 46034
rect 30196 45970 30248 45976
rect 30104 45348 30156 45354
rect 30104 45290 30156 45296
rect 30104 44396 30156 44402
rect 30104 44338 30156 44344
rect 30012 44328 30064 44334
rect 30116 44305 30144 44338
rect 30012 44270 30064 44276
rect 30102 44296 30158 44305
rect 30024 44146 30052 44270
rect 30102 44231 30158 44240
rect 30024 44118 30144 44146
rect 30012 43852 30064 43858
rect 30012 43794 30064 43800
rect 29828 40656 29880 40662
rect 29828 40598 29880 40604
rect 29656 40310 29776 40338
rect 29288 38950 29408 38978
rect 29184 38888 29236 38894
rect 29184 38830 29236 38836
rect 29276 38888 29328 38894
rect 29276 38830 29328 38836
rect 29196 36310 29224 38830
rect 29184 36304 29236 36310
rect 29184 36246 29236 36252
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 29104 35290 29132 35566
rect 29092 35284 29144 35290
rect 29092 35226 29144 35232
rect 29196 35154 29224 36246
rect 29288 35222 29316 38830
rect 29276 35216 29328 35222
rect 29276 35158 29328 35164
rect 29184 35148 29236 35154
rect 29184 35090 29236 35096
rect 29380 34406 29408 38950
rect 29656 38486 29684 40310
rect 29736 40180 29788 40186
rect 29736 40122 29788 40128
rect 29748 38842 29776 40122
rect 30024 39642 30052 43794
rect 30116 41818 30144 44118
rect 30104 41812 30156 41818
rect 30104 41754 30156 41760
rect 30104 40384 30156 40390
rect 30104 40326 30156 40332
rect 30012 39636 30064 39642
rect 30012 39578 30064 39584
rect 29828 39432 29880 39438
rect 29828 39374 29880 39380
rect 29840 38962 29868 39374
rect 29920 39296 29972 39302
rect 29920 39238 29972 39244
rect 29828 38956 29880 38962
rect 29828 38898 29880 38904
rect 29748 38814 29868 38842
rect 29644 38480 29696 38486
rect 29644 38422 29696 38428
rect 29642 35320 29698 35329
rect 29642 35255 29698 35264
rect 29460 34944 29512 34950
rect 29460 34886 29512 34892
rect 29368 34400 29420 34406
rect 29288 34360 29368 34388
rect 28908 34196 28960 34202
rect 28908 34138 28960 34144
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 28724 32224 28776 32230
rect 28724 32166 28776 32172
rect 28736 31890 28764 32166
rect 28724 31884 28776 31890
rect 28724 31826 28776 31832
rect 28724 31680 28776 31686
rect 28724 31622 28776 31628
rect 28736 30666 28764 31622
rect 28724 30660 28776 30666
rect 28724 30602 28776 30608
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 28448 28756 28500 28762
rect 28448 28698 28500 28704
rect 28356 27396 28408 27402
rect 28356 27338 28408 27344
rect 27950 27228 28258 27237
rect 27950 27226 27956 27228
rect 28012 27226 28036 27228
rect 28092 27226 28116 27228
rect 28172 27226 28196 27228
rect 28252 27226 28258 27228
rect 28012 27174 28014 27226
rect 28194 27174 28196 27226
rect 27950 27172 27956 27174
rect 28012 27172 28036 27174
rect 28092 27172 28116 27174
rect 28172 27172 28196 27174
rect 28252 27172 28258 27174
rect 27950 27163 28258 27172
rect 27950 26140 28258 26149
rect 27950 26138 27956 26140
rect 28012 26138 28036 26140
rect 28092 26138 28116 26140
rect 28172 26138 28196 26140
rect 28252 26138 28258 26140
rect 28012 26086 28014 26138
rect 28194 26086 28196 26138
rect 27950 26084 27956 26086
rect 28012 26084 28036 26086
rect 28092 26084 28116 26086
rect 28172 26084 28196 26086
rect 28252 26084 28258 26086
rect 27950 26075 28258 26084
rect 27950 25052 28258 25061
rect 27950 25050 27956 25052
rect 28012 25050 28036 25052
rect 28092 25050 28116 25052
rect 28172 25050 28196 25052
rect 28252 25050 28258 25052
rect 28012 24998 28014 25050
rect 28194 24998 28196 25050
rect 27950 24996 27956 24998
rect 28012 24996 28036 24998
rect 28092 24996 28116 24998
rect 28172 24996 28196 24998
rect 28252 24996 28258 24998
rect 27950 24987 28258 24996
rect 28460 24818 28488 28698
rect 28448 24812 28500 24818
rect 28448 24754 28500 24760
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 28736 22094 28764 30602
rect 28828 29306 28856 33934
rect 29184 32904 29236 32910
rect 29184 32846 29236 32852
rect 29092 32360 29144 32366
rect 29092 32302 29144 32308
rect 28906 31920 28962 31929
rect 29104 31890 29132 32302
rect 28906 31855 28908 31864
rect 28960 31855 28962 31864
rect 29092 31884 29144 31890
rect 28908 31826 28960 31832
rect 29092 31826 29144 31832
rect 29000 31816 29052 31822
rect 28920 31764 29000 31770
rect 28920 31758 29052 31764
rect 28920 31742 29040 31758
rect 28816 29300 28868 29306
rect 28816 29242 28868 29248
rect 28920 29170 28948 31742
rect 29196 31482 29224 32846
rect 29288 32366 29316 34360
rect 29368 34342 29420 34348
rect 29276 32360 29328 32366
rect 29276 32302 29328 32308
rect 29184 31476 29236 31482
rect 29184 31418 29236 31424
rect 29288 31278 29316 32302
rect 29472 31958 29500 34886
rect 29552 33924 29604 33930
rect 29552 33866 29604 33872
rect 29564 33522 29592 33866
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 29460 31952 29512 31958
rect 29460 31894 29512 31900
rect 29276 31272 29328 31278
rect 29276 31214 29328 31220
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 29104 29306 29132 29990
rect 29184 29504 29236 29510
rect 29184 29446 29236 29452
rect 29092 29300 29144 29306
rect 29092 29242 29144 29248
rect 28908 29164 28960 29170
rect 28908 29106 28960 29112
rect 29196 29102 29224 29446
rect 29184 29096 29236 29102
rect 29184 29038 29236 29044
rect 27632 22066 27752 22094
rect 27724 17202 27752 22066
rect 28644 22066 28764 22094
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 27080 16546 27200 16574
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 25872 3460 25924 3466
rect 25872 3402 25924 3408
rect 25412 2508 25464 2514
rect 25412 2450 25464 2456
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 25424 800 25452 2450
rect 26252 2378 26280 15438
rect 26608 11076 26660 11082
rect 26608 11018 26660 11024
rect 26620 5710 26648 11018
rect 27080 10130 27108 16546
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 27160 14340 27212 14346
rect 27160 14282 27212 14288
rect 27172 12442 27200 14282
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27160 12436 27212 12442
rect 27160 12378 27212 12384
rect 27528 12300 27580 12306
rect 27528 12242 27580 12248
rect 27068 10124 27120 10130
rect 27068 10066 27120 10072
rect 27540 8378 27568 12242
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27804 9920 27856 9926
rect 27804 9862 27856 9868
rect 27816 8430 27844 9862
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27804 8424 27856 8430
rect 27540 8350 27660 8378
rect 27804 8366 27856 8372
rect 27632 8294 27660 8350
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28368 2582 28396 14894
rect 28644 13938 28672 22066
rect 29196 17678 29224 29038
rect 29656 25974 29684 35255
rect 29840 34406 29868 38814
rect 29932 38758 29960 39238
rect 29920 38752 29972 38758
rect 29920 38694 29972 38700
rect 29920 37936 29972 37942
rect 29920 37878 29972 37884
rect 29932 37262 29960 37878
rect 30012 37324 30064 37330
rect 30012 37266 30064 37272
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 29932 36854 29960 37198
rect 29920 36848 29972 36854
rect 29920 36790 29972 36796
rect 29932 36242 29960 36790
rect 29920 36236 29972 36242
rect 29920 36178 29972 36184
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29828 34400 29880 34406
rect 29828 34342 29880 34348
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29748 32910 29776 33458
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29748 31890 29776 32846
rect 29736 31884 29788 31890
rect 29736 31826 29788 31832
rect 29840 31278 29868 34342
rect 29932 33538 29960 34546
rect 30024 34066 30052 37266
rect 30116 36582 30144 40326
rect 30208 39982 30236 45970
rect 30300 45422 30328 46310
rect 30288 45416 30340 45422
rect 30288 45358 30340 45364
rect 30380 45416 30432 45422
rect 30380 45358 30432 45364
rect 30300 44198 30328 45358
rect 30392 44538 30420 45358
rect 30380 44532 30432 44538
rect 30380 44474 30432 44480
rect 30484 44470 30512 46310
rect 30656 46164 30708 46170
rect 30656 46106 30708 46112
rect 30564 45484 30616 45490
rect 30564 45426 30616 45432
rect 30472 44464 30524 44470
rect 30472 44406 30524 44412
rect 30288 44192 30340 44198
rect 30288 44134 30340 44140
rect 30576 42906 30604 45426
rect 30668 43738 30696 46106
rect 30760 44538 30788 48486
rect 30852 48314 30880 49694
rect 31036 49162 31064 50662
rect 31116 50176 31168 50182
rect 31116 50118 31168 50124
rect 31024 49156 31076 49162
rect 31024 49098 31076 49104
rect 30852 48286 30972 48314
rect 30944 47410 30972 48286
rect 31024 48204 31076 48210
rect 31024 48146 31076 48152
rect 31036 47598 31064 48146
rect 31024 47592 31076 47598
rect 31024 47534 31076 47540
rect 30944 47382 31064 47410
rect 30932 47252 30984 47258
rect 30932 47194 30984 47200
rect 30840 46504 30892 46510
rect 30840 46446 30892 46452
rect 30852 46034 30880 46446
rect 30840 46028 30892 46034
rect 30840 45970 30892 45976
rect 30840 44736 30892 44742
rect 30840 44678 30892 44684
rect 30748 44532 30800 44538
rect 30748 44474 30800 44480
rect 30852 44266 30880 44678
rect 30840 44260 30892 44266
rect 30840 44202 30892 44208
rect 30944 43790 30972 47194
rect 31036 47122 31064 47382
rect 31024 47116 31076 47122
rect 31024 47058 31076 47064
rect 31024 46096 31076 46102
rect 31024 46038 31076 46044
rect 30932 43784 30984 43790
rect 30668 43710 30880 43738
rect 30932 43726 30984 43732
rect 31036 43722 31064 46038
rect 31128 45354 31156 50118
rect 31208 48680 31260 48686
rect 31208 48622 31260 48628
rect 31116 45348 31168 45354
rect 31116 45290 31168 45296
rect 31220 45082 31248 48622
rect 31312 48226 31340 50866
rect 31576 50720 31628 50726
rect 31576 50662 31628 50668
rect 31588 49858 31616 50662
rect 31668 50244 31720 50250
rect 31668 50186 31720 50192
rect 31680 49978 31708 50186
rect 31668 49972 31720 49978
rect 31668 49914 31720 49920
rect 31588 49830 31708 49858
rect 31680 49774 31708 49830
rect 31576 49768 31628 49774
rect 31576 49710 31628 49716
rect 31668 49768 31720 49774
rect 31668 49710 31720 49716
rect 31312 48210 31432 48226
rect 31312 48204 31444 48210
rect 31312 48198 31392 48204
rect 31392 48146 31444 48152
rect 31300 48068 31352 48074
rect 31300 48010 31352 48016
rect 31312 47734 31340 48010
rect 31300 47728 31352 47734
rect 31300 47670 31352 47676
rect 31312 46646 31340 47670
rect 31484 47116 31536 47122
rect 31484 47058 31536 47064
rect 31300 46640 31352 46646
rect 31300 46582 31352 46588
rect 31496 45914 31524 47058
rect 31588 46918 31616 49710
rect 31760 49224 31812 49230
rect 31760 49166 31812 49172
rect 31772 47802 31800 49166
rect 31864 48890 31892 51046
rect 31956 49842 31984 53994
rect 31944 49836 31996 49842
rect 31944 49778 31996 49784
rect 32036 49156 32088 49162
rect 32036 49098 32088 49104
rect 32048 48890 32076 49098
rect 31852 48884 31904 48890
rect 31852 48826 31904 48832
rect 32036 48884 32088 48890
rect 32036 48826 32088 48832
rect 31852 48748 31904 48754
rect 31852 48690 31904 48696
rect 31760 47796 31812 47802
rect 31760 47738 31812 47744
rect 31864 47530 31892 48690
rect 31944 47796 31996 47802
rect 31944 47738 31996 47744
rect 31760 47524 31812 47530
rect 31760 47466 31812 47472
rect 31852 47524 31904 47530
rect 31852 47466 31904 47472
rect 31576 46912 31628 46918
rect 31576 46854 31628 46860
rect 31668 46640 31720 46646
rect 31668 46582 31720 46588
rect 31576 46028 31628 46034
rect 31576 45970 31628 45976
rect 31588 45914 31616 45970
rect 31680 45966 31708 46582
rect 31772 46510 31800 47466
rect 31852 46572 31904 46578
rect 31852 46514 31904 46520
rect 31760 46504 31812 46510
rect 31760 46446 31812 46452
rect 31300 45892 31352 45898
rect 31300 45834 31352 45840
rect 31496 45886 31616 45914
rect 31668 45960 31720 45966
rect 31668 45902 31720 45908
rect 31312 45354 31340 45834
rect 31300 45348 31352 45354
rect 31300 45290 31352 45296
rect 31496 45234 31524 45886
rect 31864 45554 31892 46514
rect 31404 45206 31524 45234
rect 31680 45526 31892 45554
rect 31208 45076 31260 45082
rect 31208 45018 31260 45024
rect 31208 44736 31260 44742
rect 31208 44678 31260 44684
rect 30748 43648 30800 43654
rect 30748 43590 30800 43596
rect 30852 43602 30880 43710
rect 31024 43716 31076 43722
rect 31024 43658 31076 43664
rect 30564 42900 30616 42906
rect 30564 42842 30616 42848
rect 30380 41676 30432 41682
rect 30300 41636 30380 41664
rect 30300 40594 30328 41636
rect 30380 41618 30432 41624
rect 30656 41676 30708 41682
rect 30656 41618 30708 41624
rect 30288 40588 30340 40594
rect 30288 40530 30340 40536
rect 30564 40520 30616 40526
rect 30564 40462 30616 40468
rect 30196 39976 30248 39982
rect 30196 39918 30248 39924
rect 30208 39098 30236 39918
rect 30196 39092 30248 39098
rect 30196 39034 30248 39040
rect 30378 38312 30434 38321
rect 30378 38247 30434 38256
rect 30392 37126 30420 38247
rect 30472 37188 30524 37194
rect 30472 37130 30524 37136
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30484 36718 30512 37130
rect 30288 36712 30340 36718
rect 30288 36654 30340 36660
rect 30472 36712 30524 36718
rect 30472 36654 30524 36660
rect 30104 36576 30156 36582
rect 30104 36518 30156 36524
rect 30300 36242 30328 36654
rect 30288 36236 30340 36242
rect 30288 36178 30340 36184
rect 30196 35624 30248 35630
rect 30196 35566 30248 35572
rect 30012 34060 30064 34066
rect 30012 34002 30064 34008
rect 30104 33856 30156 33862
rect 30104 33798 30156 33804
rect 30010 33552 30066 33561
rect 29932 33510 30010 33538
rect 30010 33487 30012 33496
rect 30064 33487 30066 33496
rect 30012 33458 30064 33464
rect 30116 32978 30144 33798
rect 30104 32972 30156 32978
rect 30104 32914 30156 32920
rect 30104 32224 30156 32230
rect 30104 32166 30156 32172
rect 30116 32026 30144 32166
rect 30104 32020 30156 32026
rect 30104 31962 30156 31968
rect 30012 31884 30064 31890
rect 30012 31826 30064 31832
rect 30024 31754 30052 31826
rect 30012 31748 30064 31754
rect 30012 31690 30064 31696
rect 29828 31272 29880 31278
rect 29828 31214 29880 31220
rect 30208 30938 30236 35566
rect 30300 35562 30328 36178
rect 30380 35760 30432 35766
rect 30380 35702 30432 35708
rect 30288 35556 30340 35562
rect 30288 35498 30340 35504
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 30300 35154 30328 35226
rect 30288 35148 30340 35154
rect 30288 35090 30340 35096
rect 30392 35018 30420 35702
rect 30380 35012 30432 35018
rect 30380 34954 30432 34960
rect 30380 34740 30432 34746
rect 30380 34682 30432 34688
rect 30286 32872 30342 32881
rect 30286 32807 30288 32816
rect 30340 32807 30342 32816
rect 30288 32778 30340 32784
rect 30392 32366 30420 34682
rect 30472 33312 30524 33318
rect 30472 33254 30524 33260
rect 30484 32978 30512 33254
rect 30472 32972 30524 32978
rect 30472 32914 30524 32920
rect 30484 32842 30512 32914
rect 30472 32836 30524 32842
rect 30472 32778 30524 32784
rect 30484 32434 30512 32778
rect 30576 32570 30604 40462
rect 30668 40118 30696 41618
rect 30656 40112 30708 40118
rect 30656 40054 30708 40060
rect 30668 38962 30696 40054
rect 30656 38956 30708 38962
rect 30656 38898 30708 38904
rect 30760 36922 30788 43590
rect 30852 43574 30972 43602
rect 30840 42900 30892 42906
rect 30840 42842 30892 42848
rect 30852 41274 30880 42842
rect 30840 41268 30892 41274
rect 30840 41210 30892 41216
rect 30840 41064 30892 41070
rect 30840 41006 30892 41012
rect 30748 36916 30800 36922
rect 30748 36858 30800 36864
rect 30852 33862 30880 41006
rect 30944 40526 30972 43574
rect 31116 43104 31168 43110
rect 31116 43046 31168 43052
rect 31024 41064 31076 41070
rect 31024 41006 31076 41012
rect 30932 40520 30984 40526
rect 30932 40462 30984 40468
rect 30932 39024 30984 39030
rect 31036 39012 31064 41006
rect 31128 40050 31156 43046
rect 31220 42401 31248 44678
rect 31300 43988 31352 43994
rect 31300 43930 31352 43936
rect 31312 43110 31340 43930
rect 31300 43104 31352 43110
rect 31300 43046 31352 43052
rect 31206 42392 31262 42401
rect 31206 42327 31262 42336
rect 31300 42084 31352 42090
rect 31300 42026 31352 42032
rect 31206 41032 31262 41041
rect 31206 40967 31262 40976
rect 31116 40044 31168 40050
rect 31116 39986 31168 39992
rect 30984 38984 31064 39012
rect 31220 39001 31248 40967
rect 31312 39098 31340 42026
rect 31404 41070 31432 45206
rect 31576 44940 31628 44946
rect 31576 44882 31628 44888
rect 31588 43722 31616 44882
rect 31576 43716 31628 43722
rect 31576 43658 31628 43664
rect 31588 43450 31616 43658
rect 31576 43444 31628 43450
rect 31576 43386 31628 43392
rect 31574 43344 31630 43353
rect 31574 43279 31630 43288
rect 31484 42900 31536 42906
rect 31484 42842 31536 42848
rect 31496 42362 31524 42842
rect 31484 42356 31536 42362
rect 31484 42298 31536 42304
rect 31496 41818 31524 42298
rect 31484 41812 31536 41818
rect 31484 41754 31536 41760
rect 31392 41064 31444 41070
rect 31392 41006 31444 41012
rect 31392 40928 31444 40934
rect 31392 40870 31444 40876
rect 31300 39092 31352 39098
rect 31300 39034 31352 39040
rect 31206 38992 31262 39001
rect 30932 38966 30984 38972
rect 30944 38010 30972 38966
rect 31206 38927 31262 38936
rect 30932 38004 30984 38010
rect 30932 37946 30984 37952
rect 31116 37664 31168 37670
rect 31116 37606 31168 37612
rect 31128 37466 31156 37606
rect 31116 37460 31168 37466
rect 31116 37402 31168 37408
rect 30930 37360 30986 37369
rect 30930 37295 30932 37304
rect 30984 37295 30986 37304
rect 30932 37266 30984 37272
rect 31220 37233 31248 38927
rect 31300 38276 31352 38282
rect 31300 38218 31352 38224
rect 31312 37942 31340 38218
rect 31300 37936 31352 37942
rect 31300 37878 31352 37884
rect 31312 37466 31340 37878
rect 31300 37460 31352 37466
rect 31300 37402 31352 37408
rect 31206 37224 31262 37233
rect 31206 37159 31262 37168
rect 31312 36854 31340 37402
rect 31300 36848 31352 36854
rect 31300 36790 31352 36796
rect 31312 36106 31340 36790
rect 31300 36100 31352 36106
rect 31300 36042 31352 36048
rect 31024 36032 31076 36038
rect 31024 35974 31076 35980
rect 31208 36032 31260 36038
rect 31208 35974 31260 35980
rect 31036 35630 31064 35974
rect 31024 35624 31076 35630
rect 31024 35566 31076 35572
rect 31116 35556 31168 35562
rect 31116 35498 31168 35504
rect 31128 35290 31156 35498
rect 31116 35284 31168 35290
rect 31116 35226 31168 35232
rect 31024 35216 31076 35222
rect 31220 35170 31248 35974
rect 31076 35164 31248 35170
rect 31024 35158 31248 35164
rect 31036 35142 31248 35158
rect 31208 34672 31260 34678
rect 31312 34660 31340 36042
rect 31260 34632 31340 34660
rect 31208 34614 31260 34620
rect 31116 34060 31168 34066
rect 31116 34002 31168 34008
rect 30840 33856 30892 33862
rect 30840 33798 30892 33804
rect 31024 33856 31076 33862
rect 31024 33798 31076 33804
rect 30748 33584 30800 33590
rect 30748 33526 30800 33532
rect 30760 33318 30788 33526
rect 30852 33318 30880 33798
rect 30748 33312 30800 33318
rect 30748 33254 30800 33260
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30564 32564 30616 32570
rect 30564 32506 30616 32512
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30852 31210 30880 32370
rect 30840 31204 30892 31210
rect 30840 31146 30892 31152
rect 30196 30932 30248 30938
rect 30196 30874 30248 30880
rect 31036 30394 31064 33798
rect 31128 33658 31156 34002
rect 31220 33658 31248 34614
rect 31116 33652 31168 33658
rect 31116 33594 31168 33600
rect 31208 33652 31260 33658
rect 31208 33594 31260 33600
rect 31128 31958 31156 33594
rect 31220 32978 31248 33594
rect 31300 33040 31352 33046
rect 31300 32982 31352 32988
rect 31208 32972 31260 32978
rect 31208 32914 31260 32920
rect 31116 31952 31168 31958
rect 31116 31894 31168 31900
rect 31220 31890 31248 32914
rect 31312 32881 31340 32982
rect 31298 32872 31354 32881
rect 31298 32807 31354 32816
rect 31300 32496 31352 32502
rect 31300 32438 31352 32444
rect 31208 31884 31260 31890
rect 31208 31826 31260 31832
rect 31312 31822 31340 32438
rect 31404 31890 31432 40870
rect 31484 40588 31536 40594
rect 31484 40530 31536 40536
rect 31496 40186 31524 40530
rect 31484 40180 31536 40186
rect 31484 40122 31536 40128
rect 31588 39982 31616 43279
rect 31680 42634 31708 45526
rect 31760 44940 31812 44946
rect 31760 44882 31812 44888
rect 31668 42628 31720 42634
rect 31668 42570 31720 42576
rect 31680 42362 31708 42570
rect 31668 42356 31720 42362
rect 31668 42298 31720 42304
rect 31576 39976 31628 39982
rect 31576 39918 31628 39924
rect 31576 39024 31628 39030
rect 31576 38966 31628 38972
rect 31588 38282 31616 38966
rect 31576 38276 31628 38282
rect 31576 38218 31628 38224
rect 31484 38208 31536 38214
rect 31484 38150 31536 38156
rect 31496 35630 31524 38150
rect 31680 36224 31708 42298
rect 31772 41414 31800 44882
rect 31956 43858 31984 47738
rect 32048 45422 32076 48826
rect 32126 48240 32182 48249
rect 32126 48175 32182 48184
rect 32140 48142 32168 48175
rect 32128 48136 32180 48142
rect 32128 48078 32180 48084
rect 32140 47734 32168 48078
rect 32128 47728 32180 47734
rect 32128 47670 32180 47676
rect 32128 47524 32180 47530
rect 32128 47466 32180 47472
rect 32036 45416 32088 45422
rect 32036 45358 32088 45364
rect 32140 44402 32168 47466
rect 32232 44402 32260 54266
rect 32312 53984 32364 53990
rect 32312 53926 32364 53932
rect 32324 50930 32352 53926
rect 32508 51074 32536 54538
rect 32600 54194 32628 55186
rect 33244 54194 33272 55186
rect 33692 54256 33744 54262
rect 33692 54198 33744 54204
rect 32588 54188 32640 54194
rect 32588 54130 32640 54136
rect 33232 54188 33284 54194
rect 33232 54130 33284 54136
rect 33704 53990 33732 54198
rect 32588 53984 32640 53990
rect 32588 53926 32640 53932
rect 33600 53984 33652 53990
rect 33600 53926 33652 53932
rect 33692 53984 33744 53990
rect 33692 53926 33744 53932
rect 32416 51046 32536 51074
rect 32312 50924 32364 50930
rect 32312 50866 32364 50872
rect 32324 50522 32352 50866
rect 32312 50516 32364 50522
rect 32312 50458 32364 50464
rect 32312 48680 32364 48686
rect 32312 48622 32364 48628
rect 32324 48346 32352 48622
rect 32312 48340 32364 48346
rect 32312 48282 32364 48288
rect 32312 46368 32364 46374
rect 32312 46310 32364 46316
rect 32324 45626 32352 46310
rect 32312 45620 32364 45626
rect 32312 45562 32364 45568
rect 32128 44396 32180 44402
rect 32128 44338 32180 44344
rect 32220 44396 32272 44402
rect 32220 44338 32272 44344
rect 32232 44010 32260 44338
rect 32416 44334 32444 51046
rect 32600 49978 32628 53926
rect 32950 53884 33258 53893
rect 32950 53882 32956 53884
rect 33012 53882 33036 53884
rect 33092 53882 33116 53884
rect 33172 53882 33196 53884
rect 33252 53882 33258 53884
rect 33012 53830 33014 53882
rect 33194 53830 33196 53882
rect 32950 53828 32956 53830
rect 33012 53828 33036 53830
rect 33092 53828 33116 53830
rect 33172 53828 33196 53830
rect 33252 53828 33258 53830
rect 32950 53819 33258 53828
rect 32950 52796 33258 52805
rect 32950 52794 32956 52796
rect 33012 52794 33036 52796
rect 33092 52794 33116 52796
rect 33172 52794 33196 52796
rect 33252 52794 33258 52796
rect 33012 52742 33014 52794
rect 33194 52742 33196 52794
rect 32950 52740 32956 52742
rect 33012 52740 33036 52742
rect 33092 52740 33116 52742
rect 33172 52740 33196 52742
rect 33252 52740 33258 52742
rect 32950 52731 33258 52740
rect 32950 51708 33258 51717
rect 32950 51706 32956 51708
rect 33012 51706 33036 51708
rect 33092 51706 33116 51708
rect 33172 51706 33196 51708
rect 33252 51706 33258 51708
rect 33012 51654 33014 51706
rect 33194 51654 33196 51706
rect 32950 51652 32956 51654
rect 33012 51652 33036 51654
rect 33092 51652 33116 51654
rect 33172 51652 33196 51654
rect 33252 51652 33258 51654
rect 32950 51643 33258 51652
rect 32950 50620 33258 50629
rect 32950 50618 32956 50620
rect 33012 50618 33036 50620
rect 33092 50618 33116 50620
rect 33172 50618 33196 50620
rect 33252 50618 33258 50620
rect 33012 50566 33014 50618
rect 33194 50566 33196 50618
rect 32950 50564 32956 50566
rect 33012 50564 33036 50566
rect 33092 50564 33116 50566
rect 33172 50564 33196 50566
rect 33252 50564 33258 50566
rect 32950 50555 33258 50564
rect 32956 50516 33008 50522
rect 32956 50458 33008 50464
rect 32588 49972 32640 49978
rect 32588 49914 32640 49920
rect 32772 49972 32824 49978
rect 32772 49914 32824 49920
rect 32864 49972 32916 49978
rect 32864 49914 32916 49920
rect 32588 49836 32640 49842
rect 32588 49778 32640 49784
rect 32680 49836 32732 49842
rect 32680 49778 32732 49784
rect 32496 49632 32548 49638
rect 32496 49574 32548 49580
rect 32508 46578 32536 49574
rect 32600 47122 32628 49778
rect 32692 48074 32720 49778
rect 32784 48113 32812 49914
rect 32770 48104 32826 48113
rect 32680 48068 32732 48074
rect 32770 48039 32826 48048
rect 32680 48010 32732 48016
rect 32772 48000 32824 48006
rect 32772 47942 32824 47948
rect 32784 47530 32812 47942
rect 32772 47524 32824 47530
rect 32772 47466 32824 47472
rect 32588 47116 32640 47122
rect 32588 47058 32640 47064
rect 32680 47116 32732 47122
rect 32680 47058 32732 47064
rect 32588 46708 32640 46714
rect 32588 46650 32640 46656
rect 32496 46572 32548 46578
rect 32496 46514 32548 46520
rect 32600 46374 32628 46650
rect 32588 46368 32640 46374
rect 32588 46310 32640 46316
rect 32496 45960 32548 45966
rect 32496 45902 32548 45908
rect 32508 45558 32536 45902
rect 32496 45552 32548 45558
rect 32496 45494 32548 45500
rect 32692 44946 32720 47058
rect 32772 46504 32824 46510
rect 32772 46446 32824 46452
rect 32784 46170 32812 46446
rect 32772 46164 32824 46170
rect 32772 46106 32824 46112
rect 32876 45558 32904 49914
rect 32968 49842 32996 50458
rect 33508 50380 33560 50386
rect 33508 50322 33560 50328
rect 32956 49836 33008 49842
rect 32956 49778 33008 49784
rect 32950 49532 33258 49541
rect 32950 49530 32956 49532
rect 33012 49530 33036 49532
rect 33092 49530 33116 49532
rect 33172 49530 33196 49532
rect 33252 49530 33258 49532
rect 33012 49478 33014 49530
rect 33194 49478 33196 49530
rect 32950 49476 32956 49478
rect 33012 49476 33036 49478
rect 33092 49476 33116 49478
rect 33172 49476 33196 49478
rect 33252 49476 33258 49478
rect 32950 49467 33258 49476
rect 33520 49434 33548 50322
rect 33612 49910 33640 53926
rect 33796 53582 33824 56200
rect 34440 53650 34468 56200
rect 34520 54528 34572 54534
rect 34520 54470 34572 54476
rect 34428 53644 34480 53650
rect 34428 53586 34480 53592
rect 33784 53576 33836 53582
rect 33784 53518 33836 53524
rect 33692 53032 33744 53038
rect 33692 52974 33744 52980
rect 33600 49904 33652 49910
rect 33600 49846 33652 49852
rect 33508 49428 33560 49434
rect 33508 49370 33560 49376
rect 33324 49360 33376 49366
rect 33324 49302 33376 49308
rect 33336 49230 33364 49302
rect 33324 49224 33376 49230
rect 33324 49166 33376 49172
rect 33416 49088 33468 49094
rect 33416 49030 33468 49036
rect 33428 48890 33456 49030
rect 33048 48884 33100 48890
rect 33048 48826 33100 48832
rect 33416 48884 33468 48890
rect 33416 48826 33468 48832
rect 33060 48686 33088 48826
rect 33048 48680 33100 48686
rect 33048 48622 33100 48628
rect 32950 48444 33258 48453
rect 32950 48442 32956 48444
rect 33012 48442 33036 48444
rect 33092 48442 33116 48444
rect 33172 48442 33196 48444
rect 33252 48442 33258 48444
rect 33012 48390 33014 48442
rect 33194 48390 33196 48442
rect 32950 48388 32956 48390
rect 33012 48388 33036 48390
rect 33092 48388 33116 48390
rect 33172 48388 33196 48390
rect 33252 48388 33258 48390
rect 32950 48379 33258 48388
rect 33416 48000 33468 48006
rect 33416 47942 33468 47948
rect 32950 47356 33258 47365
rect 32950 47354 32956 47356
rect 33012 47354 33036 47356
rect 33092 47354 33116 47356
rect 33172 47354 33196 47356
rect 33252 47354 33258 47356
rect 33012 47302 33014 47354
rect 33194 47302 33196 47354
rect 32950 47300 32956 47302
rect 33012 47300 33036 47302
rect 33092 47300 33116 47302
rect 33172 47300 33196 47302
rect 33252 47300 33258 47302
rect 32950 47291 33258 47300
rect 33324 46912 33376 46918
rect 33324 46854 33376 46860
rect 32950 46268 33258 46277
rect 32950 46266 32956 46268
rect 33012 46266 33036 46268
rect 33092 46266 33116 46268
rect 33172 46266 33196 46268
rect 33252 46266 33258 46268
rect 33012 46214 33014 46266
rect 33194 46214 33196 46266
rect 32950 46212 32956 46214
rect 33012 46212 33036 46214
rect 33092 46212 33116 46214
rect 33172 46212 33196 46214
rect 33252 46212 33258 46214
rect 32950 46203 33258 46212
rect 32956 45892 33008 45898
rect 33232 45892 33284 45898
rect 33008 45852 33232 45880
rect 32956 45834 33008 45840
rect 33232 45834 33284 45840
rect 32864 45552 32916 45558
rect 32864 45494 32916 45500
rect 33232 45552 33284 45558
rect 33232 45494 33284 45500
rect 32772 45416 32824 45422
rect 32772 45358 32824 45364
rect 32680 44940 32732 44946
rect 32680 44882 32732 44888
rect 32496 44736 32548 44742
rect 32496 44678 32548 44684
rect 32404 44328 32456 44334
rect 32404 44270 32456 44276
rect 32140 43982 32260 44010
rect 31944 43852 31996 43858
rect 31944 43794 31996 43800
rect 31956 43314 31984 43794
rect 31944 43308 31996 43314
rect 31944 43250 31996 43256
rect 31956 42770 31984 43250
rect 31944 42764 31996 42770
rect 31944 42706 31996 42712
rect 31852 42288 31904 42294
rect 31852 42230 31904 42236
rect 31864 41546 31892 42230
rect 31956 42158 31984 42706
rect 31944 42152 31996 42158
rect 31944 42094 31996 42100
rect 31956 41682 31984 42094
rect 31944 41676 31996 41682
rect 31944 41618 31996 41624
rect 31852 41540 31904 41546
rect 31852 41482 31904 41488
rect 32140 41414 32168 43982
rect 32220 43852 32272 43858
rect 32220 43794 32272 43800
rect 31772 41386 31892 41414
rect 31760 40384 31812 40390
rect 31760 40326 31812 40332
rect 31772 40118 31800 40326
rect 31760 40112 31812 40118
rect 31760 40054 31812 40060
rect 31758 39672 31814 39681
rect 31758 39607 31760 39616
rect 31812 39607 31814 39616
rect 31864 39624 31892 41386
rect 32048 41386 32168 41414
rect 31944 39636 31996 39642
rect 31760 39578 31812 39584
rect 31864 39596 31944 39624
rect 31760 39296 31812 39302
rect 31760 39238 31812 39244
rect 31772 39098 31800 39238
rect 31760 39092 31812 39098
rect 31760 39034 31812 39040
rect 31864 39030 31892 39596
rect 31944 39578 31996 39584
rect 31942 39128 31998 39137
rect 31942 39063 31998 39072
rect 31852 39024 31904 39030
rect 31852 38966 31904 38972
rect 31956 38842 31984 39063
rect 31772 38814 31984 38842
rect 31772 37097 31800 38814
rect 31944 38412 31996 38418
rect 31944 38354 31996 38360
rect 31852 37800 31904 37806
rect 31852 37742 31904 37748
rect 31758 37088 31814 37097
rect 31758 37023 31814 37032
rect 31588 36196 31708 36224
rect 31588 35766 31616 36196
rect 31576 35760 31628 35766
rect 31576 35702 31628 35708
rect 31484 35624 31536 35630
rect 31484 35566 31536 35572
rect 31484 34944 31536 34950
rect 31484 34886 31536 34892
rect 31392 31884 31444 31890
rect 31392 31826 31444 31832
rect 31300 31816 31352 31822
rect 31300 31758 31352 31764
rect 31496 31414 31524 34886
rect 31668 34536 31720 34542
rect 31668 34478 31720 34484
rect 31576 34468 31628 34474
rect 31576 34410 31628 34416
rect 31588 33114 31616 34410
rect 31680 33454 31708 34478
rect 31668 33448 31720 33454
rect 31668 33390 31720 33396
rect 31576 33108 31628 33114
rect 31576 33050 31628 33056
rect 31680 32502 31708 33390
rect 31668 32496 31720 32502
rect 31668 32438 31720 32444
rect 31484 31408 31536 31414
rect 31484 31350 31536 31356
rect 31024 30388 31076 30394
rect 31024 30330 31076 30336
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 30024 29646 30052 30194
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28644 8838 28672 13874
rect 29196 13870 29224 17614
rect 30380 14476 30432 14482
rect 30380 14418 30432 14424
rect 29828 14408 29880 14414
rect 30392 14385 30420 14418
rect 29828 14350 29880 14356
rect 30378 14376 30434 14385
rect 29184 13864 29236 13870
rect 29184 13806 29236 13812
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28816 5636 28868 5642
rect 28816 5578 28868 5584
rect 28828 3058 28856 5578
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 26240 2372 26292 2378
rect 26240 2314 26292 2320
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28736 800 28764 2926
rect 29840 2514 29868 14350
rect 30378 14311 30434 14320
rect 31036 13326 31064 30330
rect 31772 28150 31800 37023
rect 31864 36310 31892 37742
rect 31852 36304 31904 36310
rect 31852 36246 31904 36252
rect 31852 32836 31904 32842
rect 31852 32778 31904 32784
rect 31864 32026 31892 32778
rect 31956 32230 31984 38354
rect 32048 37874 32076 41386
rect 32126 41304 32182 41313
rect 32126 41239 32182 41248
rect 32140 38554 32168 41239
rect 32232 39137 32260 43794
rect 32404 42560 32456 42566
rect 32404 42502 32456 42508
rect 32312 41472 32364 41478
rect 32312 41414 32364 41420
rect 32324 40168 32352 41414
rect 32416 40526 32444 42502
rect 32508 41313 32536 44678
rect 32680 44396 32732 44402
rect 32680 44338 32732 44344
rect 32588 44328 32640 44334
rect 32588 44270 32640 44276
rect 32600 43858 32628 44270
rect 32692 43926 32720 44338
rect 32680 43920 32732 43926
rect 32680 43862 32732 43868
rect 32588 43852 32640 43858
rect 32588 43794 32640 43800
rect 32588 43648 32640 43654
rect 32588 43590 32640 43596
rect 32600 41818 32628 43590
rect 32784 42770 32812 45358
rect 33244 45354 33272 45494
rect 33232 45348 33284 45354
rect 33232 45290 33284 45296
rect 32950 45180 33258 45189
rect 32950 45178 32956 45180
rect 33012 45178 33036 45180
rect 33092 45178 33116 45180
rect 33172 45178 33196 45180
rect 33252 45178 33258 45180
rect 33012 45126 33014 45178
rect 33194 45126 33196 45178
rect 32950 45124 32956 45126
rect 33012 45124 33036 45126
rect 33092 45124 33116 45126
rect 33172 45124 33196 45126
rect 33252 45124 33258 45126
rect 32950 45115 33258 45124
rect 33138 44976 33194 44985
rect 33138 44911 33140 44920
rect 33192 44911 33194 44920
rect 33140 44882 33192 44888
rect 33336 44810 33364 46854
rect 33428 45626 33456 47942
rect 33520 47734 33548 49370
rect 33600 49224 33652 49230
rect 33600 49166 33652 49172
rect 33508 47728 33560 47734
rect 33508 47670 33560 47676
rect 33416 45620 33468 45626
rect 33416 45562 33468 45568
rect 33508 45416 33560 45422
rect 33508 45358 33560 45364
rect 33416 44940 33468 44946
rect 33416 44882 33468 44888
rect 33324 44804 33376 44810
rect 33324 44746 33376 44752
rect 33324 44328 33376 44334
rect 33324 44270 33376 44276
rect 32950 44092 33258 44101
rect 32950 44090 32956 44092
rect 33012 44090 33036 44092
rect 33092 44090 33116 44092
rect 33172 44090 33196 44092
rect 33252 44090 33258 44092
rect 33012 44038 33014 44090
rect 33194 44038 33196 44090
rect 32950 44036 32956 44038
rect 33012 44036 33036 44038
rect 33092 44036 33116 44038
rect 33172 44036 33196 44038
rect 33252 44036 33258 44038
rect 32950 44027 33258 44036
rect 33048 43852 33100 43858
rect 33048 43794 33100 43800
rect 32864 43716 32916 43722
rect 32864 43658 32916 43664
rect 32876 43382 32904 43658
rect 32864 43376 32916 43382
rect 32864 43318 32916 43324
rect 32772 42764 32824 42770
rect 32772 42706 32824 42712
rect 32784 42294 32812 42706
rect 32876 42634 32904 43318
rect 33060 43246 33088 43794
rect 33232 43716 33284 43722
rect 33232 43658 33284 43664
rect 33244 43450 33272 43658
rect 33232 43444 33284 43450
rect 33232 43386 33284 43392
rect 33048 43240 33100 43246
rect 33048 43182 33100 43188
rect 32950 43004 33258 43013
rect 32950 43002 32956 43004
rect 33012 43002 33036 43004
rect 33092 43002 33116 43004
rect 33172 43002 33196 43004
rect 33252 43002 33258 43004
rect 33012 42950 33014 43002
rect 33194 42950 33196 43002
rect 32950 42948 32956 42950
rect 33012 42948 33036 42950
rect 33092 42948 33116 42950
rect 33172 42948 33196 42950
rect 33252 42948 33258 42950
rect 32950 42939 33258 42948
rect 32864 42628 32916 42634
rect 32864 42570 32916 42576
rect 32876 42362 32904 42570
rect 32864 42356 32916 42362
rect 32864 42298 32916 42304
rect 32772 42288 32824 42294
rect 32772 42230 32824 42236
rect 32588 41812 32640 41818
rect 32588 41754 32640 41760
rect 32784 41414 32812 42230
rect 32864 42152 32916 42158
rect 32864 42094 32916 42100
rect 32692 41386 32812 41414
rect 32494 41304 32550 41313
rect 32494 41239 32550 41248
rect 32496 41132 32548 41138
rect 32496 41074 32548 41080
rect 32508 41041 32536 41074
rect 32494 41032 32550 41041
rect 32494 40967 32550 40976
rect 32508 40934 32536 40967
rect 32496 40928 32548 40934
rect 32496 40870 32548 40876
rect 32404 40520 32456 40526
rect 32404 40462 32456 40468
rect 32324 40140 32444 40168
rect 32312 40044 32364 40050
rect 32312 39986 32364 39992
rect 32324 39506 32352 39986
rect 32312 39500 32364 39506
rect 32312 39442 32364 39448
rect 32312 39296 32364 39302
rect 32312 39238 32364 39244
rect 32218 39128 32274 39137
rect 32218 39063 32274 39072
rect 32220 38956 32272 38962
rect 32220 38898 32272 38904
rect 32128 38548 32180 38554
rect 32128 38490 32180 38496
rect 32232 38350 32260 38898
rect 32220 38344 32272 38350
rect 32220 38286 32272 38292
rect 32036 37868 32088 37874
rect 32036 37810 32088 37816
rect 32324 37262 32352 39238
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32416 37210 32444 40140
rect 32494 39808 32550 39817
rect 32494 39743 32550 39752
rect 32508 38026 32536 39743
rect 32692 38894 32720 41386
rect 32876 40594 32904 42094
rect 32950 41916 33258 41925
rect 32950 41914 32956 41916
rect 33012 41914 33036 41916
rect 33092 41914 33116 41916
rect 33172 41914 33196 41916
rect 33252 41914 33258 41916
rect 33012 41862 33014 41914
rect 33194 41862 33196 41914
rect 32950 41860 32956 41862
rect 33012 41860 33036 41862
rect 33092 41860 33116 41862
rect 33172 41860 33196 41862
rect 33252 41860 33258 41862
rect 32950 41851 33258 41860
rect 32956 41812 33008 41818
rect 32956 41754 33008 41760
rect 32968 41070 32996 41754
rect 33336 41414 33364 44270
rect 33428 41818 33456 44882
rect 33520 44334 33548 45358
rect 33612 45014 33640 49166
rect 33704 47054 33732 52974
rect 34532 50250 34560 54470
rect 35084 54194 35112 56200
rect 35256 54256 35308 54262
rect 35256 54198 35308 54204
rect 35072 54188 35124 54194
rect 35072 54130 35124 54136
rect 35164 50992 35216 50998
rect 35164 50934 35216 50940
rect 34520 50244 34572 50250
rect 34520 50186 34572 50192
rect 34428 50176 34480 50182
rect 34428 50118 34480 50124
rect 34060 49768 34112 49774
rect 34244 49768 34296 49774
rect 34112 49728 34244 49756
rect 34060 49710 34112 49716
rect 34244 49710 34296 49716
rect 34440 49434 34468 50118
rect 34532 49978 34560 50186
rect 35176 49978 35204 50934
rect 35268 50454 35296 54198
rect 35728 54176 35756 56200
rect 35900 54188 35952 54194
rect 35728 54148 35900 54176
rect 35900 54130 35952 54136
rect 36372 53582 36400 56200
rect 37016 54194 37044 56200
rect 37660 55214 37688 56200
rect 38304 55214 38332 56200
rect 37660 55186 37780 55214
rect 38304 55186 38424 55214
rect 37464 54664 37516 54670
rect 37464 54606 37516 54612
rect 37188 54256 37240 54262
rect 37188 54198 37240 54204
rect 37004 54188 37056 54194
rect 37004 54130 37056 54136
rect 36360 53576 36412 53582
rect 36360 53518 36412 53524
rect 36360 52556 36412 52562
rect 36360 52498 36412 52504
rect 35532 52420 35584 52426
rect 35532 52362 35584 52368
rect 35544 51074 35572 52362
rect 35452 51046 35572 51074
rect 36372 51074 36400 52498
rect 37200 51074 37228 54198
rect 37476 53990 37504 54606
rect 37752 54194 37780 55186
rect 37950 54428 38258 54437
rect 37950 54426 37956 54428
rect 38012 54426 38036 54428
rect 38092 54426 38116 54428
rect 38172 54426 38196 54428
rect 38252 54426 38258 54428
rect 38012 54374 38014 54426
rect 38194 54374 38196 54426
rect 37950 54372 37956 54374
rect 38012 54372 38036 54374
rect 38092 54372 38116 54374
rect 38172 54372 38196 54374
rect 38252 54372 38258 54374
rect 37950 54363 38258 54372
rect 38396 54194 38424 55186
rect 37740 54188 37792 54194
rect 37740 54130 37792 54136
rect 38384 54188 38436 54194
rect 38384 54130 38436 54136
rect 37464 53984 37516 53990
rect 37464 53926 37516 53932
rect 37556 53984 37608 53990
rect 37556 53926 37608 53932
rect 37372 53508 37424 53514
rect 37372 53450 37424 53456
rect 37280 51400 37332 51406
rect 37280 51342 37332 51348
rect 36372 51046 36492 51074
rect 35256 50448 35308 50454
rect 35256 50390 35308 50396
rect 34520 49972 34572 49978
rect 34520 49914 34572 49920
rect 35164 49972 35216 49978
rect 35164 49914 35216 49920
rect 34428 49428 34480 49434
rect 34428 49370 34480 49376
rect 34152 49292 34204 49298
rect 34152 49234 34204 49240
rect 33784 49156 33836 49162
rect 33784 49098 33836 49104
rect 33796 48754 33824 49098
rect 33784 48748 33836 48754
rect 33784 48690 33836 48696
rect 33796 48249 33824 48690
rect 34164 48686 34192 49234
rect 34704 49224 34756 49230
rect 34704 49166 34756 49172
rect 34152 48680 34204 48686
rect 34152 48622 34204 48628
rect 34336 48680 34388 48686
rect 34336 48622 34388 48628
rect 33968 48544 34020 48550
rect 33968 48486 34020 48492
rect 33782 48240 33838 48249
rect 33782 48175 33838 48184
rect 33796 47734 33824 48175
rect 33784 47728 33836 47734
rect 33784 47670 33836 47676
rect 33876 47116 33928 47122
rect 33876 47058 33928 47064
rect 33692 47048 33744 47054
rect 33692 46990 33744 46996
rect 33704 46714 33732 46990
rect 33692 46708 33744 46714
rect 33692 46650 33744 46656
rect 33600 45008 33652 45014
rect 33600 44950 33652 44956
rect 33508 44328 33560 44334
rect 33508 44270 33560 44276
rect 33600 44192 33652 44198
rect 33506 44160 33562 44169
rect 33600 44134 33652 44140
rect 33692 44192 33744 44198
rect 33692 44134 33744 44140
rect 33506 44095 33562 44104
rect 33520 43654 33548 44095
rect 33508 43648 33560 43654
rect 33508 43590 33560 43596
rect 33612 42770 33640 44134
rect 33704 43858 33732 44134
rect 33692 43852 33744 43858
rect 33692 43794 33744 43800
rect 33784 43852 33836 43858
rect 33784 43794 33836 43800
rect 33600 42764 33652 42770
rect 33600 42706 33652 42712
rect 33796 42566 33824 43794
rect 33600 42560 33652 42566
rect 33600 42502 33652 42508
rect 33692 42560 33744 42566
rect 33692 42502 33744 42508
rect 33784 42560 33836 42566
rect 33784 42502 33836 42508
rect 33416 41812 33468 41818
rect 33468 41772 33548 41800
rect 33416 41754 33468 41760
rect 33336 41386 33456 41414
rect 33428 41274 33456 41386
rect 33416 41268 33468 41274
rect 33416 41210 33468 41216
rect 33324 41132 33376 41138
rect 33324 41074 33376 41080
rect 32956 41064 33008 41070
rect 32956 41006 33008 41012
rect 32950 40828 33258 40837
rect 32950 40826 32956 40828
rect 33012 40826 33036 40828
rect 33092 40826 33116 40828
rect 33172 40826 33196 40828
rect 33252 40826 33258 40828
rect 33012 40774 33014 40826
rect 33194 40774 33196 40826
rect 32950 40772 32956 40774
rect 33012 40772 33036 40774
rect 33092 40772 33116 40774
rect 33172 40772 33196 40774
rect 33252 40772 33258 40774
rect 32950 40763 33258 40772
rect 33336 40594 33364 41074
rect 32864 40588 32916 40594
rect 32864 40530 32916 40536
rect 33324 40588 33376 40594
rect 33324 40530 33376 40536
rect 32772 40520 32824 40526
rect 32772 40462 32824 40468
rect 32784 39794 32812 40462
rect 32876 40118 32904 40530
rect 32864 40112 32916 40118
rect 32864 40054 32916 40060
rect 33414 40080 33470 40089
rect 33414 40015 33470 40024
rect 32784 39766 32904 39794
rect 32770 39672 32826 39681
rect 32770 39607 32826 39616
rect 32784 39574 32812 39607
rect 32772 39568 32824 39574
rect 32772 39510 32824 39516
rect 32680 38888 32732 38894
rect 32680 38830 32732 38836
rect 32508 37998 32628 38026
rect 32416 37182 32536 37210
rect 32508 37126 32536 37182
rect 32312 37120 32364 37126
rect 32496 37120 32548 37126
rect 32364 37080 32444 37108
rect 32312 37062 32364 37068
rect 32416 36718 32444 37080
rect 32496 37062 32548 37068
rect 32404 36712 32456 36718
rect 32456 36672 32536 36700
rect 32404 36654 32456 36660
rect 32220 36576 32272 36582
rect 32220 36518 32272 36524
rect 32036 35828 32088 35834
rect 32036 35770 32088 35776
rect 32048 35086 32076 35770
rect 32232 35766 32260 36518
rect 32312 36372 32364 36378
rect 32312 36314 32364 36320
rect 32324 36174 32352 36314
rect 32312 36168 32364 36174
rect 32312 36110 32364 36116
rect 32324 35766 32352 36110
rect 32220 35760 32272 35766
rect 32220 35702 32272 35708
rect 32312 35760 32364 35766
rect 32312 35702 32364 35708
rect 32508 35630 32536 36672
rect 32496 35624 32548 35630
rect 32496 35566 32548 35572
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 32220 34944 32272 34950
rect 32220 34886 32272 34892
rect 32128 34604 32180 34610
rect 32128 34546 32180 34552
rect 32140 34354 32168 34546
rect 32232 34542 32260 34886
rect 32220 34536 32272 34542
rect 32220 34478 32272 34484
rect 32140 34326 32260 34354
rect 32128 32768 32180 32774
rect 32128 32710 32180 32716
rect 32036 32292 32088 32298
rect 32036 32234 32088 32240
rect 31944 32224 31996 32230
rect 31944 32166 31996 32172
rect 31852 32020 31904 32026
rect 31852 31962 31904 31968
rect 31760 28144 31812 28150
rect 31760 28086 31812 28092
rect 32048 23730 32076 32234
rect 32140 31958 32168 32710
rect 32128 31952 32180 31958
rect 32128 31894 32180 31900
rect 32036 23724 32088 23730
rect 32036 23666 32088 23672
rect 32232 20874 32260 34326
rect 32402 34096 32458 34105
rect 32402 34031 32404 34040
rect 32456 34031 32458 34040
rect 32404 34002 32456 34008
rect 32508 33998 32536 35566
rect 32600 35154 32628 37998
rect 32772 37188 32824 37194
rect 32772 37130 32824 37136
rect 32680 36916 32732 36922
rect 32680 36858 32732 36864
rect 32692 36106 32720 36858
rect 32784 36718 32812 37130
rect 32772 36712 32824 36718
rect 32772 36654 32824 36660
rect 32876 36394 32904 39766
rect 32950 39740 33258 39749
rect 32950 39738 32956 39740
rect 33012 39738 33036 39740
rect 33092 39738 33116 39740
rect 33172 39738 33196 39740
rect 33252 39738 33258 39740
rect 33012 39686 33014 39738
rect 33194 39686 33196 39738
rect 32950 39684 32956 39686
rect 33012 39684 33036 39686
rect 33092 39684 33116 39686
rect 33172 39684 33196 39686
rect 33252 39684 33258 39686
rect 32950 39675 33258 39684
rect 33140 39432 33192 39438
rect 33140 39374 33192 39380
rect 33152 38826 33180 39374
rect 33428 39370 33456 40015
rect 33520 39964 33548 41772
rect 33612 40066 33640 42502
rect 33704 40458 33732 42502
rect 33692 40452 33744 40458
rect 33692 40394 33744 40400
rect 33612 40038 33732 40066
rect 33600 39976 33652 39982
rect 33520 39936 33600 39964
rect 33600 39918 33652 39924
rect 33704 39506 33732 40038
rect 33692 39500 33744 39506
rect 33692 39442 33744 39448
rect 33416 39364 33468 39370
rect 33416 39306 33468 39312
rect 33600 39296 33652 39302
rect 33600 39238 33652 39244
rect 33612 39098 33640 39238
rect 33600 39092 33652 39098
rect 33600 39034 33652 39040
rect 33600 38956 33652 38962
rect 33600 38898 33652 38904
rect 33140 38820 33192 38826
rect 33140 38762 33192 38768
rect 32950 38652 33258 38661
rect 32950 38650 32956 38652
rect 33012 38650 33036 38652
rect 33092 38650 33116 38652
rect 33172 38650 33196 38652
rect 33252 38650 33258 38652
rect 33012 38598 33014 38650
rect 33194 38598 33196 38650
rect 32950 38596 32956 38598
rect 33012 38596 33036 38598
rect 33092 38596 33116 38598
rect 33172 38596 33196 38598
rect 33252 38596 33258 38598
rect 32950 38587 33258 38596
rect 33416 38208 33468 38214
rect 33416 38150 33468 38156
rect 32950 37564 33258 37573
rect 32950 37562 32956 37564
rect 33012 37562 33036 37564
rect 33092 37562 33116 37564
rect 33172 37562 33196 37564
rect 33252 37562 33258 37564
rect 33012 37510 33014 37562
rect 33194 37510 33196 37562
rect 32950 37508 32956 37510
rect 33012 37508 33036 37510
rect 33092 37508 33116 37510
rect 33172 37508 33196 37510
rect 33252 37508 33258 37510
rect 32950 37499 33258 37508
rect 33428 37466 33456 38150
rect 33416 37460 33468 37466
rect 33416 37402 33468 37408
rect 33324 37324 33376 37330
rect 33324 37266 33376 37272
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 33152 36718 33180 37198
rect 33140 36712 33192 36718
rect 33140 36654 33192 36660
rect 32950 36476 33258 36485
rect 32950 36474 32956 36476
rect 33012 36474 33036 36476
rect 33092 36474 33116 36476
rect 33172 36474 33196 36476
rect 33252 36474 33258 36476
rect 33012 36422 33014 36474
rect 33194 36422 33196 36474
rect 32950 36420 32956 36422
rect 33012 36420 33036 36422
rect 33092 36420 33116 36422
rect 33172 36420 33196 36422
rect 33252 36420 33258 36422
rect 32950 36411 33258 36420
rect 32784 36366 32904 36394
rect 32680 36100 32732 36106
rect 32680 36042 32732 36048
rect 32588 35148 32640 35154
rect 32588 35090 32640 35096
rect 32784 34762 32812 36366
rect 32864 36304 32916 36310
rect 32864 36246 32916 36252
rect 32876 35154 32904 36246
rect 32950 35388 33258 35397
rect 32950 35386 32956 35388
rect 33012 35386 33036 35388
rect 33092 35386 33116 35388
rect 33172 35386 33196 35388
rect 33252 35386 33258 35388
rect 33012 35334 33014 35386
rect 33194 35334 33196 35386
rect 32950 35332 32956 35334
rect 33012 35332 33036 35334
rect 33092 35332 33116 35334
rect 33172 35332 33196 35334
rect 33252 35332 33258 35334
rect 32950 35323 33258 35332
rect 32864 35148 32916 35154
rect 32864 35090 32916 35096
rect 32692 34734 32812 34762
rect 32864 34740 32916 34746
rect 32588 34468 32640 34474
rect 32588 34410 32640 34416
rect 32496 33992 32548 33998
rect 32496 33934 32548 33940
rect 32404 33924 32456 33930
rect 32404 33866 32456 33872
rect 32416 33522 32444 33866
rect 32508 33561 32536 33934
rect 32494 33552 32550 33561
rect 32404 33516 32456 33522
rect 32494 33487 32550 33496
rect 32404 33458 32456 33464
rect 32312 31680 32364 31686
rect 32312 31622 32364 31628
rect 32324 29578 32352 31622
rect 32312 29572 32364 29578
rect 32312 29514 32364 29520
rect 32404 29232 32456 29238
rect 32404 29174 32456 29180
rect 32220 20868 32272 20874
rect 32220 20810 32272 20816
rect 32416 19378 32444 29174
rect 32508 22094 32536 33487
rect 32600 33454 32628 34410
rect 32588 33448 32640 33454
rect 32588 33390 32640 33396
rect 32600 32978 32628 33390
rect 32588 32972 32640 32978
rect 32588 32914 32640 32920
rect 32692 32586 32720 34734
rect 32864 34682 32916 34688
rect 32772 34536 32824 34542
rect 32876 34524 32904 34682
rect 32824 34496 32904 34524
rect 32772 34478 32824 34484
rect 32950 34300 33258 34309
rect 32950 34298 32956 34300
rect 33012 34298 33036 34300
rect 33092 34298 33116 34300
rect 33172 34298 33196 34300
rect 33252 34298 33258 34300
rect 33012 34246 33014 34298
rect 33194 34246 33196 34298
rect 32950 34244 32956 34246
rect 33012 34244 33036 34246
rect 33092 34244 33116 34246
rect 33172 34244 33196 34246
rect 33252 34244 33258 34246
rect 32950 34235 33258 34244
rect 33336 34066 33364 37266
rect 33416 37188 33468 37194
rect 33416 37130 33468 37136
rect 33324 34060 33376 34066
rect 33324 34002 33376 34008
rect 33140 33924 33192 33930
rect 33140 33866 33192 33872
rect 33048 33856 33100 33862
rect 33048 33798 33100 33804
rect 33060 33318 33088 33798
rect 33152 33658 33180 33866
rect 33232 33856 33284 33862
rect 33232 33798 33284 33804
rect 33140 33652 33192 33658
rect 33140 33594 33192 33600
rect 33244 33402 33272 33798
rect 33244 33374 33364 33402
rect 33048 33312 33100 33318
rect 33048 33254 33100 33260
rect 32950 33212 33258 33221
rect 32950 33210 32956 33212
rect 33012 33210 33036 33212
rect 33092 33210 33116 33212
rect 33172 33210 33196 33212
rect 33252 33210 33258 33212
rect 33012 33158 33014 33210
rect 33194 33158 33196 33210
rect 32950 33156 32956 33158
rect 33012 33156 33036 33158
rect 33092 33156 33116 33158
rect 33172 33156 33196 33158
rect 33252 33156 33258 33158
rect 32950 33147 33258 33156
rect 33336 32994 33364 33374
rect 33152 32966 33364 32994
rect 33152 32842 33180 32966
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 32692 32558 32904 32586
rect 32876 32434 32904 32558
rect 32680 32428 32732 32434
rect 32680 32370 32732 32376
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 32692 31346 32720 32370
rect 32772 32360 32824 32366
rect 32772 32302 32824 32308
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 32784 29238 32812 32302
rect 32950 32124 33258 32133
rect 32950 32122 32956 32124
rect 33012 32122 33036 32124
rect 33092 32122 33116 32124
rect 33172 32122 33196 32124
rect 33252 32122 33258 32124
rect 33012 32070 33014 32122
rect 33194 32070 33196 32122
rect 32950 32068 32956 32070
rect 33012 32068 33036 32070
rect 33092 32068 33116 32070
rect 33172 32068 33196 32070
rect 33252 32068 33258 32070
rect 32950 32059 33258 32068
rect 32950 31036 33258 31045
rect 32950 31034 32956 31036
rect 33012 31034 33036 31036
rect 33092 31034 33116 31036
rect 33172 31034 33196 31036
rect 33252 31034 33258 31036
rect 33012 30982 33014 31034
rect 33194 30982 33196 31034
rect 32950 30980 32956 30982
rect 33012 30980 33036 30982
rect 33092 30980 33116 30982
rect 33172 30980 33196 30982
rect 33252 30980 33258 30982
rect 32950 30971 33258 30980
rect 32950 29948 33258 29957
rect 32950 29946 32956 29948
rect 33012 29946 33036 29948
rect 33092 29946 33116 29948
rect 33172 29946 33196 29948
rect 33252 29946 33258 29948
rect 33012 29894 33014 29946
rect 33194 29894 33196 29946
rect 32950 29892 32956 29894
rect 33012 29892 33036 29894
rect 33092 29892 33116 29894
rect 33172 29892 33196 29894
rect 33252 29892 33258 29894
rect 32950 29883 33258 29892
rect 32772 29232 32824 29238
rect 32772 29174 32824 29180
rect 32950 28860 33258 28869
rect 32950 28858 32956 28860
rect 33012 28858 33036 28860
rect 33092 28858 33116 28860
rect 33172 28858 33196 28860
rect 33252 28858 33258 28860
rect 33012 28806 33014 28858
rect 33194 28806 33196 28858
rect 32950 28804 32956 28806
rect 33012 28804 33036 28806
rect 33092 28804 33116 28806
rect 33172 28804 33196 28806
rect 33252 28804 33258 28806
rect 32950 28795 33258 28804
rect 32950 27772 33258 27781
rect 32950 27770 32956 27772
rect 33012 27770 33036 27772
rect 33092 27770 33116 27772
rect 33172 27770 33196 27772
rect 33252 27770 33258 27772
rect 33012 27718 33014 27770
rect 33194 27718 33196 27770
rect 32950 27716 32956 27718
rect 33012 27716 33036 27718
rect 33092 27716 33116 27718
rect 33172 27716 33196 27718
rect 33252 27716 33258 27718
rect 32950 27707 33258 27716
rect 32950 26684 33258 26693
rect 32950 26682 32956 26684
rect 33012 26682 33036 26684
rect 33092 26682 33116 26684
rect 33172 26682 33196 26684
rect 33252 26682 33258 26684
rect 33012 26630 33014 26682
rect 33194 26630 33196 26682
rect 32950 26628 32956 26630
rect 33012 26628 33036 26630
rect 33092 26628 33116 26630
rect 33172 26628 33196 26630
rect 33252 26628 33258 26630
rect 32950 26619 33258 26628
rect 32950 25596 33258 25605
rect 32950 25594 32956 25596
rect 33012 25594 33036 25596
rect 33092 25594 33116 25596
rect 33172 25594 33196 25596
rect 33252 25594 33258 25596
rect 33012 25542 33014 25594
rect 33194 25542 33196 25594
rect 32950 25540 32956 25542
rect 33012 25540 33036 25542
rect 33092 25540 33116 25542
rect 33172 25540 33196 25542
rect 33252 25540 33258 25542
rect 32950 25531 33258 25540
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32508 22066 32720 22094
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 30760 7410 30788 8570
rect 31036 8498 31064 13262
rect 32692 8498 32720 22066
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33336 9994 33364 32370
rect 33428 32026 33456 37130
rect 33508 36916 33560 36922
rect 33508 36858 33560 36864
rect 33520 36378 33548 36858
rect 33508 36372 33560 36378
rect 33508 36314 33560 36320
rect 33520 34542 33548 36314
rect 33508 34536 33560 34542
rect 33508 34478 33560 34484
rect 33508 32972 33560 32978
rect 33508 32914 33560 32920
rect 33416 32020 33468 32026
rect 33416 31962 33468 31968
rect 33520 31754 33548 32914
rect 33612 32570 33640 38898
rect 33692 38888 33744 38894
rect 33692 38830 33744 38836
rect 33704 35630 33732 38830
rect 33796 37806 33824 42502
rect 33888 41682 33916 47058
rect 33980 44878 34008 48486
rect 34348 47122 34376 48622
rect 34520 48612 34572 48618
rect 34520 48554 34572 48560
rect 34532 48249 34560 48554
rect 34518 48240 34574 48249
rect 34518 48175 34574 48184
rect 34336 47116 34388 47122
rect 34336 47058 34388 47064
rect 34428 47116 34480 47122
rect 34428 47058 34480 47064
rect 34440 46374 34468 47058
rect 34532 46578 34560 48175
rect 34612 47456 34664 47462
rect 34612 47398 34664 47404
rect 34520 46572 34572 46578
rect 34520 46514 34572 46520
rect 34428 46368 34480 46374
rect 34428 46310 34480 46316
rect 34532 46034 34560 46514
rect 34520 46028 34572 46034
rect 34520 45970 34572 45976
rect 34152 45960 34204 45966
rect 34152 45902 34204 45908
rect 34164 45626 34192 45902
rect 34244 45892 34296 45898
rect 34244 45834 34296 45840
rect 34256 45626 34284 45834
rect 34152 45620 34204 45626
rect 34152 45562 34204 45568
rect 34244 45620 34296 45626
rect 34244 45562 34296 45568
rect 34336 45552 34388 45558
rect 34336 45494 34388 45500
rect 34060 45484 34112 45490
rect 34060 45426 34112 45432
rect 34072 44946 34100 45426
rect 34152 45348 34204 45354
rect 34152 45290 34204 45296
rect 34164 45082 34192 45290
rect 34152 45076 34204 45082
rect 34152 45018 34204 45024
rect 34060 44940 34112 44946
rect 34060 44882 34112 44888
rect 33968 44872 34020 44878
rect 33968 44814 34020 44820
rect 34348 44554 34376 45494
rect 34164 44526 34376 44554
rect 33968 43920 34020 43926
rect 33968 43862 34020 43868
rect 33980 43654 34008 43862
rect 33968 43648 34020 43654
rect 33968 43590 34020 43596
rect 33876 41676 33928 41682
rect 33876 41618 33928 41624
rect 33968 40384 34020 40390
rect 33968 40326 34020 40332
rect 33876 40112 33928 40118
rect 33874 40080 33876 40089
rect 33928 40080 33930 40089
rect 33874 40015 33930 40024
rect 33876 39976 33928 39982
rect 33876 39918 33928 39924
rect 33888 38894 33916 39918
rect 33980 39302 34008 40326
rect 34060 39840 34112 39846
rect 34060 39782 34112 39788
rect 34072 39642 34100 39782
rect 34060 39636 34112 39642
rect 34060 39578 34112 39584
rect 34060 39500 34112 39506
rect 34060 39442 34112 39448
rect 33968 39296 34020 39302
rect 33966 39264 33968 39273
rect 34020 39264 34022 39273
rect 33966 39199 34022 39208
rect 33968 38956 34020 38962
rect 33968 38898 34020 38904
rect 33876 38888 33928 38894
rect 33876 38830 33928 38836
rect 33876 38208 33928 38214
rect 33876 38150 33928 38156
rect 33784 37800 33836 37806
rect 33784 37742 33836 37748
rect 33888 35834 33916 38150
rect 33876 35828 33928 35834
rect 33876 35770 33928 35776
rect 33692 35624 33744 35630
rect 33692 35566 33744 35572
rect 33980 35562 34008 38898
rect 34072 35834 34100 39442
rect 34164 39370 34192 44526
rect 34336 44328 34388 44334
rect 34336 44270 34388 44276
rect 34428 44328 34480 44334
rect 34428 44270 34480 44276
rect 34348 43110 34376 44270
rect 34336 43104 34388 43110
rect 34336 43046 34388 43052
rect 34244 42356 34296 42362
rect 34244 42298 34296 42304
rect 34256 41206 34284 42298
rect 34336 41676 34388 41682
rect 34336 41618 34388 41624
rect 34244 41200 34296 41206
rect 34244 41142 34296 41148
rect 34348 40662 34376 41618
rect 34336 40656 34388 40662
rect 34336 40598 34388 40604
rect 34348 39574 34376 40598
rect 34440 40186 34468 44270
rect 34624 44198 34652 47398
rect 34716 47138 34744 49166
rect 35268 48890 35296 50390
rect 35348 49088 35400 49094
rect 35348 49030 35400 49036
rect 35256 48884 35308 48890
rect 35256 48826 35308 48832
rect 35360 48346 35388 49030
rect 34796 48340 34848 48346
rect 34796 48282 34848 48288
rect 35348 48340 35400 48346
rect 35348 48282 35400 48288
rect 34808 47802 34836 48282
rect 35348 48204 35400 48210
rect 35348 48146 35400 48152
rect 34980 48000 35032 48006
rect 34980 47942 35032 47948
rect 34796 47796 34848 47802
rect 34796 47738 34848 47744
rect 34888 47592 34940 47598
rect 34888 47534 34940 47540
rect 34900 47258 34928 47534
rect 34992 47462 35020 47942
rect 35256 47660 35308 47666
rect 35256 47602 35308 47608
rect 34980 47456 35032 47462
rect 34980 47398 35032 47404
rect 34888 47252 34940 47258
rect 34888 47194 34940 47200
rect 34716 47110 34836 47138
rect 34704 47048 34756 47054
rect 34704 46990 34756 46996
rect 34612 44192 34664 44198
rect 34612 44134 34664 44140
rect 34716 42378 34744 46990
rect 34808 46889 34836 47110
rect 34794 46880 34850 46889
rect 34794 46815 34850 46824
rect 34796 46504 34848 46510
rect 34796 46446 34848 46452
rect 34808 45422 34836 46446
rect 34888 46028 34940 46034
rect 34888 45970 34940 45976
rect 34796 45416 34848 45422
rect 34796 45358 34848 45364
rect 34808 45082 34836 45358
rect 34796 45076 34848 45082
rect 34796 45018 34848 45024
rect 34900 44946 34928 45970
rect 34888 44940 34940 44946
rect 34888 44882 34940 44888
rect 34900 43897 34928 44882
rect 34886 43888 34942 43897
rect 34886 43823 34888 43832
rect 34940 43823 34942 43832
rect 34888 43794 34940 43800
rect 34900 42770 34928 43794
rect 34888 42764 34940 42770
rect 34888 42706 34940 42712
rect 34624 42350 34744 42378
rect 34624 41414 34652 42350
rect 34900 41682 34928 42706
rect 34888 41676 34940 41682
rect 34888 41618 34940 41624
rect 34992 41414 35020 47398
rect 35268 47054 35296 47602
rect 35256 47048 35308 47054
rect 35256 46990 35308 46996
rect 35360 46510 35388 48146
rect 35452 48006 35480 51046
rect 36358 48104 36414 48113
rect 36358 48039 36360 48048
rect 36412 48039 36414 48048
rect 36360 48010 36412 48016
rect 35440 48000 35492 48006
rect 35440 47942 35492 47948
rect 35716 48000 35768 48006
rect 35716 47942 35768 47948
rect 36268 48000 36320 48006
rect 36268 47942 36320 47948
rect 35348 46504 35400 46510
rect 35348 46446 35400 46452
rect 35360 45898 35388 46446
rect 35452 46170 35480 47942
rect 35728 47462 35756 47942
rect 35808 47592 35860 47598
rect 35808 47534 35860 47540
rect 35716 47456 35768 47462
rect 35716 47398 35768 47404
rect 35820 47122 35848 47534
rect 35808 47116 35860 47122
rect 35808 47058 35860 47064
rect 36084 46980 36136 46986
rect 36084 46922 36136 46928
rect 35440 46164 35492 46170
rect 35440 46106 35492 46112
rect 35440 46028 35492 46034
rect 35440 45970 35492 45976
rect 35348 45892 35400 45898
rect 35348 45834 35400 45840
rect 35256 45280 35308 45286
rect 35256 45222 35308 45228
rect 35164 44804 35216 44810
rect 35164 44746 35216 44752
rect 35176 44169 35204 44746
rect 35162 44160 35218 44169
rect 35162 44095 35218 44104
rect 35164 43376 35216 43382
rect 35164 43318 35216 43324
rect 35176 42294 35204 43318
rect 35164 42288 35216 42294
rect 35164 42230 35216 42236
rect 35176 42106 35204 42230
rect 35268 42226 35296 45222
rect 35348 44396 35400 44402
rect 35348 44338 35400 44344
rect 35360 43314 35388 44338
rect 35348 43308 35400 43314
rect 35348 43250 35400 43256
rect 35256 42220 35308 42226
rect 35256 42162 35308 42168
rect 35176 42078 35296 42106
rect 35164 42016 35216 42022
rect 34624 41386 34744 41414
rect 34520 41064 34572 41070
rect 34520 41006 34572 41012
rect 34532 40526 34560 41006
rect 34612 40928 34664 40934
rect 34612 40870 34664 40876
rect 34520 40520 34572 40526
rect 34520 40462 34572 40468
rect 34428 40180 34480 40186
rect 34428 40122 34480 40128
rect 34532 40050 34560 40462
rect 34520 40044 34572 40050
rect 34520 39986 34572 39992
rect 34428 39976 34480 39982
rect 34428 39918 34480 39924
rect 34336 39568 34388 39574
rect 34256 39528 34336 39556
rect 34152 39364 34204 39370
rect 34152 39306 34204 39312
rect 34256 38214 34284 39528
rect 34336 39510 34388 39516
rect 34440 38654 34468 39918
rect 34532 39438 34560 39986
rect 34520 39432 34572 39438
rect 34520 39374 34572 39380
rect 34624 39030 34652 40870
rect 34612 39024 34664 39030
rect 34612 38966 34664 38972
rect 34440 38626 34560 38654
rect 34244 38208 34296 38214
rect 34244 38150 34296 38156
rect 34428 37936 34480 37942
rect 34428 37878 34480 37884
rect 34244 37664 34296 37670
rect 34244 37606 34296 37612
rect 34256 37369 34284 37606
rect 34242 37360 34298 37369
rect 34242 37295 34298 37304
rect 34152 37256 34204 37262
rect 34152 37198 34204 37204
rect 34164 36718 34192 37198
rect 34440 36786 34468 37878
rect 34428 36780 34480 36786
rect 34428 36722 34480 36728
rect 34152 36712 34204 36718
rect 34152 36654 34204 36660
rect 34164 36106 34192 36654
rect 34152 36100 34204 36106
rect 34152 36042 34204 36048
rect 34060 35828 34112 35834
rect 34060 35770 34112 35776
rect 34164 35630 34192 36042
rect 34152 35624 34204 35630
rect 34152 35566 34204 35572
rect 33968 35556 34020 35562
rect 33968 35498 34020 35504
rect 33784 35488 33836 35494
rect 33784 35430 33836 35436
rect 33796 35086 33824 35430
rect 34164 35086 34192 35566
rect 34440 35494 34468 36722
rect 34428 35488 34480 35494
rect 34428 35430 34480 35436
rect 33784 35080 33836 35086
rect 33784 35022 33836 35028
rect 34152 35080 34204 35086
rect 34152 35022 34204 35028
rect 34428 35080 34480 35086
rect 34428 35022 34480 35028
rect 33692 35012 33744 35018
rect 33692 34954 33744 34960
rect 34244 35012 34296 35018
rect 34244 34954 34296 34960
rect 33704 34406 33732 34954
rect 34060 34672 34112 34678
rect 34060 34614 34112 34620
rect 33692 34400 33744 34406
rect 33692 34342 33744 34348
rect 33692 33652 33744 33658
rect 33692 33594 33744 33600
rect 33704 33454 33732 33594
rect 33784 33584 33836 33590
rect 33784 33526 33836 33532
rect 33692 33448 33744 33454
rect 33692 33390 33744 33396
rect 33600 32564 33652 32570
rect 33600 32506 33652 32512
rect 33704 31890 33732 33390
rect 33796 32960 33824 33526
rect 34072 33454 34100 34614
rect 34150 34096 34206 34105
rect 34150 34031 34206 34040
rect 34164 33998 34192 34031
rect 34152 33992 34204 33998
rect 34152 33934 34204 33940
rect 34060 33448 34112 33454
rect 34060 33390 34112 33396
rect 33796 32932 33916 32960
rect 33796 32434 33824 32932
rect 33888 32842 33916 32932
rect 33876 32836 33928 32842
rect 33876 32778 33928 32784
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33876 32428 33928 32434
rect 33876 32370 33928 32376
rect 33784 32020 33836 32026
rect 33784 31962 33836 31968
rect 33692 31884 33744 31890
rect 33692 31826 33744 31832
rect 33600 31816 33652 31822
rect 33600 31758 33652 31764
rect 33508 31748 33560 31754
rect 33508 31690 33560 31696
rect 33612 31414 33640 31758
rect 33600 31408 33652 31414
rect 33600 31350 33652 31356
rect 33612 30394 33640 31350
rect 33600 30388 33652 30394
rect 33600 30330 33652 30336
rect 33414 24848 33470 24857
rect 33414 24783 33470 24792
rect 33428 23798 33456 24783
rect 33796 24206 33824 31962
rect 33888 31142 33916 32370
rect 34256 32230 34284 34954
rect 34336 34604 34388 34610
rect 34336 34546 34388 34552
rect 34348 34202 34376 34546
rect 34440 34542 34468 35022
rect 34428 34536 34480 34542
rect 34428 34478 34480 34484
rect 34336 34196 34388 34202
rect 34336 34138 34388 34144
rect 34336 34060 34388 34066
rect 34336 34002 34388 34008
rect 34348 33386 34376 34002
rect 34336 33380 34388 33386
rect 34336 33322 34388 33328
rect 34244 32224 34296 32230
rect 34244 32166 34296 32172
rect 34532 31929 34560 38626
rect 34716 37670 34744 41386
rect 34900 41386 35020 41414
rect 35084 41976 35164 42004
rect 34900 39506 34928 41386
rect 35084 41290 35112 41976
rect 35164 41958 35216 41964
rect 35164 41676 35216 41682
rect 35164 41618 35216 41624
rect 34992 41262 35112 41290
rect 34888 39500 34940 39506
rect 34888 39442 34940 39448
rect 34888 38276 34940 38282
rect 34888 38218 34940 38224
rect 34704 37664 34756 37670
rect 34704 37606 34756 37612
rect 34716 36582 34744 37606
rect 34704 36576 34756 36582
rect 34704 36518 34756 36524
rect 34900 36174 34928 38218
rect 34888 36168 34940 36174
rect 34888 36110 34940 36116
rect 34704 35760 34756 35766
rect 34704 35702 34756 35708
rect 34716 34134 34744 35702
rect 34796 35216 34848 35222
rect 34796 35158 34848 35164
rect 34612 34128 34664 34134
rect 34612 34070 34664 34076
rect 34704 34128 34756 34134
rect 34704 34070 34756 34076
rect 34624 32230 34652 34070
rect 34612 32224 34664 32230
rect 34612 32166 34664 32172
rect 34518 31920 34574 31929
rect 34518 31855 34574 31864
rect 33876 31136 33928 31142
rect 33876 31078 33928 31084
rect 34808 28558 34836 35158
rect 34992 34950 35020 41262
rect 35072 40996 35124 41002
rect 35072 40938 35124 40944
rect 35084 40730 35112 40938
rect 35072 40724 35124 40730
rect 35072 40666 35124 40672
rect 35176 40526 35204 41618
rect 35268 41546 35296 42078
rect 35256 41540 35308 41546
rect 35256 41482 35308 41488
rect 35268 41206 35296 41482
rect 35256 41200 35308 41206
rect 35256 41142 35308 41148
rect 35164 40520 35216 40526
rect 35164 40462 35216 40468
rect 35268 40118 35296 41142
rect 35452 41138 35480 45970
rect 35532 45824 35584 45830
rect 35532 45766 35584 45772
rect 35544 43450 35572 45766
rect 35900 44940 35952 44946
rect 35900 44882 35952 44888
rect 35808 44736 35860 44742
rect 35808 44678 35860 44684
rect 35820 44418 35848 44678
rect 35636 44390 35848 44418
rect 35636 44198 35664 44390
rect 35716 44328 35768 44334
rect 35912 44282 35940 44882
rect 35716 44270 35768 44276
rect 35624 44192 35676 44198
rect 35624 44134 35676 44140
rect 35728 43858 35756 44270
rect 35820 44254 35940 44282
rect 35820 44198 35848 44254
rect 35808 44192 35860 44198
rect 35808 44134 35860 44140
rect 35716 43852 35768 43858
rect 35716 43794 35768 43800
rect 35532 43444 35584 43450
rect 35532 43386 35584 43392
rect 36096 42158 36124 46922
rect 36176 45280 36228 45286
rect 36176 45222 36228 45228
rect 36188 44266 36216 45222
rect 36176 44260 36228 44266
rect 36176 44202 36228 44208
rect 36280 43450 36308 47942
rect 36464 46986 36492 51046
rect 37108 51046 37228 51074
rect 37004 49904 37056 49910
rect 37004 49846 37056 49852
rect 36636 49768 36688 49774
rect 36636 49710 36688 49716
rect 36544 49360 36596 49366
rect 36544 49302 36596 49308
rect 36556 47122 36584 49302
rect 36648 47122 36676 49710
rect 36820 48204 36872 48210
rect 36820 48146 36872 48152
rect 36726 48104 36782 48113
rect 36726 48039 36728 48048
rect 36780 48039 36782 48048
rect 36728 48010 36780 48016
rect 36544 47116 36596 47122
rect 36544 47058 36596 47064
rect 36636 47116 36688 47122
rect 36636 47058 36688 47064
rect 36452 46980 36504 46986
rect 36452 46922 36504 46928
rect 36464 45422 36492 46922
rect 36544 46640 36596 46646
rect 36544 46582 36596 46588
rect 36556 45966 36584 46582
rect 36544 45960 36596 45966
rect 36544 45902 36596 45908
rect 36452 45416 36504 45422
rect 36452 45358 36504 45364
rect 36464 44985 36492 45358
rect 36450 44976 36506 44985
rect 36450 44911 36506 44920
rect 36556 44810 36584 45902
rect 36544 44804 36596 44810
rect 36544 44746 36596 44752
rect 36556 43858 36584 44746
rect 36544 43852 36596 43858
rect 36544 43794 36596 43800
rect 36360 43648 36412 43654
rect 36360 43590 36412 43596
rect 36268 43444 36320 43450
rect 36268 43386 36320 43392
rect 36176 43240 36228 43246
rect 36176 43182 36228 43188
rect 36084 42152 36136 42158
rect 36084 42094 36136 42100
rect 36084 41472 36136 41478
rect 36084 41414 36136 41420
rect 36096 41206 36124 41414
rect 36084 41200 36136 41206
rect 36084 41142 36136 41148
rect 35440 41132 35492 41138
rect 35360 41092 35440 41120
rect 35256 40112 35308 40118
rect 35256 40054 35308 40060
rect 35360 39982 35388 41092
rect 35440 41074 35492 41080
rect 35992 41064 36044 41070
rect 35992 41006 36044 41012
rect 35440 40180 35492 40186
rect 35440 40122 35492 40128
rect 35348 39976 35400 39982
rect 35348 39918 35400 39924
rect 35348 39500 35400 39506
rect 35348 39442 35400 39448
rect 35164 39364 35216 39370
rect 35164 39306 35216 39312
rect 35256 39364 35308 39370
rect 35256 39306 35308 39312
rect 35176 38962 35204 39306
rect 35268 39098 35296 39306
rect 35256 39092 35308 39098
rect 35256 39034 35308 39040
rect 35164 38956 35216 38962
rect 35164 38898 35216 38904
rect 35072 38820 35124 38826
rect 35072 38762 35124 38768
rect 35084 36582 35112 38762
rect 35176 38282 35204 38898
rect 35164 38276 35216 38282
rect 35164 38218 35216 38224
rect 35176 38010 35204 38218
rect 35164 38004 35216 38010
rect 35164 37946 35216 37952
rect 35360 36922 35388 39442
rect 35452 38894 35480 40122
rect 35440 38888 35492 38894
rect 35440 38830 35492 38836
rect 35452 38418 35480 38830
rect 35440 38412 35492 38418
rect 35440 38354 35492 38360
rect 35440 37800 35492 37806
rect 35440 37742 35492 37748
rect 35716 37800 35768 37806
rect 35716 37742 35768 37748
rect 35808 37800 35860 37806
rect 35808 37742 35860 37748
rect 35348 36916 35400 36922
rect 35348 36858 35400 36864
rect 35072 36576 35124 36582
rect 35072 36518 35124 36524
rect 35360 36106 35388 36858
rect 35348 36100 35400 36106
rect 35348 36042 35400 36048
rect 35164 35624 35216 35630
rect 35164 35566 35216 35572
rect 35176 35154 35204 35566
rect 35164 35148 35216 35154
rect 35164 35090 35216 35096
rect 34980 34944 35032 34950
rect 34980 34886 35032 34892
rect 35452 32570 35480 37742
rect 35728 37670 35756 37742
rect 35716 37664 35768 37670
rect 35716 37606 35768 37612
rect 35820 37210 35848 37742
rect 36004 37369 36032 41006
rect 36096 40458 36124 41142
rect 36084 40452 36136 40458
rect 36084 40394 36136 40400
rect 36096 40066 36124 40394
rect 36188 40186 36216 43182
rect 36266 42392 36322 42401
rect 36266 42327 36322 42336
rect 36280 42294 36308 42327
rect 36268 42288 36320 42294
rect 36268 42230 36320 42236
rect 36372 41414 36400 43590
rect 36556 42702 36584 43794
rect 36544 42696 36596 42702
rect 36464 42656 36544 42684
rect 36464 41546 36492 42656
rect 36544 42638 36596 42644
rect 36648 42242 36676 47058
rect 36832 46034 36860 48146
rect 36820 46028 36872 46034
rect 36820 45970 36872 45976
rect 36912 44940 36964 44946
rect 36912 44882 36964 44888
rect 36820 44328 36872 44334
rect 36820 44270 36872 44276
rect 36832 43654 36860 44270
rect 36820 43648 36872 43654
rect 36820 43590 36872 43596
rect 36832 42906 36860 43590
rect 36820 42900 36872 42906
rect 36820 42842 36872 42848
rect 36556 42214 36676 42242
rect 36556 41818 36584 42214
rect 36636 42152 36688 42158
rect 36636 42094 36688 42100
rect 36544 41812 36596 41818
rect 36544 41754 36596 41760
rect 36452 41540 36504 41546
rect 36452 41482 36504 41488
rect 36372 41386 36584 41414
rect 36556 41274 36584 41386
rect 36544 41268 36596 41274
rect 36544 41210 36596 41216
rect 36176 40180 36228 40186
rect 36176 40122 36228 40128
rect 36096 40038 36308 40066
rect 36280 39370 36308 40038
rect 36268 39364 36320 39370
rect 36188 39324 36268 39352
rect 36084 39296 36136 39302
rect 36084 39238 36136 39244
rect 35990 37360 36046 37369
rect 35990 37295 36046 37304
rect 35636 37182 35848 37210
rect 35636 35170 35664 37182
rect 35808 37120 35860 37126
rect 35808 37062 35860 37068
rect 35544 35142 35664 35170
rect 35544 33862 35572 35142
rect 35820 34542 35848 37062
rect 35992 35828 36044 35834
rect 35992 35770 36044 35776
rect 35808 34536 35860 34542
rect 35808 34478 35860 34484
rect 36004 34406 36032 35770
rect 35992 34400 36044 34406
rect 35992 34342 36044 34348
rect 36096 33998 36124 39238
rect 36188 39030 36216 39324
rect 36268 39306 36320 39312
rect 36176 39024 36228 39030
rect 36176 38966 36228 38972
rect 36188 38654 36216 38966
rect 36188 38626 36400 38654
rect 36176 38276 36228 38282
rect 36176 38218 36228 38224
rect 36084 33992 36136 33998
rect 36084 33934 36136 33940
rect 35532 33856 35584 33862
rect 35532 33798 35584 33804
rect 36188 33318 36216 38218
rect 36372 37194 36400 38626
rect 36648 38350 36676 42094
rect 36924 41818 36952 44882
rect 37016 44810 37044 49846
rect 37108 49842 37136 51046
rect 37096 49836 37148 49842
rect 37096 49778 37148 49784
rect 37108 48113 37136 49778
rect 37188 49156 37240 49162
rect 37188 49098 37240 49104
rect 37094 48104 37150 48113
rect 37094 48039 37150 48048
rect 37200 47258 37228 49098
rect 37292 48249 37320 51342
rect 37384 51074 37412 53450
rect 37384 51046 37504 51074
rect 37372 48272 37424 48278
rect 37278 48240 37334 48249
rect 37372 48214 37424 48220
rect 37278 48175 37334 48184
rect 37188 47252 37240 47258
rect 37188 47194 37240 47200
rect 37096 47184 37148 47190
rect 37096 47126 37148 47132
rect 37108 44878 37136 47126
rect 37188 45824 37240 45830
rect 37188 45766 37240 45772
rect 37096 44872 37148 44878
rect 37096 44814 37148 44820
rect 37004 44804 37056 44810
rect 37004 44746 37056 44752
rect 37200 44334 37228 45766
rect 37384 45286 37412 48214
rect 37476 47462 37504 51046
rect 37568 47666 37596 53926
rect 38660 53712 38712 53718
rect 38660 53654 38712 53660
rect 38292 53644 38344 53650
rect 38292 53586 38344 53592
rect 37950 53340 38258 53349
rect 37950 53338 37956 53340
rect 38012 53338 38036 53340
rect 38092 53338 38116 53340
rect 38172 53338 38196 53340
rect 38252 53338 38258 53340
rect 38012 53286 38014 53338
rect 38194 53286 38196 53338
rect 37950 53284 37956 53286
rect 38012 53284 38036 53286
rect 38092 53284 38116 53286
rect 38172 53284 38196 53286
rect 38252 53284 38258 53286
rect 37950 53275 38258 53284
rect 37950 52252 38258 52261
rect 37950 52250 37956 52252
rect 38012 52250 38036 52252
rect 38092 52250 38116 52252
rect 38172 52250 38196 52252
rect 38252 52250 38258 52252
rect 38012 52198 38014 52250
rect 38194 52198 38196 52250
rect 37950 52196 37956 52198
rect 38012 52196 38036 52198
rect 38092 52196 38116 52198
rect 38172 52196 38196 52198
rect 38252 52196 38258 52198
rect 37950 52187 38258 52196
rect 37950 51164 38258 51173
rect 37950 51162 37956 51164
rect 38012 51162 38036 51164
rect 38092 51162 38116 51164
rect 38172 51162 38196 51164
rect 38252 51162 38258 51164
rect 38012 51110 38014 51162
rect 38194 51110 38196 51162
rect 37950 51108 37956 51110
rect 38012 51108 38036 51110
rect 38092 51108 38116 51110
rect 38172 51108 38196 51110
rect 38252 51108 38258 51110
rect 37950 51099 38258 51108
rect 37950 50076 38258 50085
rect 37950 50074 37956 50076
rect 38012 50074 38036 50076
rect 38092 50074 38116 50076
rect 38172 50074 38196 50076
rect 38252 50074 38258 50076
rect 38012 50022 38014 50074
rect 38194 50022 38196 50074
rect 37950 50020 37956 50022
rect 38012 50020 38036 50022
rect 38092 50020 38116 50022
rect 38172 50020 38196 50022
rect 38252 50020 38258 50022
rect 37950 50011 38258 50020
rect 37950 48988 38258 48997
rect 37950 48986 37956 48988
rect 38012 48986 38036 48988
rect 38092 48986 38116 48988
rect 38172 48986 38196 48988
rect 38252 48986 38258 48988
rect 38012 48934 38014 48986
rect 38194 48934 38196 48986
rect 37950 48932 37956 48934
rect 38012 48932 38036 48934
rect 38092 48932 38116 48934
rect 38172 48932 38196 48934
rect 38252 48932 38258 48934
rect 37950 48923 38258 48932
rect 37950 47900 38258 47909
rect 37950 47898 37956 47900
rect 38012 47898 38036 47900
rect 38092 47898 38116 47900
rect 38172 47898 38196 47900
rect 38252 47898 38258 47900
rect 38012 47846 38014 47898
rect 38194 47846 38196 47898
rect 37950 47844 37956 47846
rect 38012 47844 38036 47846
rect 38092 47844 38116 47846
rect 38172 47844 38196 47846
rect 38252 47844 38258 47846
rect 37950 47835 38258 47844
rect 37556 47660 37608 47666
rect 37556 47602 37608 47608
rect 37464 47456 37516 47462
rect 37464 47398 37516 47404
rect 37464 45416 37516 45422
rect 37464 45358 37516 45364
rect 37372 45280 37424 45286
rect 37372 45222 37424 45228
rect 37372 45008 37424 45014
rect 37372 44950 37424 44956
rect 37188 44328 37240 44334
rect 37188 44270 37240 44276
rect 37278 43888 37334 43897
rect 37278 43823 37280 43832
rect 37332 43823 37334 43832
rect 37280 43794 37332 43800
rect 37004 43104 37056 43110
rect 37004 43046 37056 43052
rect 36728 41812 36780 41818
rect 36728 41754 36780 41760
rect 36912 41812 36964 41818
rect 36912 41754 36964 41760
rect 36740 41070 36768 41754
rect 36912 41676 36964 41682
rect 36912 41618 36964 41624
rect 36728 41064 36780 41070
rect 36728 41006 36780 41012
rect 36924 39302 36952 41618
rect 36912 39296 36964 39302
rect 36912 39238 36964 39244
rect 36924 38894 36952 39238
rect 36912 38888 36964 38894
rect 36912 38830 36964 38836
rect 36820 38412 36872 38418
rect 36820 38354 36872 38360
rect 36636 38344 36688 38350
rect 36636 38286 36688 38292
rect 36452 38208 36504 38214
rect 36452 38150 36504 38156
rect 36636 38208 36688 38214
rect 36636 38150 36688 38156
rect 36728 38208 36780 38214
rect 36728 38150 36780 38156
rect 36464 37942 36492 38150
rect 36452 37936 36504 37942
rect 36452 37878 36504 37884
rect 36542 37904 36598 37913
rect 36542 37839 36598 37848
rect 36360 37188 36412 37194
rect 36360 37130 36412 37136
rect 36372 36786 36400 37130
rect 36556 36854 36584 37839
rect 36544 36848 36596 36854
rect 36544 36790 36596 36796
rect 36360 36780 36412 36786
rect 36360 36722 36412 36728
rect 36372 36174 36400 36722
rect 36360 36168 36412 36174
rect 36360 36110 36412 36116
rect 36372 35630 36400 36110
rect 36360 35624 36412 35630
rect 36360 35566 36412 35572
rect 36268 35080 36320 35086
rect 36372 35068 36400 35566
rect 36320 35040 36400 35068
rect 36268 35022 36320 35028
rect 36280 34678 36308 35022
rect 36648 34746 36676 38150
rect 36740 38010 36768 38150
rect 36728 38004 36780 38010
rect 36728 37946 36780 37952
rect 36832 37330 36860 38354
rect 37016 37874 37044 43046
rect 37292 41138 37320 43794
rect 37188 41132 37240 41138
rect 37188 41074 37240 41080
rect 37280 41132 37332 41138
rect 37280 41074 37332 41080
rect 37200 40730 37228 41074
rect 37096 40724 37148 40730
rect 37096 40666 37148 40672
rect 37188 40724 37240 40730
rect 37188 40666 37240 40672
rect 37108 40594 37136 40666
rect 37096 40588 37148 40594
rect 37096 40530 37148 40536
rect 37384 39642 37412 44950
rect 37476 44266 37504 45358
rect 37568 44826 37596 47602
rect 37832 47456 37884 47462
rect 37832 47398 37884 47404
rect 37844 45966 37872 47398
rect 38304 47054 38332 53586
rect 38292 47048 38344 47054
rect 38292 46990 38344 46996
rect 37950 46812 38258 46821
rect 37950 46810 37956 46812
rect 38012 46810 38036 46812
rect 38092 46810 38116 46812
rect 38172 46810 38196 46812
rect 38252 46810 38258 46812
rect 38012 46758 38014 46810
rect 38194 46758 38196 46810
rect 37950 46756 37956 46758
rect 38012 46756 38036 46758
rect 38092 46756 38116 46758
rect 38172 46756 38196 46758
rect 38252 46756 38258 46758
rect 37950 46747 38258 46756
rect 37832 45960 37884 45966
rect 37832 45902 37884 45908
rect 37740 45824 37792 45830
rect 37740 45766 37792 45772
rect 37752 44946 37780 45766
rect 37950 45724 38258 45733
rect 37950 45722 37956 45724
rect 38012 45722 38036 45724
rect 38092 45722 38116 45724
rect 38172 45722 38196 45724
rect 38252 45722 38258 45724
rect 38012 45670 38014 45722
rect 38194 45670 38196 45722
rect 37950 45668 37956 45670
rect 38012 45668 38036 45670
rect 38092 45668 38116 45670
rect 38172 45668 38196 45670
rect 38252 45668 38258 45670
rect 37950 45659 38258 45668
rect 38016 45416 38068 45422
rect 38016 45358 38068 45364
rect 38028 45082 38056 45358
rect 38016 45076 38068 45082
rect 38016 45018 38068 45024
rect 37740 44940 37792 44946
rect 37740 44882 37792 44888
rect 37568 44798 37780 44826
rect 37556 44736 37608 44742
rect 37556 44678 37608 44684
rect 37568 44538 37596 44678
rect 37556 44532 37608 44538
rect 37556 44474 37608 44480
rect 37648 44532 37700 44538
rect 37648 44474 37700 44480
rect 37464 44260 37516 44266
rect 37464 44202 37516 44208
rect 37556 44260 37608 44266
rect 37556 44202 37608 44208
rect 37568 43722 37596 44202
rect 37556 43716 37608 43722
rect 37556 43658 37608 43664
rect 37568 43353 37596 43658
rect 37554 43344 37610 43353
rect 37554 43279 37610 43288
rect 37660 41414 37688 44474
rect 37752 44402 37780 44798
rect 37950 44636 38258 44645
rect 37950 44634 37956 44636
rect 38012 44634 38036 44636
rect 38092 44634 38116 44636
rect 38172 44634 38196 44636
rect 38252 44634 38258 44636
rect 38012 44582 38014 44634
rect 38194 44582 38196 44634
rect 37950 44580 37956 44582
rect 38012 44580 38036 44582
rect 38092 44580 38116 44582
rect 38172 44580 38196 44582
rect 38252 44580 38258 44582
rect 37950 44571 38258 44580
rect 38304 44538 38332 46990
rect 38672 45626 38700 53654
rect 38948 53582 38976 56200
rect 39120 54256 39172 54262
rect 39120 54198 39172 54204
rect 38936 53576 38988 53582
rect 38936 53518 38988 53524
rect 39028 53440 39080 53446
rect 39028 53382 39080 53388
rect 38936 51808 38988 51814
rect 38936 51750 38988 51756
rect 38948 47598 38976 51750
rect 39040 49978 39068 53382
rect 39028 49972 39080 49978
rect 39028 49914 39080 49920
rect 39028 48000 39080 48006
rect 39028 47942 39080 47948
rect 38936 47592 38988 47598
rect 38936 47534 38988 47540
rect 39040 47122 39068 47942
rect 39028 47116 39080 47122
rect 39028 47058 39080 47064
rect 39132 45830 39160 54198
rect 39592 54194 39620 56200
rect 40236 55214 40264 56200
rect 40236 55186 40356 55214
rect 40328 54194 40356 55186
rect 40684 54528 40736 54534
rect 40684 54470 40736 54476
rect 39580 54188 39632 54194
rect 39580 54130 39632 54136
rect 40316 54188 40368 54194
rect 40316 54130 40368 54136
rect 40696 54058 40724 54470
rect 42168 54262 42196 56200
rect 40776 54256 40828 54262
rect 40776 54198 40828 54204
rect 42156 54256 42208 54262
rect 42156 54198 42208 54204
rect 40788 54058 40816 54198
rect 40684 54052 40736 54058
rect 40684 53994 40736 54000
rect 40776 54052 40828 54058
rect 40776 53994 40828 54000
rect 43904 53984 43956 53990
rect 43904 53926 43956 53932
rect 42950 53884 43258 53893
rect 42950 53882 42956 53884
rect 43012 53882 43036 53884
rect 43092 53882 43116 53884
rect 43172 53882 43196 53884
rect 43252 53882 43258 53884
rect 43012 53830 43014 53882
rect 43194 53830 43196 53882
rect 42950 53828 42956 53830
rect 43012 53828 43036 53830
rect 43092 53828 43116 53830
rect 43172 53828 43196 53830
rect 43252 53828 43258 53830
rect 42950 53819 43258 53828
rect 42950 52796 43258 52805
rect 42950 52794 42956 52796
rect 43012 52794 43036 52796
rect 43092 52794 43116 52796
rect 43172 52794 43196 52796
rect 43252 52794 43258 52796
rect 43012 52742 43014 52794
rect 43194 52742 43196 52794
rect 42950 52740 42956 52742
rect 43012 52740 43036 52742
rect 43092 52740 43116 52742
rect 43172 52740 43196 52742
rect 43252 52740 43258 52742
rect 42950 52731 43258 52740
rect 43444 51808 43496 51814
rect 43444 51750 43496 51756
rect 42950 51708 43258 51717
rect 42950 51706 42956 51708
rect 43012 51706 43036 51708
rect 43092 51706 43116 51708
rect 43172 51706 43196 51708
rect 43252 51706 43258 51708
rect 43012 51654 43014 51706
rect 43194 51654 43196 51706
rect 42950 51652 42956 51654
rect 43012 51652 43036 51654
rect 43092 51652 43116 51654
rect 43172 51652 43196 51654
rect 43252 51652 43258 51654
rect 42950 51643 43258 51652
rect 42156 51604 42208 51610
rect 42156 51546 42208 51552
rect 42168 51338 42196 51546
rect 43456 51406 43484 51750
rect 43916 51610 43944 53926
rect 44100 53582 44128 56200
rect 44744 54194 44772 56200
rect 45388 54618 45416 56200
rect 46032 55214 46060 56200
rect 46032 55186 46152 55214
rect 45388 54590 45692 54618
rect 45664 54262 45692 54590
rect 45836 54596 45888 54602
rect 45836 54538 45888 54544
rect 45848 54330 45876 54538
rect 45836 54324 45888 54330
rect 45836 54266 45888 54272
rect 45652 54256 45704 54262
rect 45652 54198 45704 54204
rect 46124 54194 46152 55186
rect 44732 54188 44784 54194
rect 44732 54130 44784 54136
rect 46112 54188 46164 54194
rect 46112 54130 46164 54136
rect 46676 53582 46704 56200
rect 47320 54194 47348 56200
rect 47964 55214 47992 56200
rect 47872 55186 47992 55214
rect 47766 54632 47822 54641
rect 47766 54567 47822 54576
rect 47308 54188 47360 54194
rect 47308 54130 47360 54136
rect 44088 53576 44140 53582
rect 44088 53518 44140 53524
rect 46664 53576 46716 53582
rect 46664 53518 46716 53524
rect 47780 53174 47808 54567
rect 47872 54194 47900 55186
rect 47950 54428 48258 54437
rect 47950 54426 47956 54428
rect 48012 54426 48036 54428
rect 48092 54426 48116 54428
rect 48172 54426 48196 54428
rect 48252 54426 48258 54428
rect 48012 54374 48014 54426
rect 48194 54374 48196 54426
rect 47950 54372 47956 54374
rect 48012 54372 48036 54374
rect 48092 54372 48116 54374
rect 48172 54372 48196 54374
rect 48252 54372 48258 54374
rect 47950 54363 48258 54372
rect 47860 54188 47912 54194
rect 47860 54130 47912 54136
rect 48318 53816 48374 53825
rect 48318 53751 48374 53760
rect 48332 53582 48360 53751
rect 48608 53582 48636 56200
rect 48688 53984 48740 53990
rect 48688 53926 48740 53932
rect 48320 53576 48372 53582
rect 48320 53518 48372 53524
rect 48596 53576 48648 53582
rect 48596 53518 48648 53524
rect 47950 53340 48258 53349
rect 47950 53338 47956 53340
rect 48012 53338 48036 53340
rect 48092 53338 48116 53340
rect 48172 53338 48196 53340
rect 48252 53338 48258 53340
rect 48012 53286 48014 53338
rect 48194 53286 48196 53338
rect 47950 53284 47956 53286
rect 48012 53284 48036 53286
rect 48092 53284 48116 53286
rect 48172 53284 48196 53286
rect 48252 53284 48258 53286
rect 47950 53275 48258 53284
rect 47768 53168 47820 53174
rect 47768 53110 47820 53116
rect 48504 53032 48556 53038
rect 48502 53000 48504 53009
rect 48556 53000 48558 53009
rect 48502 52935 48558 52944
rect 46204 52896 46256 52902
rect 46204 52838 46256 52844
rect 43904 51604 43956 51610
rect 43904 51546 43956 51552
rect 43444 51400 43496 51406
rect 43444 51342 43496 51348
rect 39304 51332 39356 51338
rect 39304 51274 39356 51280
rect 42156 51332 42208 51338
rect 42156 51274 42208 51280
rect 39316 46646 39344 51274
rect 42800 50720 42852 50726
rect 42800 50662 42852 50668
rect 42812 47802 42840 50662
rect 42950 50620 43258 50629
rect 42950 50618 42956 50620
rect 43012 50618 43036 50620
rect 43092 50618 43116 50620
rect 43172 50618 43196 50620
rect 43252 50618 43258 50620
rect 43012 50566 43014 50618
rect 43194 50566 43196 50618
rect 42950 50564 42956 50566
rect 43012 50564 43036 50566
rect 43092 50564 43116 50566
rect 43172 50564 43196 50566
rect 43252 50564 43258 50566
rect 42950 50555 43258 50564
rect 43444 49768 43496 49774
rect 43444 49710 43496 49716
rect 42950 49532 43258 49541
rect 42950 49530 42956 49532
rect 43012 49530 43036 49532
rect 43092 49530 43116 49532
rect 43172 49530 43196 49532
rect 43252 49530 43258 49532
rect 43012 49478 43014 49530
rect 43194 49478 43196 49530
rect 42950 49476 42956 49478
rect 43012 49476 43036 49478
rect 43092 49476 43116 49478
rect 43172 49476 43196 49478
rect 43252 49476 43258 49478
rect 42950 49467 43258 49476
rect 42950 48444 43258 48453
rect 42950 48442 42956 48444
rect 43012 48442 43036 48444
rect 43092 48442 43116 48444
rect 43172 48442 43196 48444
rect 43252 48442 43258 48444
rect 43012 48390 43014 48442
rect 43194 48390 43196 48442
rect 42950 48388 42956 48390
rect 43012 48388 43036 48390
rect 43092 48388 43116 48390
rect 43172 48388 43196 48390
rect 43252 48388 43258 48390
rect 42950 48379 43258 48388
rect 43352 48000 43404 48006
rect 43352 47942 43404 47948
rect 42800 47796 42852 47802
rect 42800 47738 42852 47744
rect 40132 47728 40184 47734
rect 40132 47670 40184 47676
rect 39764 47660 39816 47666
rect 39764 47602 39816 47608
rect 39304 46640 39356 46646
rect 39304 46582 39356 46588
rect 39120 45824 39172 45830
rect 39120 45766 39172 45772
rect 38660 45620 38712 45626
rect 38660 45562 38712 45568
rect 38672 45098 38700 45562
rect 38580 45070 38700 45098
rect 38384 44736 38436 44742
rect 38384 44678 38436 44684
rect 38292 44532 38344 44538
rect 38292 44474 38344 44480
rect 38396 44470 38424 44678
rect 38384 44464 38436 44470
rect 38384 44406 38436 44412
rect 37740 44396 37792 44402
rect 37740 44338 37792 44344
rect 38016 44328 38068 44334
rect 38016 44270 38068 44276
rect 38028 44169 38056 44270
rect 38014 44160 38070 44169
rect 38014 44095 38070 44104
rect 38580 43738 38608 45070
rect 38660 44940 38712 44946
rect 38660 44882 38712 44888
rect 38672 44198 38700 44882
rect 38752 44736 38804 44742
rect 38752 44678 38804 44684
rect 38660 44192 38712 44198
rect 38660 44134 38712 44140
rect 38672 43926 38700 44134
rect 38660 43920 38712 43926
rect 38660 43862 38712 43868
rect 38580 43710 38700 43738
rect 37950 43548 38258 43557
rect 37950 43546 37956 43548
rect 38012 43546 38036 43548
rect 38092 43546 38116 43548
rect 38172 43546 38196 43548
rect 38252 43546 38258 43548
rect 38012 43494 38014 43546
rect 38194 43494 38196 43546
rect 37950 43492 37956 43494
rect 38012 43492 38036 43494
rect 38092 43492 38116 43494
rect 38172 43492 38196 43494
rect 38252 43492 38258 43494
rect 37950 43483 38258 43492
rect 37832 42560 37884 42566
rect 37832 42502 37884 42508
rect 37568 41386 37688 41414
rect 37568 39846 37596 41386
rect 37740 41064 37792 41070
rect 37740 41006 37792 41012
rect 37646 40624 37702 40633
rect 37646 40559 37648 40568
rect 37700 40559 37702 40568
rect 37648 40530 37700 40536
rect 37660 40390 37688 40530
rect 37648 40384 37700 40390
rect 37648 40326 37700 40332
rect 37556 39840 37608 39846
rect 37556 39782 37608 39788
rect 37372 39636 37424 39642
rect 37372 39578 37424 39584
rect 37646 39536 37702 39545
rect 37646 39471 37702 39480
rect 37462 39400 37518 39409
rect 37462 39335 37464 39344
rect 37516 39335 37518 39344
rect 37464 39306 37516 39312
rect 37660 39030 37688 39471
rect 37648 39024 37700 39030
rect 37648 38966 37700 38972
rect 37004 37868 37056 37874
rect 37004 37810 37056 37816
rect 36820 37324 36872 37330
rect 36820 37266 36872 37272
rect 36912 37324 36964 37330
rect 36912 37266 36964 37272
rect 36832 36922 36860 37266
rect 36820 36916 36872 36922
rect 36820 36858 36872 36864
rect 36924 35834 36952 37266
rect 37660 37262 37688 38966
rect 37752 38418 37780 41006
rect 37844 40594 37872 42502
rect 37950 42460 38258 42469
rect 37950 42458 37956 42460
rect 38012 42458 38036 42460
rect 38092 42458 38116 42460
rect 38172 42458 38196 42460
rect 38252 42458 38258 42460
rect 38012 42406 38014 42458
rect 38194 42406 38196 42458
rect 37950 42404 37956 42406
rect 38012 42404 38036 42406
rect 38092 42404 38116 42406
rect 38172 42404 38196 42406
rect 38252 42404 38258 42406
rect 37950 42395 38258 42404
rect 37950 41372 38258 41381
rect 37950 41370 37956 41372
rect 38012 41370 38036 41372
rect 38092 41370 38116 41372
rect 38172 41370 38196 41372
rect 38252 41370 38258 41372
rect 38012 41318 38014 41370
rect 38194 41318 38196 41370
rect 37950 41316 37956 41318
rect 38012 41316 38036 41318
rect 38092 41316 38116 41318
rect 38172 41316 38196 41318
rect 38252 41316 38258 41318
rect 37950 41307 38258 41316
rect 37832 40588 37884 40594
rect 37832 40530 37884 40536
rect 37950 40284 38258 40293
rect 37950 40282 37956 40284
rect 38012 40282 38036 40284
rect 38092 40282 38116 40284
rect 38172 40282 38196 40284
rect 38252 40282 38258 40284
rect 38012 40230 38014 40282
rect 38194 40230 38196 40282
rect 37950 40228 37956 40230
rect 38012 40228 38036 40230
rect 38092 40228 38116 40230
rect 38172 40228 38196 40230
rect 38252 40228 38258 40230
rect 37950 40219 38258 40228
rect 38476 39840 38528 39846
rect 38476 39782 38528 39788
rect 38488 39302 38516 39782
rect 38476 39296 38528 39302
rect 38476 39238 38528 39244
rect 37950 39196 38258 39205
rect 37950 39194 37956 39196
rect 38012 39194 38036 39196
rect 38092 39194 38116 39196
rect 38172 39194 38196 39196
rect 38252 39194 38258 39196
rect 38012 39142 38014 39194
rect 38194 39142 38196 39194
rect 37950 39140 37956 39142
rect 38012 39140 38036 39142
rect 38092 39140 38116 39142
rect 38172 39140 38196 39142
rect 38252 39140 38258 39142
rect 37950 39131 38258 39140
rect 37832 39092 37884 39098
rect 37832 39034 37884 39040
rect 37740 38412 37792 38418
rect 37740 38354 37792 38360
rect 37844 37806 37872 39034
rect 38106 38992 38162 39001
rect 38106 38927 38108 38936
rect 38160 38927 38162 38936
rect 38108 38898 38160 38904
rect 38488 38321 38516 39238
rect 38672 39098 38700 43710
rect 38764 40934 38792 44678
rect 38844 43648 38896 43654
rect 38844 43590 38896 43596
rect 38856 41138 38884 43590
rect 38844 41132 38896 41138
rect 38844 41074 38896 41080
rect 38752 40928 38804 40934
rect 38752 40870 38804 40876
rect 38752 40180 38804 40186
rect 38752 40122 38804 40128
rect 38660 39092 38712 39098
rect 38660 39034 38712 39040
rect 38660 38752 38712 38758
rect 38660 38694 38712 38700
rect 38672 38350 38700 38694
rect 38660 38344 38712 38350
rect 38474 38312 38530 38321
rect 38660 38286 38712 38292
rect 38474 38247 38530 38256
rect 37950 38108 38258 38117
rect 37950 38106 37956 38108
rect 38012 38106 38036 38108
rect 38092 38106 38116 38108
rect 38172 38106 38196 38108
rect 38252 38106 38258 38108
rect 38012 38054 38014 38106
rect 38194 38054 38196 38106
rect 37950 38052 37956 38054
rect 38012 38052 38036 38054
rect 38092 38052 38116 38054
rect 38172 38052 38196 38054
rect 38252 38052 38258 38054
rect 37950 38043 38258 38052
rect 37832 37800 37884 37806
rect 37832 37742 37884 37748
rect 38568 37800 38620 37806
rect 38568 37742 38620 37748
rect 37648 37256 37700 37262
rect 37648 37198 37700 37204
rect 37556 37120 37608 37126
rect 37648 37120 37700 37126
rect 37556 37062 37608 37068
rect 37646 37088 37648 37097
rect 37700 37088 37702 37097
rect 37108 36230 37504 36258
rect 37108 36174 37136 36230
rect 37096 36168 37148 36174
rect 37096 36110 37148 36116
rect 37476 36106 37504 36230
rect 37372 36100 37424 36106
rect 37372 36042 37424 36048
rect 37464 36100 37516 36106
rect 37464 36042 37516 36048
rect 37096 36032 37148 36038
rect 37096 35974 37148 35980
rect 36912 35828 36964 35834
rect 36912 35770 36964 35776
rect 37108 34950 37136 35974
rect 37188 35284 37240 35290
rect 37188 35226 37240 35232
rect 37096 34944 37148 34950
rect 37096 34886 37148 34892
rect 36636 34740 36688 34746
rect 36636 34682 36688 34688
rect 36268 34672 36320 34678
rect 36268 34614 36320 34620
rect 36268 34400 36320 34406
rect 36268 34342 36320 34348
rect 36280 33658 36308 34342
rect 36268 33652 36320 33658
rect 36268 33594 36320 33600
rect 36176 33312 36228 33318
rect 36176 33254 36228 33260
rect 36728 32768 36780 32774
rect 36728 32710 36780 32716
rect 35440 32564 35492 32570
rect 35440 32506 35492 32512
rect 36544 32428 36596 32434
rect 36544 32370 36596 32376
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 36556 27946 36584 32370
rect 36740 32366 36768 32710
rect 36728 32360 36780 32366
rect 36728 32302 36780 32308
rect 37200 31346 37228 35226
rect 37188 31340 37240 31346
rect 37188 31282 37240 31288
rect 37384 30258 37412 36042
rect 37568 34746 37596 37062
rect 37646 37023 37702 37032
rect 37950 37020 38258 37029
rect 37950 37018 37956 37020
rect 38012 37018 38036 37020
rect 38092 37018 38116 37020
rect 38172 37018 38196 37020
rect 38252 37018 38258 37020
rect 38012 36966 38014 37018
rect 38194 36966 38196 37018
rect 37950 36964 37956 36966
rect 38012 36964 38036 36966
rect 38092 36964 38116 36966
rect 38172 36964 38196 36966
rect 38252 36964 38258 36966
rect 37950 36955 38258 36964
rect 38580 36378 38608 37742
rect 38660 37188 38712 37194
rect 38660 37130 38712 37136
rect 38568 36372 38620 36378
rect 38568 36314 38620 36320
rect 38672 36242 38700 37130
rect 38764 36922 38792 40122
rect 39132 40050 39160 45766
rect 39776 45558 39804 47602
rect 40144 46986 40172 47670
rect 42800 47456 42852 47462
rect 42800 47398 42852 47404
rect 40132 46980 40184 46986
rect 40132 46922 40184 46928
rect 39764 45552 39816 45558
rect 39764 45494 39816 45500
rect 39488 45416 39540 45422
rect 39488 45358 39540 45364
rect 39500 44334 39528 45358
rect 39672 44804 39724 44810
rect 39672 44746 39724 44752
rect 39684 44538 39712 44746
rect 39672 44532 39724 44538
rect 39672 44474 39724 44480
rect 39488 44328 39540 44334
rect 39488 44270 39540 44276
rect 39488 42016 39540 42022
rect 39488 41958 39540 41964
rect 39212 40928 39264 40934
rect 39212 40870 39264 40876
rect 39224 40458 39252 40870
rect 39212 40452 39264 40458
rect 39212 40394 39264 40400
rect 39120 40044 39172 40050
rect 39120 39986 39172 39992
rect 39224 39506 39252 40394
rect 39396 39976 39448 39982
rect 39396 39918 39448 39924
rect 39304 39636 39356 39642
rect 39304 39578 39356 39584
rect 38936 39500 38988 39506
rect 38936 39442 38988 39448
rect 39212 39500 39264 39506
rect 39212 39442 39264 39448
rect 38844 38820 38896 38826
rect 38844 38762 38896 38768
rect 38856 38282 38884 38762
rect 38948 38418 38976 39442
rect 39316 39370 39344 39578
rect 39120 39364 39172 39370
rect 39120 39306 39172 39312
rect 39304 39364 39356 39370
rect 39304 39306 39356 39312
rect 38936 38412 38988 38418
rect 38936 38354 38988 38360
rect 38844 38276 38896 38282
rect 38844 38218 38896 38224
rect 39132 38010 39160 39306
rect 39212 39296 39264 39302
rect 39212 39238 39264 39244
rect 39224 38554 39252 39238
rect 39304 38956 39356 38962
rect 39304 38898 39356 38904
rect 39212 38548 39264 38554
rect 39212 38490 39264 38496
rect 39120 38004 39172 38010
rect 39120 37946 39172 37952
rect 38752 36916 38804 36922
rect 38752 36858 38804 36864
rect 38844 36712 38896 36718
rect 38844 36654 38896 36660
rect 38660 36236 38712 36242
rect 38660 36178 38712 36184
rect 38856 36038 38884 36654
rect 38844 36032 38896 36038
rect 38844 35974 38896 35980
rect 37950 35932 38258 35941
rect 37950 35930 37956 35932
rect 38012 35930 38036 35932
rect 38092 35930 38116 35932
rect 38172 35930 38196 35932
rect 38252 35930 38258 35932
rect 38012 35878 38014 35930
rect 38194 35878 38196 35930
rect 37950 35876 37956 35878
rect 38012 35876 38036 35878
rect 38092 35876 38116 35878
rect 38172 35876 38196 35878
rect 38252 35876 38258 35878
rect 37950 35867 38258 35876
rect 37950 34844 38258 34853
rect 37950 34842 37956 34844
rect 38012 34842 38036 34844
rect 38092 34842 38116 34844
rect 38172 34842 38196 34844
rect 38252 34842 38258 34844
rect 38012 34790 38014 34842
rect 38194 34790 38196 34842
rect 37950 34788 37956 34790
rect 38012 34788 38036 34790
rect 38092 34788 38116 34790
rect 38172 34788 38196 34790
rect 38252 34788 38258 34790
rect 37950 34779 38258 34788
rect 37556 34740 37608 34746
rect 37556 34682 37608 34688
rect 38568 34604 38620 34610
rect 38568 34546 38620 34552
rect 37950 33756 38258 33765
rect 37950 33754 37956 33756
rect 38012 33754 38036 33756
rect 38092 33754 38116 33756
rect 38172 33754 38196 33756
rect 38252 33754 38258 33756
rect 38012 33702 38014 33754
rect 38194 33702 38196 33754
rect 37950 33700 37956 33702
rect 38012 33700 38036 33702
rect 38092 33700 38116 33702
rect 38172 33700 38196 33702
rect 38252 33700 38258 33702
rect 37950 33691 38258 33700
rect 37950 32668 38258 32677
rect 37950 32666 37956 32668
rect 38012 32666 38036 32668
rect 38092 32666 38116 32668
rect 38172 32666 38196 32668
rect 38252 32666 38258 32668
rect 38012 32614 38014 32666
rect 38194 32614 38196 32666
rect 37950 32612 37956 32614
rect 38012 32612 38036 32614
rect 38092 32612 38116 32614
rect 38172 32612 38196 32614
rect 38252 32612 38258 32614
rect 37950 32603 38258 32612
rect 37832 32292 37884 32298
rect 37832 32234 37884 32240
rect 37372 30252 37424 30258
rect 37372 30194 37424 30200
rect 36544 27940 36596 27946
rect 36544 27882 36596 27888
rect 37844 25906 37872 32234
rect 37950 31580 38258 31589
rect 37950 31578 37956 31580
rect 38012 31578 38036 31580
rect 38092 31578 38116 31580
rect 38172 31578 38196 31580
rect 38252 31578 38258 31580
rect 38012 31526 38014 31578
rect 38194 31526 38196 31578
rect 37950 31524 37956 31526
rect 38012 31524 38036 31526
rect 38092 31524 38116 31526
rect 38172 31524 38196 31526
rect 38252 31524 38258 31526
rect 37950 31515 38258 31524
rect 38580 31278 38608 34546
rect 38568 31272 38620 31278
rect 38568 31214 38620 31220
rect 37950 30492 38258 30501
rect 37950 30490 37956 30492
rect 38012 30490 38036 30492
rect 38092 30490 38116 30492
rect 38172 30490 38196 30492
rect 38252 30490 38258 30492
rect 38012 30438 38014 30490
rect 38194 30438 38196 30490
rect 37950 30436 37956 30438
rect 38012 30436 38036 30438
rect 38092 30436 38116 30438
rect 38172 30436 38196 30438
rect 38252 30436 38258 30438
rect 37950 30427 38258 30436
rect 37950 29404 38258 29413
rect 37950 29402 37956 29404
rect 38012 29402 38036 29404
rect 38092 29402 38116 29404
rect 38172 29402 38196 29404
rect 38252 29402 38258 29404
rect 38012 29350 38014 29402
rect 38194 29350 38196 29402
rect 37950 29348 37956 29350
rect 38012 29348 38036 29350
rect 38092 29348 38116 29350
rect 38172 29348 38196 29350
rect 38252 29348 38258 29350
rect 37950 29339 38258 29348
rect 37950 28316 38258 28325
rect 37950 28314 37956 28316
rect 38012 28314 38036 28316
rect 38092 28314 38116 28316
rect 38172 28314 38196 28316
rect 38252 28314 38258 28316
rect 38012 28262 38014 28314
rect 38194 28262 38196 28314
rect 37950 28260 37956 28262
rect 38012 28260 38036 28262
rect 38092 28260 38116 28262
rect 38172 28260 38196 28262
rect 38252 28260 38258 28262
rect 37950 28251 38258 28260
rect 37950 27228 38258 27237
rect 37950 27226 37956 27228
rect 38012 27226 38036 27228
rect 38092 27226 38116 27228
rect 38172 27226 38196 27228
rect 38252 27226 38258 27228
rect 38012 27174 38014 27226
rect 38194 27174 38196 27226
rect 37950 27172 37956 27174
rect 38012 27172 38036 27174
rect 38092 27172 38116 27174
rect 38172 27172 38196 27174
rect 38252 27172 38258 27174
rect 37950 27163 38258 27172
rect 37950 26140 38258 26149
rect 37950 26138 37956 26140
rect 38012 26138 38036 26140
rect 38092 26138 38116 26140
rect 38172 26138 38196 26140
rect 38252 26138 38258 26140
rect 38012 26086 38014 26138
rect 38194 26086 38196 26138
rect 37950 26084 37956 26086
rect 38012 26084 38036 26086
rect 38092 26084 38116 26086
rect 38172 26084 38196 26086
rect 38252 26084 38258 26086
rect 37950 26075 38258 26084
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 37950 25052 38258 25061
rect 37950 25050 37956 25052
rect 38012 25050 38036 25052
rect 38092 25050 38116 25052
rect 38172 25050 38196 25052
rect 38252 25050 38258 25052
rect 38012 24998 38014 25050
rect 38194 24998 38196 25050
rect 37950 24996 37956 24998
rect 38012 24996 38036 24998
rect 38092 24996 38116 24998
rect 38172 24996 38196 24998
rect 38252 24996 38258 24998
rect 37950 24987 38258 24996
rect 39316 24750 39344 38898
rect 39408 37194 39436 39918
rect 39396 37188 39448 37194
rect 39396 37130 39448 37136
rect 39500 35086 39528 41958
rect 39776 41414 39804 45494
rect 40144 44334 40172 46922
rect 42812 45490 42840 47398
rect 42950 47356 43258 47365
rect 42950 47354 42956 47356
rect 43012 47354 43036 47356
rect 43092 47354 43116 47356
rect 43172 47354 43196 47356
rect 43252 47354 43258 47356
rect 43012 47302 43014 47354
rect 43194 47302 43196 47354
rect 42950 47300 42956 47302
rect 43012 47300 43036 47302
rect 43092 47300 43116 47302
rect 43172 47300 43196 47302
rect 43252 47300 43258 47302
rect 42950 47291 43258 47300
rect 42950 46268 43258 46277
rect 42950 46266 42956 46268
rect 43012 46266 43036 46268
rect 43092 46266 43116 46268
rect 43172 46266 43196 46268
rect 43252 46266 43258 46268
rect 43012 46214 43014 46266
rect 43194 46214 43196 46266
rect 42950 46212 42956 46214
rect 43012 46212 43036 46214
rect 43092 46212 43116 46214
rect 43172 46212 43196 46214
rect 43252 46212 43258 46214
rect 42950 46203 43258 46212
rect 42800 45484 42852 45490
rect 42800 45426 42852 45432
rect 42950 45180 43258 45189
rect 42950 45178 42956 45180
rect 43012 45178 43036 45180
rect 43092 45178 43116 45180
rect 43172 45178 43196 45180
rect 43252 45178 43258 45180
rect 43012 45126 43014 45178
rect 43194 45126 43196 45178
rect 42950 45124 42956 45126
rect 43012 45124 43036 45126
rect 43092 45124 43116 45126
rect 43172 45124 43196 45126
rect 43252 45124 43258 45126
rect 42950 45115 43258 45124
rect 43364 44878 43392 47942
rect 43456 47054 43484 49710
rect 43444 47048 43496 47054
rect 43444 46990 43496 46996
rect 46216 45286 46244 52838
rect 48504 52488 48556 52494
rect 48504 52430 48556 52436
rect 47950 52252 48258 52261
rect 47950 52250 47956 52252
rect 48012 52250 48036 52252
rect 48092 52250 48116 52252
rect 48172 52250 48196 52252
rect 48252 52250 48258 52252
rect 48012 52198 48014 52250
rect 48194 52198 48196 52250
rect 47950 52196 47956 52198
rect 48012 52196 48036 52198
rect 48092 52196 48116 52198
rect 48172 52196 48196 52198
rect 48252 52196 48258 52198
rect 47950 52187 48258 52196
rect 48516 52193 48544 52430
rect 48502 52184 48558 52193
rect 48502 52119 48558 52128
rect 48504 51400 48556 51406
rect 48502 51368 48504 51377
rect 48556 51368 48558 51377
rect 48502 51303 48558 51312
rect 47950 51164 48258 51173
rect 47950 51162 47956 51164
rect 48012 51162 48036 51164
rect 48092 51162 48116 51164
rect 48172 51162 48196 51164
rect 48252 51162 48258 51164
rect 48012 51110 48014 51162
rect 48194 51110 48196 51162
rect 47950 51108 47956 51110
rect 48012 51108 48036 51110
rect 48092 51108 48116 51110
rect 48172 51108 48196 51110
rect 48252 51108 48258 51110
rect 47950 51099 48258 51108
rect 47950 50076 48258 50085
rect 47950 50074 47956 50076
rect 48012 50074 48036 50076
rect 48092 50074 48116 50076
rect 48172 50074 48196 50076
rect 48252 50074 48258 50076
rect 48012 50022 48014 50074
rect 48194 50022 48196 50074
rect 47950 50020 47956 50022
rect 48012 50020 48036 50022
rect 48092 50020 48116 50022
rect 48172 50020 48196 50022
rect 48252 50020 48258 50022
rect 47950 50011 48258 50020
rect 47950 48988 48258 48997
rect 47950 48986 47956 48988
rect 48012 48986 48036 48988
rect 48092 48986 48116 48988
rect 48172 48986 48196 48988
rect 48252 48986 48258 48988
rect 48012 48934 48014 48986
rect 48194 48934 48196 48986
rect 47950 48932 47956 48934
rect 48012 48932 48036 48934
rect 48092 48932 48116 48934
rect 48172 48932 48196 48934
rect 48252 48932 48258 48934
rect 47950 48923 48258 48932
rect 47950 47900 48258 47909
rect 47950 47898 47956 47900
rect 48012 47898 48036 47900
rect 48092 47898 48116 47900
rect 48172 47898 48196 47900
rect 48252 47898 48258 47900
rect 48012 47846 48014 47898
rect 48194 47846 48196 47898
rect 47950 47844 47956 47846
rect 48012 47844 48036 47846
rect 48092 47844 48116 47846
rect 48172 47844 48196 47846
rect 48252 47844 48258 47846
rect 47950 47835 48258 47844
rect 48700 47666 48728 53926
rect 48872 53440 48924 53446
rect 48872 53382 48924 53388
rect 48884 47734 48912 53382
rect 49252 52018 49280 56200
rect 49240 52012 49292 52018
rect 49240 51954 49292 51960
rect 49148 51808 49200 51814
rect 49148 51750 49200 51756
rect 49160 51474 49188 51750
rect 49148 51468 49200 51474
rect 49148 51410 49200 51416
rect 49332 50924 49384 50930
rect 49332 50866 49384 50872
rect 49344 50561 49372 50866
rect 49330 50552 49386 50561
rect 49330 50487 49386 50496
rect 49332 49836 49384 49842
rect 49332 49778 49384 49784
rect 49344 49745 49372 49778
rect 49330 49736 49386 49745
rect 49330 49671 49386 49680
rect 49056 49224 49108 49230
rect 49056 49166 49108 49172
rect 49068 48929 49096 49166
rect 49054 48920 49110 48929
rect 49054 48855 49110 48864
rect 49332 48136 49384 48142
rect 49330 48104 49332 48113
rect 49384 48104 49386 48113
rect 49330 48039 49386 48048
rect 48872 47728 48924 47734
rect 48872 47670 48924 47676
rect 48688 47660 48740 47666
rect 48688 47602 48740 47608
rect 49332 47660 49384 47666
rect 49332 47602 49384 47608
rect 49344 47297 49372 47602
rect 49330 47288 49386 47297
rect 49330 47223 49386 47232
rect 47950 46812 48258 46821
rect 47950 46810 47956 46812
rect 48012 46810 48036 46812
rect 48092 46810 48116 46812
rect 48172 46810 48196 46812
rect 48252 46810 48258 46812
rect 48012 46758 48014 46810
rect 48194 46758 48196 46810
rect 47950 46756 47956 46758
rect 48012 46756 48036 46758
rect 48092 46756 48116 46758
rect 48172 46756 48196 46758
rect 48252 46756 48258 46758
rect 47950 46747 48258 46756
rect 49056 46572 49108 46578
rect 49056 46514 49108 46520
rect 49068 46481 49096 46514
rect 49054 46472 49110 46481
rect 49054 46407 49110 46416
rect 49056 45960 49108 45966
rect 49056 45902 49108 45908
rect 48596 45824 48648 45830
rect 48596 45766 48648 45772
rect 47950 45724 48258 45733
rect 47950 45722 47956 45724
rect 48012 45722 48036 45724
rect 48092 45722 48116 45724
rect 48172 45722 48196 45724
rect 48252 45722 48258 45724
rect 48012 45670 48014 45722
rect 48194 45670 48196 45722
rect 47950 45668 47956 45670
rect 48012 45668 48036 45670
rect 48092 45668 48116 45670
rect 48172 45668 48196 45670
rect 48252 45668 48258 45670
rect 47950 45659 48258 45668
rect 46204 45280 46256 45286
rect 46204 45222 46256 45228
rect 47400 45008 47452 45014
rect 47400 44950 47452 44956
rect 43352 44872 43404 44878
rect 43352 44814 43404 44820
rect 40132 44328 40184 44334
rect 40132 44270 40184 44276
rect 39684 41386 39804 41414
rect 39684 39953 39712 41386
rect 39670 39944 39726 39953
rect 39670 39879 39726 39888
rect 40144 38865 40172 44270
rect 42950 44092 43258 44101
rect 42950 44090 42956 44092
rect 43012 44090 43036 44092
rect 43092 44090 43116 44092
rect 43172 44090 43196 44092
rect 43252 44090 43258 44092
rect 43012 44038 43014 44090
rect 43194 44038 43196 44090
rect 42950 44036 42956 44038
rect 43012 44036 43036 44038
rect 43092 44036 43116 44038
rect 43172 44036 43196 44038
rect 43252 44036 43258 44038
rect 42950 44027 43258 44036
rect 42950 43004 43258 43013
rect 42950 43002 42956 43004
rect 43012 43002 43036 43004
rect 43092 43002 43116 43004
rect 43172 43002 43196 43004
rect 43252 43002 43258 43004
rect 43012 42950 43014 43002
rect 43194 42950 43196 43002
rect 42950 42948 42956 42950
rect 43012 42948 43036 42950
rect 43092 42948 43116 42950
rect 43172 42948 43196 42950
rect 43252 42948 43258 42950
rect 42950 42939 43258 42948
rect 47216 42560 47268 42566
rect 47216 42502 47268 42508
rect 42950 41916 43258 41925
rect 42950 41914 42956 41916
rect 43012 41914 43036 41916
rect 43092 41914 43116 41916
rect 43172 41914 43196 41916
rect 43252 41914 43258 41916
rect 43012 41862 43014 41914
rect 43194 41862 43196 41914
rect 42950 41860 42956 41862
rect 43012 41860 43036 41862
rect 43092 41860 43116 41862
rect 43172 41860 43196 41862
rect 43252 41860 43258 41862
rect 42950 41851 43258 41860
rect 42950 40828 43258 40837
rect 42950 40826 42956 40828
rect 43012 40826 43036 40828
rect 43092 40826 43116 40828
rect 43172 40826 43196 40828
rect 43252 40826 43258 40828
rect 43012 40774 43014 40826
rect 43194 40774 43196 40826
rect 42950 40772 42956 40774
rect 43012 40772 43036 40774
rect 43092 40772 43116 40774
rect 43172 40772 43196 40774
rect 43252 40772 43258 40774
rect 42950 40763 43258 40772
rect 47228 40458 47256 42502
rect 47412 40730 47440 44950
rect 48608 44742 48636 45766
rect 49068 45665 49096 45902
rect 49054 45656 49110 45665
rect 49054 45591 49110 45600
rect 49056 44872 49108 44878
rect 49054 44840 49056 44849
rect 49108 44840 49110 44849
rect 49054 44775 49110 44784
rect 48596 44736 48648 44742
rect 48596 44678 48648 44684
rect 47950 44636 48258 44645
rect 47950 44634 47956 44636
rect 48012 44634 48036 44636
rect 48092 44634 48116 44636
rect 48172 44634 48196 44636
rect 48252 44634 48258 44636
rect 48012 44582 48014 44634
rect 48194 44582 48196 44634
rect 47950 44580 47956 44582
rect 48012 44580 48036 44582
rect 48092 44580 48116 44582
rect 48172 44580 48196 44582
rect 48252 44580 48258 44582
rect 47950 44571 48258 44580
rect 49332 44396 49384 44402
rect 49332 44338 49384 44344
rect 49344 44033 49372 44338
rect 49330 44024 49386 44033
rect 49240 43988 49292 43994
rect 49330 43959 49386 43968
rect 49240 43930 49292 43936
rect 47950 43548 48258 43557
rect 47950 43546 47956 43548
rect 48012 43546 48036 43548
rect 48092 43546 48116 43548
rect 48172 43546 48196 43548
rect 48252 43546 48258 43548
rect 48012 43494 48014 43546
rect 48194 43494 48196 43546
rect 47950 43492 47956 43494
rect 48012 43492 48036 43494
rect 48092 43492 48116 43494
rect 48172 43492 48196 43494
rect 48252 43492 48258 43494
rect 47950 43483 48258 43492
rect 49252 43450 49280 43930
rect 49240 43444 49292 43450
rect 49240 43386 49292 43392
rect 49148 43308 49200 43314
rect 49148 43250 49200 43256
rect 49160 43217 49188 43250
rect 49146 43208 49202 43217
rect 49146 43143 49202 43152
rect 49056 42696 49108 42702
rect 49056 42638 49108 42644
rect 47950 42460 48258 42469
rect 47950 42458 47956 42460
rect 48012 42458 48036 42460
rect 48092 42458 48116 42460
rect 48172 42458 48196 42460
rect 48252 42458 48258 42460
rect 48012 42406 48014 42458
rect 48194 42406 48196 42458
rect 47950 42404 47956 42406
rect 48012 42404 48036 42406
rect 48092 42404 48116 42406
rect 48172 42404 48196 42406
rect 48252 42404 48258 42406
rect 47950 42395 48258 42404
rect 49068 42401 49096 42638
rect 49054 42392 49110 42401
rect 49054 42327 49110 42336
rect 49056 41608 49108 41614
rect 49054 41576 49056 41585
rect 49108 41576 49110 41585
rect 49054 41511 49110 41520
rect 49240 41472 49292 41478
rect 49240 41414 49292 41420
rect 47950 41372 48258 41381
rect 47950 41370 47956 41372
rect 48012 41370 48036 41372
rect 48092 41370 48116 41372
rect 48172 41370 48196 41372
rect 48252 41370 48258 41372
rect 48012 41318 48014 41370
rect 48194 41318 48196 41370
rect 47950 41316 47956 41318
rect 48012 41316 48036 41318
rect 48092 41316 48116 41318
rect 48172 41316 48196 41318
rect 48252 41316 48258 41318
rect 47950 41307 48258 41316
rect 49148 40928 49200 40934
rect 49148 40870 49200 40876
rect 47400 40724 47452 40730
rect 47400 40666 47452 40672
rect 49160 40526 49188 40870
rect 49148 40520 49200 40526
rect 49148 40462 49200 40468
rect 47216 40452 47268 40458
rect 47216 40394 47268 40400
rect 47950 40284 48258 40293
rect 47950 40282 47956 40284
rect 48012 40282 48036 40284
rect 48092 40282 48116 40284
rect 48172 40282 48196 40284
rect 48252 40282 48258 40284
rect 48012 40230 48014 40282
rect 48194 40230 48196 40282
rect 47950 40228 47956 40230
rect 48012 40228 48036 40230
rect 48092 40228 48116 40230
rect 48172 40228 48196 40230
rect 48252 40228 48258 40230
rect 47950 40219 48258 40228
rect 49056 40044 49108 40050
rect 49056 39986 49108 39992
rect 49068 39953 49096 39986
rect 49054 39944 49110 39953
rect 49054 39879 49110 39888
rect 42950 39740 43258 39749
rect 42950 39738 42956 39740
rect 43012 39738 43036 39740
rect 43092 39738 43116 39740
rect 43172 39738 43196 39740
rect 43252 39738 43258 39740
rect 43012 39686 43014 39738
rect 43194 39686 43196 39738
rect 42950 39684 42956 39686
rect 43012 39684 43036 39686
rect 43092 39684 43116 39686
rect 43172 39684 43196 39686
rect 43252 39684 43258 39686
rect 42950 39675 43258 39684
rect 41328 39568 41380 39574
rect 41328 39510 41380 39516
rect 40130 38856 40186 38865
rect 40130 38791 40186 38800
rect 39672 38480 39724 38486
rect 39672 38422 39724 38428
rect 39488 35080 39540 35086
rect 39488 35022 39540 35028
rect 39684 33522 39712 38422
rect 39856 37664 39908 37670
rect 39856 37606 39908 37612
rect 39868 33522 39896 37606
rect 39948 35488 40000 35494
rect 39948 35430 40000 35436
rect 39672 33516 39724 33522
rect 39672 33458 39724 33464
rect 39856 33516 39908 33522
rect 39856 33458 39908 33464
rect 39960 31414 39988 35430
rect 41340 34610 41368 39510
rect 49252 39438 49280 41414
rect 49332 41132 49384 41138
rect 49332 41074 49384 41080
rect 49344 40769 49372 41074
rect 49330 40760 49386 40769
rect 49330 40695 49386 40704
rect 49240 39432 49292 39438
rect 49240 39374 49292 39380
rect 49148 39364 49200 39370
rect 49148 39306 49200 39312
rect 47950 39196 48258 39205
rect 47950 39194 47956 39196
rect 48012 39194 48036 39196
rect 48092 39194 48116 39196
rect 48172 39194 48196 39196
rect 48252 39194 48258 39196
rect 48012 39142 48014 39194
rect 48194 39142 48196 39194
rect 47950 39140 47956 39142
rect 48012 39140 48036 39142
rect 48092 39140 48116 39142
rect 48172 39140 48196 39142
rect 48252 39140 48258 39142
rect 47950 39131 48258 39140
rect 49160 39137 49188 39306
rect 49240 39296 49292 39302
rect 49240 39238 49292 39244
rect 49146 39128 49202 39137
rect 49146 39063 49202 39072
rect 49252 38962 49280 39238
rect 49240 38956 49292 38962
rect 49240 38898 49292 38904
rect 42950 38652 43258 38661
rect 42950 38650 42956 38652
rect 43012 38650 43036 38652
rect 43092 38650 43116 38652
rect 43172 38650 43196 38652
rect 43252 38650 43258 38652
rect 43012 38598 43014 38650
rect 43194 38598 43196 38650
rect 42950 38596 42956 38598
rect 43012 38596 43036 38598
rect 43092 38596 43116 38598
rect 43172 38596 43196 38598
rect 43252 38596 43258 38598
rect 42950 38587 43258 38596
rect 49146 38312 49202 38321
rect 49146 38247 49148 38256
rect 49200 38247 49202 38256
rect 49148 38218 49200 38224
rect 49240 38208 49292 38214
rect 49240 38150 49292 38156
rect 47950 38108 48258 38117
rect 47950 38106 47956 38108
rect 48012 38106 48036 38108
rect 48092 38106 48116 38108
rect 48172 38106 48196 38108
rect 48252 38106 48258 38108
rect 48012 38054 48014 38106
rect 48194 38054 48196 38106
rect 47950 38052 47956 38054
rect 48012 38052 48036 38054
rect 48092 38052 48116 38054
rect 48172 38052 48196 38054
rect 48252 38052 48258 38054
rect 47950 38043 48258 38052
rect 49252 37942 49280 38150
rect 49240 37936 49292 37942
rect 49240 37878 49292 37884
rect 49332 37868 49384 37874
rect 49332 37810 49384 37816
rect 42950 37564 43258 37573
rect 42950 37562 42956 37564
rect 43012 37562 43036 37564
rect 43092 37562 43116 37564
rect 43172 37562 43196 37564
rect 43252 37562 43258 37564
rect 43012 37510 43014 37562
rect 43194 37510 43196 37562
rect 42950 37508 42956 37510
rect 43012 37508 43036 37510
rect 43092 37508 43116 37510
rect 43172 37508 43196 37510
rect 43252 37508 43258 37510
rect 42950 37499 43258 37508
rect 49344 37505 49372 37810
rect 49330 37496 49386 37505
rect 49330 37431 49386 37440
rect 47950 37020 48258 37029
rect 47950 37018 47956 37020
rect 48012 37018 48036 37020
rect 48092 37018 48116 37020
rect 48172 37018 48196 37020
rect 48252 37018 48258 37020
rect 48012 36966 48014 37018
rect 48194 36966 48196 37018
rect 47950 36964 47956 36966
rect 48012 36964 48036 36966
rect 48092 36964 48116 36966
rect 48172 36964 48196 36966
rect 48252 36964 48258 36966
rect 47950 36955 48258 36964
rect 49240 36848 49292 36854
rect 49240 36790 49292 36796
rect 47400 36780 47452 36786
rect 47400 36722 47452 36728
rect 49056 36780 49108 36786
rect 49056 36722 49108 36728
rect 42950 36476 43258 36485
rect 42950 36474 42956 36476
rect 43012 36474 43036 36476
rect 43092 36474 43116 36476
rect 43172 36474 43196 36476
rect 43252 36474 43258 36476
rect 43012 36422 43014 36474
rect 43194 36422 43196 36474
rect 42950 36420 42956 36422
rect 43012 36420 43036 36422
rect 43092 36420 43116 36422
rect 43172 36420 43196 36422
rect 43252 36420 43258 36422
rect 42950 36411 43258 36420
rect 42950 35388 43258 35397
rect 42950 35386 42956 35388
rect 43012 35386 43036 35388
rect 43092 35386 43116 35388
rect 43172 35386 43196 35388
rect 43252 35386 43258 35388
rect 43012 35334 43014 35386
rect 43194 35334 43196 35386
rect 42950 35332 42956 35334
rect 43012 35332 43036 35334
rect 43092 35332 43116 35334
rect 43172 35332 43196 35334
rect 43252 35332 43258 35334
rect 42950 35323 43258 35332
rect 42616 34944 42668 34950
rect 42616 34886 42668 34892
rect 41328 34604 41380 34610
rect 41328 34546 41380 34552
rect 39948 31408 40000 31414
rect 39948 31350 40000 31356
rect 42628 30734 42656 34886
rect 47412 34746 47440 36722
rect 49068 36689 49096 36722
rect 48318 36680 48374 36689
rect 48318 36615 48320 36624
rect 48372 36615 48374 36624
rect 49054 36680 49110 36689
rect 49054 36615 49110 36624
rect 48320 36586 48372 36592
rect 49252 36378 49280 36790
rect 49240 36372 49292 36378
rect 49240 36314 49292 36320
rect 48320 36168 48372 36174
rect 48320 36110 48372 36116
rect 47950 35932 48258 35941
rect 47950 35930 47956 35932
rect 48012 35930 48036 35932
rect 48092 35930 48116 35932
rect 48172 35930 48196 35932
rect 48252 35930 48258 35932
rect 48012 35878 48014 35930
rect 48194 35878 48196 35930
rect 47950 35876 47956 35878
rect 48012 35876 48036 35878
rect 48092 35876 48116 35878
rect 48172 35876 48196 35878
rect 48252 35876 48258 35878
rect 47950 35867 48258 35876
rect 48332 35894 48360 36110
rect 48332 35873 48452 35894
rect 48332 35866 48466 35873
rect 48410 35864 48466 35866
rect 48410 35799 48466 35808
rect 49056 35080 49108 35086
rect 48318 35048 48374 35057
rect 48318 34983 48374 34992
rect 49054 35048 49056 35057
rect 49108 35048 49110 35057
rect 49054 34983 49110 34992
rect 48332 34950 48360 34983
rect 48320 34944 48372 34950
rect 48320 34886 48372 34892
rect 47950 34844 48258 34853
rect 47950 34842 47956 34844
rect 48012 34842 48036 34844
rect 48092 34842 48116 34844
rect 48172 34842 48196 34844
rect 48252 34842 48258 34844
rect 48012 34790 48014 34842
rect 48194 34790 48196 34842
rect 47950 34788 47956 34790
rect 48012 34788 48036 34790
rect 48092 34788 48116 34790
rect 48172 34788 48196 34790
rect 48252 34788 48258 34790
rect 47950 34779 48258 34788
rect 44180 34740 44232 34746
rect 44180 34682 44232 34688
rect 47400 34740 47452 34746
rect 47400 34682 47452 34688
rect 42950 34300 43258 34309
rect 42950 34298 42956 34300
rect 43012 34298 43036 34300
rect 43092 34298 43116 34300
rect 43172 34298 43196 34300
rect 43252 34298 43258 34300
rect 43012 34246 43014 34298
rect 43194 34246 43196 34298
rect 42950 34244 42956 34246
rect 43012 34244 43036 34246
rect 43092 34244 43116 34246
rect 43172 34244 43196 34246
rect 43252 34244 43258 34246
rect 42950 34235 43258 34244
rect 44088 33380 44140 33386
rect 44088 33322 44140 33328
rect 42950 33212 43258 33221
rect 42950 33210 42956 33212
rect 43012 33210 43036 33212
rect 43092 33210 43116 33212
rect 43172 33210 43196 33212
rect 43252 33210 43258 33212
rect 43012 33158 43014 33210
rect 43194 33158 43196 33210
rect 42950 33156 42956 33158
rect 43012 33156 43036 33158
rect 43092 33156 43116 33158
rect 43172 33156 43196 33158
rect 43252 33156 43258 33158
rect 42950 33147 43258 33156
rect 42950 32124 43258 32133
rect 42950 32122 42956 32124
rect 43012 32122 43036 32124
rect 43092 32122 43116 32124
rect 43172 32122 43196 32124
rect 43252 32122 43258 32124
rect 43012 32070 43014 32122
rect 43194 32070 43196 32122
rect 42950 32068 42956 32070
rect 43012 32068 43036 32070
rect 43092 32068 43116 32070
rect 43172 32068 43196 32070
rect 43252 32068 43258 32070
rect 42950 32059 43258 32068
rect 42950 31036 43258 31045
rect 42950 31034 42956 31036
rect 43012 31034 43036 31036
rect 43092 31034 43116 31036
rect 43172 31034 43196 31036
rect 43252 31034 43258 31036
rect 43012 30982 43014 31034
rect 43194 30982 43196 31034
rect 42950 30980 42956 30982
rect 43012 30980 43036 30982
rect 43092 30980 43116 30982
rect 43172 30980 43196 30982
rect 43252 30980 43258 30982
rect 42950 30971 43258 30980
rect 42616 30728 42668 30734
rect 42616 30670 42668 30676
rect 40132 30388 40184 30394
rect 40132 30330 40184 30336
rect 39396 30048 39448 30054
rect 39396 29990 39448 29996
rect 39304 24744 39356 24750
rect 39304 24686 39356 24692
rect 39408 24206 39436 29990
rect 39948 25696 40000 25702
rect 39948 25638 40000 25644
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 33416 23792 33468 23798
rect 33416 23734 33468 23740
rect 33428 18698 33456 23734
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 33416 18692 33468 18698
rect 33416 18634 33468 18640
rect 36740 15094 36768 23462
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 39960 19446 39988 25638
rect 39948 19440 40000 19446
rect 39948 19382 40000 19388
rect 40144 18766 40172 30330
rect 42950 29948 43258 29957
rect 42950 29946 42956 29948
rect 43012 29946 43036 29948
rect 43092 29946 43116 29948
rect 43172 29946 43196 29948
rect 43252 29946 43258 29948
rect 43012 29894 43014 29946
rect 43194 29894 43196 29946
rect 42950 29892 42956 29894
rect 43012 29892 43036 29894
rect 43092 29892 43116 29894
rect 43172 29892 43196 29894
rect 43252 29892 43258 29894
rect 42950 29883 43258 29892
rect 42950 28860 43258 28869
rect 42950 28858 42956 28860
rect 43012 28858 43036 28860
rect 43092 28858 43116 28860
rect 43172 28858 43196 28860
rect 43252 28858 43258 28860
rect 43012 28806 43014 28858
rect 43194 28806 43196 28858
rect 42950 28804 42956 28806
rect 43012 28804 43036 28806
rect 43092 28804 43116 28806
rect 43172 28804 43196 28806
rect 43252 28804 43258 28806
rect 42950 28795 43258 28804
rect 43904 28416 43956 28422
rect 43904 28358 43956 28364
rect 42950 27772 43258 27781
rect 42950 27770 42956 27772
rect 43012 27770 43036 27772
rect 43092 27770 43116 27772
rect 43172 27770 43196 27772
rect 43252 27770 43258 27772
rect 43012 27718 43014 27770
rect 43194 27718 43196 27770
rect 42950 27716 42956 27718
rect 43012 27716 43036 27718
rect 43092 27716 43116 27718
rect 43172 27716 43196 27718
rect 43252 27716 43258 27718
rect 42950 27707 43258 27716
rect 42950 26684 43258 26693
rect 42950 26682 42956 26684
rect 43012 26682 43036 26684
rect 43092 26682 43116 26684
rect 43172 26682 43196 26684
rect 43252 26682 43258 26684
rect 43012 26630 43014 26682
rect 43194 26630 43196 26682
rect 42950 26628 42956 26630
rect 43012 26628 43036 26630
rect 43092 26628 43116 26630
rect 43172 26628 43196 26630
rect 43252 26628 43258 26630
rect 42950 26619 43258 26628
rect 42950 25596 43258 25605
rect 42950 25594 42956 25596
rect 43012 25594 43036 25596
rect 43092 25594 43116 25596
rect 43172 25594 43196 25596
rect 43252 25594 43258 25596
rect 43012 25542 43014 25594
rect 43194 25542 43196 25594
rect 42950 25540 42956 25542
rect 43012 25540 43036 25542
rect 43092 25540 43116 25542
rect 43172 25540 43196 25542
rect 43252 25540 43258 25542
rect 42950 25531 43258 25540
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 43444 24064 43496 24070
rect 43444 24006 43496 24012
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42800 21412 42852 21418
rect 42800 21354 42852 21360
rect 40132 18760 40184 18766
rect 40132 18702 40184 18708
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 42812 17202 42840 21354
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 43352 17604 43404 17610
rect 43352 17546 43404 17552
rect 42800 17196 42852 17202
rect 42800 17138 42852 17144
rect 38292 17060 38344 17066
rect 38292 17002 38344 17008
rect 38304 16574 38332 17002
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 38568 16652 38620 16658
rect 38568 16594 38620 16600
rect 37844 16546 38332 16574
rect 36728 15088 36780 15094
rect 36728 15030 36780 15036
rect 37740 13864 37792 13870
rect 37740 13806 37792 13812
rect 37464 11076 37516 11082
rect 37464 11018 37516 11024
rect 33324 9988 33376 9994
rect 33324 9930 33376 9936
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 33336 8634 33364 9930
rect 36452 9444 36504 9450
rect 36452 9386 36504 9392
rect 33324 8628 33376 8634
rect 33324 8570 33376 8576
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 30748 7404 30800 7410
rect 30748 7346 30800 7352
rect 29828 2508 29880 2514
rect 29828 2450 29880 2456
rect 30760 2106 30788 7346
rect 34440 7206 34468 8230
rect 34428 7200 34480 7206
rect 34428 7142 34480 7148
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 34440 2650 34468 7142
rect 36464 3534 36492 9386
rect 37476 5234 37504 11018
rect 37752 8498 37780 13806
rect 37844 11762 37872 16546
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 38580 16130 38608 16594
rect 38304 16102 38608 16130
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 37832 11756 37884 11762
rect 37832 11698 37884 11704
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 38304 10674 38332 16102
rect 38476 15972 38528 15978
rect 38476 15914 38528 15920
rect 38384 12640 38436 12646
rect 38384 12582 38436 12588
rect 38292 10668 38344 10674
rect 38292 10610 38344 10616
rect 37832 10532 37884 10538
rect 37832 10474 37884 10480
rect 37740 8492 37792 8498
rect 37740 8434 37792 8440
rect 37464 5228 37516 5234
rect 37464 5170 37516 5176
rect 37844 4146 37872 10474
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 38396 6798 38424 12582
rect 38488 10062 38516 15914
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 43364 13326 43392 17546
rect 43456 16590 43484 24006
rect 43916 22030 43944 28358
rect 44100 28150 44128 33322
rect 44192 29510 44220 34682
rect 49332 34604 49384 34610
rect 49332 34546 49384 34552
rect 49344 34241 49372 34546
rect 49330 34232 49386 34241
rect 49330 34167 49386 34176
rect 47950 33756 48258 33765
rect 47950 33754 47956 33756
rect 48012 33754 48036 33756
rect 48092 33754 48116 33756
rect 48172 33754 48196 33756
rect 48252 33754 48258 33756
rect 48012 33702 48014 33754
rect 48194 33702 48196 33754
rect 47950 33700 47956 33702
rect 48012 33700 48036 33702
rect 48092 33700 48116 33702
rect 48172 33700 48196 33702
rect 48252 33700 48258 33702
rect 47950 33691 48258 33700
rect 49148 33516 49200 33522
rect 49148 33458 49200 33464
rect 49160 33425 49188 33458
rect 49146 33416 49202 33425
rect 49146 33351 49202 33360
rect 45836 33312 45888 33318
rect 45836 33254 45888 33260
rect 44548 31136 44600 31142
rect 44548 31078 44600 31084
rect 44180 29504 44232 29510
rect 44180 29446 44232 29452
rect 44088 28144 44140 28150
rect 44088 28086 44140 28092
rect 44560 27062 44588 31078
rect 45848 29578 45876 33254
rect 49056 32904 49108 32910
rect 49056 32846 49108 32852
rect 47950 32668 48258 32677
rect 47950 32666 47956 32668
rect 48012 32666 48036 32668
rect 48092 32666 48116 32668
rect 48172 32666 48196 32668
rect 48252 32666 48258 32668
rect 48012 32614 48014 32666
rect 48194 32614 48196 32666
rect 47950 32612 47956 32614
rect 48012 32612 48036 32614
rect 48092 32612 48116 32614
rect 48172 32612 48196 32614
rect 48252 32612 48258 32614
rect 47950 32603 48258 32612
rect 49068 32609 49096 32846
rect 49054 32600 49110 32609
rect 49054 32535 49110 32544
rect 49056 31816 49108 31822
rect 49054 31784 49056 31793
rect 49108 31784 49110 31793
rect 49054 31719 49110 31728
rect 47950 31580 48258 31589
rect 47950 31578 47956 31580
rect 48012 31578 48036 31580
rect 48092 31578 48116 31580
rect 48172 31578 48196 31580
rect 48252 31578 48258 31580
rect 48012 31526 48014 31578
rect 48194 31526 48196 31578
rect 47950 31524 47956 31526
rect 48012 31524 48036 31526
rect 48092 31524 48116 31526
rect 48172 31524 48196 31526
rect 48252 31524 48258 31526
rect 47950 31515 48258 31524
rect 49332 31340 49384 31346
rect 49332 31282 49384 31288
rect 46756 31204 46808 31210
rect 46756 31146 46808 31152
rect 46480 30660 46532 30666
rect 46480 30602 46532 30608
rect 45836 29572 45888 29578
rect 45836 29514 45888 29520
rect 45928 29504 45980 29510
rect 45928 29446 45980 29452
rect 45284 27872 45336 27878
rect 45284 27814 45336 27820
rect 44548 27056 44600 27062
rect 44548 26998 44600 27004
rect 44732 26852 44784 26858
rect 44732 26794 44784 26800
rect 44272 25764 44324 25770
rect 44272 25706 44324 25712
rect 44180 24676 44232 24682
rect 44180 24618 44232 24624
rect 43904 22024 43956 22030
rect 43904 21966 43956 21972
rect 44192 20466 44220 24618
rect 44284 21554 44312 25706
rect 44744 22030 44772 26794
rect 45100 24132 45152 24138
rect 45100 24074 45152 24080
rect 44732 22024 44784 22030
rect 44732 21966 44784 21972
rect 44824 21956 44876 21962
rect 44824 21898 44876 21904
rect 44272 21548 44324 21554
rect 44272 21490 44324 21496
rect 44180 20460 44232 20466
rect 44180 20402 44232 20408
rect 44272 19236 44324 19242
rect 44272 19178 44324 19184
rect 43444 16584 43496 16590
rect 43444 16526 43496 16532
rect 44284 15026 44312 19178
rect 44836 15502 44864 21898
rect 45112 18766 45140 24074
rect 45296 23118 45324 27814
rect 45940 25294 45968 29446
rect 46492 26382 46520 30602
rect 46768 26994 46796 31146
rect 49344 30977 49372 31282
rect 49330 30968 49386 30977
rect 49330 30903 49386 30912
rect 47950 30492 48258 30501
rect 47950 30490 47956 30492
rect 48012 30490 48036 30492
rect 48092 30490 48116 30492
rect 48172 30490 48196 30492
rect 48252 30490 48258 30492
rect 48012 30438 48014 30490
rect 48194 30438 48196 30490
rect 47950 30436 47956 30438
rect 48012 30436 48036 30438
rect 48092 30436 48116 30438
rect 48172 30436 48196 30438
rect 48252 30436 48258 30438
rect 47950 30427 48258 30436
rect 49056 30252 49108 30258
rect 49056 30194 49108 30200
rect 49068 30161 49096 30194
rect 49054 30152 49110 30161
rect 49054 30087 49110 30096
rect 49240 30048 49292 30054
rect 49240 29990 49292 29996
rect 49252 29850 49280 29990
rect 49240 29844 49292 29850
rect 49240 29786 49292 29792
rect 47768 29572 47820 29578
rect 47768 29514 47820 29520
rect 49148 29572 49200 29578
rect 49148 29514 49200 29520
rect 46848 27396 46900 27402
rect 46848 27338 46900 27344
rect 46756 26988 46808 26994
rect 46756 26930 46808 26936
rect 46480 26376 46532 26382
rect 46480 26318 46532 26324
rect 45928 25288 45980 25294
rect 45928 25230 45980 25236
rect 46860 23730 46888 27338
rect 47780 24818 47808 29514
rect 47950 29404 48258 29413
rect 47950 29402 47956 29404
rect 48012 29402 48036 29404
rect 48092 29402 48116 29404
rect 48172 29402 48196 29404
rect 48252 29402 48258 29404
rect 48012 29350 48014 29402
rect 48194 29350 48196 29402
rect 47950 29348 47956 29350
rect 48012 29348 48036 29350
rect 48092 29348 48116 29350
rect 48172 29348 48196 29350
rect 48252 29348 48258 29350
rect 47950 29339 48258 29348
rect 49160 29345 49188 29514
rect 49146 29336 49202 29345
rect 49146 29271 49202 29280
rect 49056 28552 49108 28558
rect 49054 28520 49056 28529
rect 49108 28520 49110 28529
rect 49054 28455 49110 28464
rect 47950 28316 48258 28325
rect 47950 28314 47956 28316
rect 48012 28314 48036 28316
rect 48092 28314 48116 28316
rect 48172 28314 48196 28316
rect 48252 28314 48258 28316
rect 48012 28262 48014 28314
rect 48194 28262 48196 28314
rect 47950 28260 47956 28262
rect 48012 28260 48036 28262
rect 48092 28260 48116 28262
rect 48172 28260 48196 28262
rect 48252 28260 48258 28262
rect 47950 28251 48258 28260
rect 49332 28076 49384 28082
rect 49332 28018 49384 28024
rect 49344 27713 49372 28018
rect 49330 27704 49386 27713
rect 49330 27639 49386 27648
rect 47950 27228 48258 27237
rect 47950 27226 47956 27228
rect 48012 27226 48036 27228
rect 48092 27226 48116 27228
rect 48172 27226 48196 27228
rect 48252 27226 48258 27228
rect 48012 27174 48014 27226
rect 48194 27174 48196 27226
rect 47950 27172 47956 27174
rect 48012 27172 48036 27174
rect 48092 27172 48116 27174
rect 48172 27172 48196 27174
rect 48252 27172 48258 27174
rect 47950 27163 48258 27172
rect 49148 26920 49200 26926
rect 49146 26888 49148 26897
rect 49200 26888 49202 26897
rect 49146 26823 49202 26832
rect 48228 26444 48280 26450
rect 48228 26386 48280 26392
rect 48240 26234 48268 26386
rect 48240 26206 48360 26234
rect 47950 26140 48258 26149
rect 47950 26138 47956 26140
rect 48012 26138 48036 26140
rect 48092 26138 48116 26140
rect 48172 26138 48196 26140
rect 48252 26138 48258 26140
rect 48012 26086 48014 26138
rect 48194 26086 48196 26138
rect 47950 26084 47956 26086
rect 48012 26084 48036 26086
rect 48092 26084 48116 26086
rect 48172 26084 48196 26086
rect 48252 26084 48258 26086
rect 47950 26075 48258 26084
rect 48332 26058 48360 26206
rect 48410 26072 48466 26081
rect 48332 26030 48410 26058
rect 48410 26007 48466 26016
rect 49148 25288 49200 25294
rect 49146 25256 49148 25265
rect 49200 25256 49202 25265
rect 49146 25191 49202 25200
rect 47950 25052 48258 25061
rect 47950 25050 47956 25052
rect 48012 25050 48036 25052
rect 48092 25050 48116 25052
rect 48172 25050 48196 25052
rect 48252 25050 48258 25052
rect 48012 24998 48014 25050
rect 48194 24998 48196 25050
rect 47950 24996 47956 24998
rect 48012 24996 48036 24998
rect 48092 24996 48116 24998
rect 48172 24996 48196 24998
rect 48252 24996 48258 24998
rect 47950 24987 48258 24996
rect 47768 24812 47820 24818
rect 47768 24754 47820 24760
rect 49148 24744 49200 24750
rect 49148 24686 49200 24692
rect 46940 24608 46992 24614
rect 46940 24550 46992 24556
rect 46848 23724 46900 23730
rect 46848 23666 46900 23672
rect 45284 23112 45336 23118
rect 45284 23054 45336 23060
rect 46952 19854 46980 24550
rect 49160 24449 49188 24686
rect 49146 24440 49202 24449
rect 49146 24375 49202 24384
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 49148 23656 49200 23662
rect 49146 23624 49148 23633
rect 49200 23624 49202 23633
rect 47032 23588 47084 23594
rect 49146 23559 49202 23568
rect 47032 23530 47084 23536
rect 46940 19848 46992 19854
rect 46940 19790 46992 19796
rect 46940 19236 46992 19242
rect 46940 19178 46992 19184
rect 45100 18760 45152 18766
rect 45100 18702 45152 18708
rect 46204 16652 46256 16658
rect 46204 16594 46256 16600
rect 44824 15496 44876 15502
rect 44824 15438 44876 15444
rect 44272 15020 44324 15026
rect 44272 14962 44324 14968
rect 43812 14816 43864 14822
rect 43812 14758 43864 14764
rect 43352 13320 43404 13326
rect 43352 13262 43404 13268
rect 38568 13252 38620 13258
rect 38568 13194 38620 13200
rect 38476 10056 38528 10062
rect 38476 9998 38528 10004
rect 38580 7410 38608 13194
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 38568 7404 38620 7410
rect 38568 7346 38620 7352
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 38384 6792 38436 6798
rect 38384 6734 38436 6740
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43824 5710 43852 14758
rect 46216 8974 46244 16594
rect 46952 12238 46980 19178
rect 47044 18290 47072 23530
rect 49148 23044 49200 23050
rect 49148 22986 49200 22992
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 49160 22817 49188 22986
rect 49146 22808 49202 22817
rect 49146 22743 49202 22752
rect 49148 22024 49200 22030
rect 49146 21992 49148 22001
rect 49200 21992 49202 22001
rect 49146 21927 49202 21936
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21185 49188 21422
rect 49146 21176 49202 21185
rect 49146 21111 49202 21120
rect 47768 20868 47820 20874
rect 47768 20810 47820 20816
rect 47032 18284 47084 18290
rect 47032 18226 47084 18232
rect 47780 16590 47808 20810
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 49148 20392 49200 20398
rect 49146 20360 49148 20369
rect 49200 20360 49202 20369
rect 49146 20295 49202 20304
rect 49148 19780 49200 19786
rect 49148 19722 49200 19728
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 49160 19553 49188 19722
rect 49146 19544 49202 19553
rect 49146 19479 49202 19488
rect 49148 18760 49200 18766
rect 49146 18728 49148 18737
rect 49200 18728 49202 18737
rect 47860 18692 47912 18698
rect 49146 18663 49202 18672
rect 47860 18634 47912 18640
rect 47768 16584 47820 16590
rect 47768 16526 47820 16532
rect 47872 13938 47900 18634
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 49148 18216 49200 18222
rect 49148 18158 49200 18164
rect 49160 17921 49188 18158
rect 49146 17912 49202 17921
rect 49146 17847 49202 17856
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 49148 17128 49200 17134
rect 49146 17096 49148 17105
rect 49200 17096 49202 17105
rect 49146 17031 49202 17040
rect 49148 16516 49200 16522
rect 49148 16458 49200 16464
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 49160 16289 49188 16458
rect 49146 16280 49202 16289
rect 49146 16215 49202 16224
rect 49148 15496 49200 15502
rect 49146 15464 49148 15473
rect 49200 15464 49202 15473
rect 49146 15399 49202 15408
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 49148 14952 49200 14958
rect 49148 14894 49200 14900
rect 49160 14657 49188 14894
rect 49146 14648 49202 14657
rect 49146 14583 49202 14592
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47860 13932 47912 13938
rect 47860 13874 47912 13880
rect 49148 13864 49200 13870
rect 49146 13832 49148 13841
rect 49200 13832 49202 13841
rect 49146 13767 49202 13776
rect 49148 13252 49200 13258
rect 49148 13194 49200 13200
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 49160 13025 49188 13194
rect 49146 13016 49202 13025
rect 49146 12951 49202 12960
rect 46940 12232 46992 12238
rect 49148 12232 49200 12238
rect 46940 12174 46992 12180
rect 49146 12200 49148 12209
rect 49200 12200 49202 12209
rect 49146 12135 49202 12144
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 49148 11688 49200 11694
rect 49148 11630 49200 11636
rect 49160 11393 49188 11630
rect 49146 11384 49202 11393
rect 49146 11319 49202 11328
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 49148 10600 49200 10606
rect 49146 10568 49148 10577
rect 49200 10568 49202 10577
rect 49146 10503 49202 10512
rect 49148 9988 49200 9994
rect 49148 9930 49200 9936
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 49160 9761 49188 9930
rect 49146 9752 49202 9761
rect 49146 9687 49202 9696
rect 46204 8968 46256 8974
rect 49148 8968 49200 8974
rect 46204 8910 46256 8916
rect 49146 8936 49148 8945
rect 49200 8936 49202 8945
rect 49146 8871 49202 8880
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 49148 8424 49200 8430
rect 49148 8366 49200 8372
rect 49160 8129 49188 8366
rect 49146 8120 49202 8129
rect 49146 8055 49202 8064
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49148 7336 49200 7342
rect 49146 7304 49148 7313
rect 49200 7304 49202 7313
rect 49146 7239 49202 7248
rect 49148 6724 49200 6730
rect 49148 6666 49200 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 49160 6497 49188 6666
rect 49146 6488 49202 6497
rect 49146 6423 49202 6432
rect 43812 5704 43864 5710
rect 49148 5704 49200 5710
rect 43812 5646 43864 5652
rect 49146 5672 49148 5681
rect 49200 5672 49202 5681
rect 49146 5607 49202 5616
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49148 5160 49200 5166
rect 49148 5102 49200 5108
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 49160 4865 49188 5102
rect 49146 4856 49202 4865
rect 49146 4791 49202 4800
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 49148 4072 49200 4078
rect 49146 4040 49148 4049
rect 49200 4040 49202 4049
rect 49146 3975 49202 3984
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 36452 3528 36504 3534
rect 36452 3470 36504 3476
rect 48596 3460 48648 3466
rect 48596 3402 48648 3408
rect 49148 3460 49200 3466
rect 49148 3402 49200 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 34428 2644 34480 2650
rect 34428 2586 34480 2592
rect 32036 2440 32088 2446
rect 32036 2382 32088 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 30748 2100 30800 2106
rect 30748 2042 30800 2048
rect 32048 800 32076 2382
rect 35360 800 35388 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38672 800 38700 2382
rect 41984 800 42012 2382
rect 45284 2372 45336 2378
rect 45284 2314 45336 2320
rect 45296 800 45324 2314
rect 45560 2304 45612 2310
rect 45560 2246 45612 2252
rect 45572 2106 45600 2246
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 45560 2100 45612 2106
rect 45560 2042 45612 2048
rect 48608 800 48636 3402
rect 49160 3233 49188 3402
rect 49146 3224 49202 3233
rect 49146 3159 49202 3168
rect 49146 2408 49202 2417
rect 49146 2343 49148 2352
rect 49200 2343 49202 2352
rect 49148 2314 49200 2320
rect 2226 0 2282 800
rect 5538 0 5594 800
rect 8850 0 8906 800
rect 12162 0 12218 800
rect 15474 0 15530 800
rect 18786 0 18842 800
rect 22098 0 22154 800
rect 25410 0 25466 800
rect 28722 0 28778 800
rect 32034 0 32090 800
rect 35346 0 35402 800
rect 38658 0 38714 800
rect 41970 0 42026 800
rect 45282 0 45338 800
rect 48594 0 48650 800
<< via2 >>
rect 1306 51312 1362 51368
rect 1306 50496 1362 50552
rect 1306 49716 1308 49736
rect 1308 49716 1360 49736
rect 1360 49716 1362 49736
rect 1306 49680 1362 49716
rect 1306 48864 1362 48920
rect 1306 48048 1362 48104
rect 1306 47232 1362 47288
rect 1306 46452 1308 46472
rect 1308 46452 1360 46472
rect 1360 46452 1362 46472
rect 1306 46416 1362 46452
rect 1306 45600 1362 45656
rect 1306 44784 1362 44840
rect 1306 43188 1308 43208
rect 1308 43188 1360 43208
rect 1360 43188 1362 43208
rect 1306 43152 1362 43188
rect 1306 42336 1362 42392
rect 1306 41520 1362 41576
rect 1306 40704 1362 40760
rect 3422 54576 3478 54632
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 3330 53624 3386 53680
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2042 43968 2098 44024
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2042 39924 2044 39944
rect 2044 39924 2096 39944
rect 2096 39924 2098 39944
rect 2042 39888 2098 39924
rect 3606 52944 3662 53000
rect 3514 44376 3570 44432
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 1306 39072 1362 39128
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 1306 38256 1362 38312
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 1306 37440 1362 37496
rect 1306 36660 1308 36680
rect 1308 36660 1360 36680
rect 1360 36660 1362 36680
rect 1306 36624 1362 36660
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 2778 35808 2834 35864
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 1306 34992 1362 35048
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2042 34176 2098 34232
rect 1306 33396 1308 33416
rect 1308 33396 1360 33416
rect 1360 33396 1362 33416
rect 1306 33360 1362 33396
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 1306 32544 1362 32600
rect 1306 31728 1362 31784
rect 1306 30912 1362 30968
rect 1306 30132 1308 30152
rect 1308 30132 1360 30152
rect 1360 30132 1362 30152
rect 1306 30096 1362 30132
rect 1306 29280 1362 29336
rect 1306 28464 1362 28520
rect 1306 27648 1362 27704
rect 938 26832 994 26888
rect 1674 26016 1730 26072
rect 938 25236 940 25256
rect 940 25236 992 25256
rect 992 25236 994 25256
rect 938 25200 994 25236
rect 938 24384 994 24440
rect 938 23568 994 23624
rect 938 22752 994 22808
rect 938 21956 994 21992
rect 938 21936 940 21956
rect 940 21936 992 21956
rect 992 21936 994 21956
rect 938 21120 994 21176
rect 938 20304 994 20360
rect 938 19488 994 19544
rect 938 18708 940 18728
rect 940 18708 992 18728
rect 992 18708 994 18728
rect 938 18672 994 18708
rect 1582 17856 1638 17912
rect 938 17040 994 17096
rect 938 16224 994 16280
rect 938 15428 994 15464
rect 938 15408 940 15428
rect 940 15408 992 15428
rect 992 15408 994 15428
rect 938 14592 994 14648
rect 938 13776 994 13832
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 13634 45892 13690 45928
rect 13634 45872 13636 45892
rect 13636 45872 13688 45892
rect 13688 45872 13690 45892
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 13450 44104 13506 44160
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 11978 36624 12034 36680
rect 11058 35944 11114 36000
rect 10874 35128 10930 35184
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 13634 40432 13690 40488
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 14554 38120 14610 38176
rect 14646 35708 14648 35728
rect 14648 35708 14700 35728
rect 14700 35708 14702 35728
rect 14646 35672 14702 35708
rect 14646 35128 14702 35184
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 15106 36352 15162 36408
rect 15106 36080 15162 36136
rect 14922 35672 14978 35728
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 2042 17040 2098 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 938 12960 994 13016
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 938 12164 994 12200
rect 938 12144 940 12164
rect 940 12144 992 12164
rect 992 12144 994 12164
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 938 11328 994 11384
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 938 10512 994 10568
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 938 9696 994 9752
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 1582 8064 1638 8120
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 938 7248 994 7304
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 938 6432 994 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 16118 39072 16174 39128
rect 938 5636 994 5672
rect 938 5616 940 5636
rect 940 5616 992 5636
rect 992 5616 994 5636
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 938 4800 994 4856
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 938 3984 994 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 938 3168 994 3224
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 15934 36352 15990 36408
rect 16302 37712 16358 37768
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 16762 36780 16818 36816
rect 16762 36760 16764 36780
rect 16764 36760 16816 36780
rect 16816 36760 16818 36780
rect 16026 35672 16082 35728
rect 16026 29164 16082 29200
rect 16026 29144 16028 29164
rect 16028 29144 16080 29164
rect 16080 29144 16082 29164
rect 16946 36352 17002 36408
rect 16854 36236 16910 36272
rect 16854 36216 16856 36236
rect 16856 36216 16908 36236
rect 16908 36216 16910 36236
rect 16302 29144 16358 29200
rect 17406 38156 17408 38176
rect 17408 38156 17460 38176
rect 17460 38156 17462 38176
rect 17406 38120 17462 38156
rect 17314 37168 17370 37224
rect 16946 27512 17002 27568
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 18418 39888 18474 39944
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17774 39092 17830 39128
rect 17774 39072 17776 39092
rect 17776 39072 17828 39092
rect 17828 39072 17830 39092
rect 18418 39092 18474 39128
rect 18418 39072 18420 39092
rect 18420 39072 18472 39092
rect 18472 39072 18474 39092
rect 17498 36488 17554 36544
rect 17314 35944 17370 36000
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 18970 39888 19026 39944
rect 18602 39244 18604 39264
rect 18604 39244 18656 39264
rect 18656 39244 18658 39264
rect 18602 39208 18658 39244
rect 18234 34992 18290 35048
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 18234 34176 18290 34232
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 27956 54426 28012 54428
rect 28036 54426 28092 54428
rect 28116 54426 28172 54428
rect 28196 54426 28252 54428
rect 27956 54374 28002 54426
rect 28002 54374 28012 54426
rect 28036 54374 28066 54426
rect 28066 54374 28078 54426
rect 28078 54374 28092 54426
rect 28116 54374 28130 54426
rect 28130 54374 28142 54426
rect 28142 54374 28172 54426
rect 28196 54374 28206 54426
rect 28206 54374 28252 54426
rect 27956 54372 28012 54374
rect 28036 54372 28092 54374
rect 28116 54372 28172 54374
rect 28196 54372 28252 54374
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 19154 40432 19210 40488
rect 19062 39480 19118 39536
rect 18786 37168 18842 37224
rect 18694 36216 18750 36272
rect 18878 36760 18934 36816
rect 19062 36760 19118 36816
rect 18694 34856 18750 34912
rect 19706 38528 19762 38584
rect 19430 38120 19486 38176
rect 19246 36524 19248 36544
rect 19248 36524 19300 36544
rect 19300 36524 19302 36544
rect 19246 36488 19302 36524
rect 18970 34176 19026 34232
rect 20350 41520 20406 41576
rect 20074 40588 20130 40624
rect 20074 40568 20076 40588
rect 20076 40568 20128 40588
rect 20128 40568 20130 40588
rect 19982 38392 20038 38448
rect 20074 38256 20130 38312
rect 19614 36080 19670 36136
rect 19798 35536 19854 35592
rect 20258 36896 20314 36952
rect 20442 40568 20498 40624
rect 20902 41384 20958 41440
rect 21178 41384 21234 41440
rect 20902 36624 20958 36680
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 20718 31728 20774 31784
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 21914 43152 21970 43208
rect 21730 38528 21786 38584
rect 21362 31728 21418 31784
rect 22374 44376 22430 44432
rect 22558 40588 22614 40624
rect 22558 40568 22560 40588
rect 22560 40568 22612 40588
rect 22612 40568 22614 40588
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22834 40160 22890 40216
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22742 38972 22744 38992
rect 22744 38972 22796 38992
rect 22796 38972 22798 38992
rect 22742 38936 22798 38972
rect 23018 39516 23020 39536
rect 23020 39516 23072 39536
rect 23072 39516 23074 39536
rect 23018 39480 23074 39516
rect 22926 38800 22982 38856
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 23386 38936 23442 38992
rect 22374 32952 22430 33008
rect 22650 33088 22706 33144
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 23386 37868 23442 37904
rect 23386 37848 23388 37868
rect 23388 37848 23440 37868
rect 23440 37848 23442 37868
rect 23846 44240 23902 44296
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 23202 34584 23258 34640
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22926 32952 22982 33008
rect 22098 29144 22154 29200
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 23386 35572 23388 35592
rect 23388 35572 23440 35592
rect 23440 35572 23442 35592
rect 23386 35536 23442 35572
rect 23386 35436 23388 35456
rect 23388 35436 23440 35456
rect 23440 35436 23442 35456
rect 23386 35400 23442 35436
rect 23386 34720 23442 34776
rect 23846 35944 23902 36000
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 25318 46996 25320 47016
rect 25320 46996 25372 47016
rect 25372 46996 25374 47016
rect 25318 46960 25374 46996
rect 24858 41384 24914 41440
rect 24398 39480 24454 39536
rect 24582 38800 24638 38856
rect 24398 37848 24454 37904
rect 25318 41384 25374 41440
rect 25226 41268 25282 41304
rect 25226 41248 25228 41268
rect 25228 41248 25280 41268
rect 25280 41248 25282 41268
rect 26238 46688 26294 46744
rect 24766 37868 24822 37904
rect 24766 37848 24768 37868
rect 24768 37848 24820 37868
rect 24820 37848 24822 37868
rect 24398 35944 24454 36000
rect 25226 36896 25282 36952
rect 25410 38120 25466 38176
rect 25502 35944 25558 36000
rect 25686 38256 25742 38312
rect 25870 37868 25926 37904
rect 25870 37848 25872 37868
rect 25872 37848 25924 37868
rect 25924 37848 25926 37868
rect 26238 40452 26294 40488
rect 26238 40432 26240 40452
rect 26240 40432 26292 40452
rect 26292 40432 26294 40452
rect 26882 47096 26938 47152
rect 26330 39752 26386 39808
rect 26330 38936 26386 38992
rect 26698 43152 26754 43208
rect 26606 41520 26662 41576
rect 27618 47132 27620 47152
rect 27620 47132 27672 47152
rect 27672 47132 27674 47152
rect 27618 47096 27674 47132
rect 27618 46688 27674 46744
rect 27342 46008 27398 46064
rect 26054 36080 26110 36136
rect 25686 35944 25742 36000
rect 26330 35400 26386 35456
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 26698 35128 26754 35184
rect 27956 53338 28012 53340
rect 28036 53338 28092 53340
rect 28116 53338 28172 53340
rect 28196 53338 28252 53340
rect 27956 53286 28002 53338
rect 28002 53286 28012 53338
rect 28036 53286 28066 53338
rect 28066 53286 28078 53338
rect 28078 53286 28092 53338
rect 28116 53286 28130 53338
rect 28130 53286 28142 53338
rect 28142 53286 28172 53338
rect 28196 53286 28206 53338
rect 28206 53286 28252 53338
rect 27956 53284 28012 53286
rect 28036 53284 28092 53286
rect 28116 53284 28172 53286
rect 28196 53284 28252 53286
rect 27956 52250 28012 52252
rect 28036 52250 28092 52252
rect 28116 52250 28172 52252
rect 28196 52250 28252 52252
rect 27956 52198 28002 52250
rect 28002 52198 28012 52250
rect 28036 52198 28066 52250
rect 28066 52198 28078 52250
rect 28078 52198 28092 52250
rect 28116 52198 28130 52250
rect 28130 52198 28142 52250
rect 28142 52198 28172 52250
rect 28196 52198 28206 52250
rect 28206 52198 28252 52250
rect 27956 52196 28012 52198
rect 28036 52196 28092 52198
rect 28116 52196 28172 52198
rect 28196 52196 28252 52198
rect 27956 51162 28012 51164
rect 28036 51162 28092 51164
rect 28116 51162 28172 51164
rect 28196 51162 28252 51164
rect 27956 51110 28002 51162
rect 28002 51110 28012 51162
rect 28036 51110 28066 51162
rect 28066 51110 28078 51162
rect 28078 51110 28092 51162
rect 28116 51110 28130 51162
rect 28130 51110 28142 51162
rect 28142 51110 28172 51162
rect 28196 51110 28206 51162
rect 28206 51110 28252 51162
rect 27956 51108 28012 51110
rect 28036 51108 28092 51110
rect 28116 51108 28172 51110
rect 28196 51108 28252 51110
rect 27956 50074 28012 50076
rect 28036 50074 28092 50076
rect 28116 50074 28172 50076
rect 28196 50074 28252 50076
rect 27956 50022 28002 50074
rect 28002 50022 28012 50074
rect 28036 50022 28066 50074
rect 28066 50022 28078 50074
rect 28078 50022 28092 50074
rect 28116 50022 28130 50074
rect 28130 50022 28142 50074
rect 28142 50022 28172 50074
rect 28196 50022 28206 50074
rect 28206 50022 28252 50074
rect 27956 50020 28012 50022
rect 28036 50020 28092 50022
rect 28116 50020 28172 50022
rect 28196 50020 28252 50022
rect 27956 48986 28012 48988
rect 28036 48986 28092 48988
rect 28116 48986 28172 48988
rect 28196 48986 28252 48988
rect 27956 48934 28002 48986
rect 28002 48934 28012 48986
rect 28036 48934 28066 48986
rect 28066 48934 28078 48986
rect 28078 48934 28092 48986
rect 28116 48934 28130 48986
rect 28130 48934 28142 48986
rect 28142 48934 28172 48986
rect 28196 48934 28206 48986
rect 28206 48934 28252 48986
rect 27956 48932 28012 48934
rect 28036 48932 28092 48934
rect 28116 48932 28172 48934
rect 28196 48932 28252 48934
rect 27956 47898 28012 47900
rect 28036 47898 28092 47900
rect 28116 47898 28172 47900
rect 28196 47898 28252 47900
rect 27956 47846 28002 47898
rect 28002 47846 28012 47898
rect 28036 47846 28066 47898
rect 28066 47846 28078 47898
rect 28078 47846 28092 47898
rect 28116 47846 28130 47898
rect 28130 47846 28142 47898
rect 28142 47846 28172 47898
rect 28196 47846 28206 47898
rect 28206 47846 28252 47898
rect 27956 47844 28012 47846
rect 28036 47844 28092 47846
rect 28116 47844 28172 47846
rect 28196 47844 28252 47846
rect 27956 46810 28012 46812
rect 28036 46810 28092 46812
rect 28116 46810 28172 46812
rect 28196 46810 28252 46812
rect 27956 46758 28002 46810
rect 28002 46758 28012 46810
rect 28036 46758 28066 46810
rect 28066 46758 28078 46810
rect 28078 46758 28092 46810
rect 28116 46758 28130 46810
rect 28130 46758 28142 46810
rect 28142 46758 28172 46810
rect 28196 46758 28206 46810
rect 28206 46758 28252 46810
rect 27956 46756 28012 46758
rect 28036 46756 28092 46758
rect 28116 46756 28172 46758
rect 28196 46756 28252 46758
rect 27894 45872 27950 45928
rect 27956 45722 28012 45724
rect 28036 45722 28092 45724
rect 28116 45722 28172 45724
rect 28196 45722 28252 45724
rect 27956 45670 28002 45722
rect 28002 45670 28012 45722
rect 28036 45670 28066 45722
rect 28066 45670 28078 45722
rect 28078 45670 28092 45722
rect 28116 45670 28130 45722
rect 28130 45670 28142 45722
rect 28142 45670 28172 45722
rect 28196 45670 28206 45722
rect 28206 45670 28252 45722
rect 27956 45668 28012 45670
rect 28036 45668 28092 45670
rect 28116 45668 28172 45670
rect 28196 45668 28252 45670
rect 28538 46824 28594 46880
rect 27956 44634 28012 44636
rect 28036 44634 28092 44636
rect 28116 44634 28172 44636
rect 28196 44634 28252 44636
rect 27956 44582 28002 44634
rect 28002 44582 28012 44634
rect 28036 44582 28066 44634
rect 28066 44582 28078 44634
rect 28078 44582 28092 44634
rect 28116 44582 28130 44634
rect 28130 44582 28142 44634
rect 28142 44582 28172 44634
rect 28196 44582 28206 44634
rect 28206 44582 28252 44634
rect 27956 44580 28012 44582
rect 28036 44580 28092 44582
rect 28116 44580 28172 44582
rect 28196 44580 28252 44582
rect 27342 39924 27344 39944
rect 27344 39924 27396 39944
rect 27396 39924 27398 39944
rect 27342 39888 27398 39924
rect 27434 39208 27490 39264
rect 27342 39072 27398 39128
rect 27434 38800 27490 38856
rect 27956 43546 28012 43548
rect 28036 43546 28092 43548
rect 28116 43546 28172 43548
rect 28196 43546 28252 43548
rect 27956 43494 28002 43546
rect 28002 43494 28012 43546
rect 28036 43494 28066 43546
rect 28066 43494 28078 43546
rect 28078 43494 28092 43546
rect 28116 43494 28130 43546
rect 28130 43494 28142 43546
rect 28142 43494 28172 43546
rect 28196 43494 28206 43546
rect 28206 43494 28252 43546
rect 27956 43492 28012 43494
rect 28036 43492 28092 43494
rect 28116 43492 28172 43494
rect 28196 43492 28252 43494
rect 28538 44276 28540 44296
rect 28540 44276 28592 44296
rect 28592 44276 28594 44296
rect 28538 44240 28594 44276
rect 27956 42458 28012 42460
rect 28036 42458 28092 42460
rect 28116 42458 28172 42460
rect 28196 42458 28252 42460
rect 27956 42406 28002 42458
rect 28002 42406 28012 42458
rect 28036 42406 28066 42458
rect 28066 42406 28078 42458
rect 28078 42406 28092 42458
rect 28116 42406 28130 42458
rect 28130 42406 28142 42458
rect 28142 42406 28172 42458
rect 28196 42406 28206 42458
rect 28206 42406 28252 42458
rect 27956 42404 28012 42406
rect 28036 42404 28092 42406
rect 28116 42404 28172 42406
rect 28196 42404 28252 42406
rect 27342 37712 27398 37768
rect 27956 41370 28012 41372
rect 28036 41370 28092 41372
rect 28116 41370 28172 41372
rect 28196 41370 28252 41372
rect 27956 41318 28002 41370
rect 28002 41318 28012 41370
rect 28036 41318 28066 41370
rect 28066 41318 28078 41370
rect 28078 41318 28092 41370
rect 28116 41318 28130 41370
rect 28130 41318 28142 41370
rect 28142 41318 28172 41370
rect 28196 41318 28206 41370
rect 28206 41318 28252 41370
rect 27956 41316 28012 41318
rect 28036 41316 28092 41318
rect 28116 41316 28172 41318
rect 28196 41316 28252 41318
rect 27956 40282 28012 40284
rect 28036 40282 28092 40284
rect 28116 40282 28172 40284
rect 28196 40282 28252 40284
rect 27956 40230 28002 40282
rect 28002 40230 28012 40282
rect 28036 40230 28066 40282
rect 28066 40230 28078 40282
rect 28078 40230 28092 40282
rect 28116 40230 28130 40282
rect 28130 40230 28142 40282
rect 28142 40230 28172 40282
rect 28196 40230 28206 40282
rect 28206 40230 28252 40282
rect 27956 40228 28012 40230
rect 28036 40228 28092 40230
rect 28116 40228 28172 40230
rect 28196 40228 28252 40230
rect 27956 39194 28012 39196
rect 28036 39194 28092 39196
rect 28116 39194 28172 39196
rect 28196 39194 28252 39196
rect 27956 39142 28002 39194
rect 28002 39142 28012 39194
rect 28036 39142 28066 39194
rect 28066 39142 28078 39194
rect 28078 39142 28092 39194
rect 28116 39142 28130 39194
rect 28130 39142 28142 39194
rect 28142 39142 28172 39194
rect 28196 39142 28206 39194
rect 28206 39142 28252 39194
rect 27956 39140 28012 39142
rect 28036 39140 28092 39142
rect 28116 39140 28172 39142
rect 28196 39140 28252 39142
rect 27956 38106 28012 38108
rect 28036 38106 28092 38108
rect 28116 38106 28172 38108
rect 28196 38106 28252 38108
rect 27956 38054 28002 38106
rect 28002 38054 28012 38106
rect 28036 38054 28066 38106
rect 28066 38054 28078 38106
rect 28078 38054 28092 38106
rect 28116 38054 28130 38106
rect 28130 38054 28142 38106
rect 28142 38054 28172 38106
rect 28196 38054 28206 38106
rect 28206 38054 28252 38106
rect 27956 38052 28012 38054
rect 28036 38052 28092 38054
rect 28116 38052 28172 38054
rect 28196 38052 28252 38054
rect 28262 37712 28318 37768
rect 28814 46996 28816 47016
rect 28816 46996 28868 47016
rect 28868 46996 28870 47016
rect 28814 46960 28870 46996
rect 29274 46008 29330 46064
rect 28630 40840 28686 40896
rect 28538 40704 28594 40760
rect 28538 40432 28594 40488
rect 27956 37018 28012 37020
rect 28036 37018 28092 37020
rect 28116 37018 28172 37020
rect 28196 37018 28252 37020
rect 27956 36966 28002 37018
rect 28002 36966 28012 37018
rect 28036 36966 28066 37018
rect 28066 36966 28078 37018
rect 28078 36966 28092 37018
rect 28116 36966 28130 37018
rect 28130 36966 28142 37018
rect 28142 36966 28172 37018
rect 28196 36966 28206 37018
rect 28206 36966 28252 37018
rect 27956 36964 28012 36966
rect 28036 36964 28092 36966
rect 28116 36964 28172 36966
rect 28196 36964 28252 36966
rect 27342 34584 27398 34640
rect 28170 36100 28226 36136
rect 28170 36080 28172 36100
rect 28172 36080 28224 36100
rect 28224 36080 28226 36100
rect 27956 35930 28012 35932
rect 28036 35930 28092 35932
rect 28116 35930 28172 35932
rect 28196 35930 28252 35932
rect 27956 35878 28002 35930
rect 28002 35878 28012 35930
rect 28036 35878 28066 35930
rect 28066 35878 28078 35930
rect 28078 35878 28092 35930
rect 28116 35878 28130 35930
rect 28130 35878 28142 35930
rect 28142 35878 28172 35930
rect 28196 35878 28206 35930
rect 28206 35878 28252 35930
rect 27956 35876 28012 35878
rect 28036 35876 28092 35878
rect 28116 35876 28172 35878
rect 28196 35876 28252 35878
rect 27986 35264 28042 35320
rect 27986 34992 28042 35048
rect 27956 34842 28012 34844
rect 28036 34842 28092 34844
rect 28116 34842 28172 34844
rect 28196 34842 28252 34844
rect 27956 34790 28002 34842
rect 28002 34790 28012 34842
rect 28036 34790 28066 34842
rect 28066 34790 28078 34842
rect 28078 34790 28092 34842
rect 28116 34790 28130 34842
rect 28130 34790 28142 34842
rect 28142 34790 28172 34842
rect 28196 34790 28206 34842
rect 28206 34790 28252 34842
rect 27956 34788 28012 34790
rect 28036 34788 28092 34790
rect 28116 34788 28172 34790
rect 28196 34788 28252 34790
rect 27956 33754 28012 33756
rect 28036 33754 28092 33756
rect 28116 33754 28172 33756
rect 28196 33754 28252 33756
rect 27956 33702 28002 33754
rect 28002 33702 28012 33754
rect 28036 33702 28066 33754
rect 28066 33702 28078 33754
rect 28078 33702 28092 33754
rect 28116 33702 28130 33754
rect 28130 33702 28142 33754
rect 28142 33702 28172 33754
rect 28196 33702 28206 33754
rect 28206 33702 28252 33754
rect 27956 33700 28012 33702
rect 28036 33700 28092 33702
rect 28116 33700 28172 33702
rect 28196 33700 28252 33702
rect 28630 36080 28686 36136
rect 27956 32666 28012 32668
rect 28036 32666 28092 32668
rect 28116 32666 28172 32668
rect 28196 32666 28252 32668
rect 27956 32614 28002 32666
rect 28002 32614 28012 32666
rect 28036 32614 28066 32666
rect 28066 32614 28078 32666
rect 28078 32614 28092 32666
rect 28116 32614 28130 32666
rect 28130 32614 28142 32666
rect 28142 32614 28172 32666
rect 28196 32614 28206 32666
rect 28206 32614 28252 32666
rect 27956 32612 28012 32614
rect 28036 32612 28092 32614
rect 28116 32612 28172 32614
rect 28196 32612 28252 32614
rect 27956 31578 28012 31580
rect 28036 31578 28092 31580
rect 28116 31578 28172 31580
rect 28196 31578 28252 31580
rect 27956 31526 28002 31578
rect 28002 31526 28012 31578
rect 28036 31526 28066 31578
rect 28066 31526 28078 31578
rect 28078 31526 28092 31578
rect 28116 31526 28130 31578
rect 28130 31526 28142 31578
rect 28142 31526 28172 31578
rect 28196 31526 28206 31578
rect 28206 31526 28252 31578
rect 27956 31524 28012 31526
rect 28036 31524 28092 31526
rect 28116 31524 28172 31526
rect 28196 31524 28252 31526
rect 27956 30490 28012 30492
rect 28036 30490 28092 30492
rect 28116 30490 28172 30492
rect 28196 30490 28252 30492
rect 27956 30438 28002 30490
rect 28002 30438 28012 30490
rect 28036 30438 28066 30490
rect 28066 30438 28078 30490
rect 28078 30438 28092 30490
rect 28116 30438 28130 30490
rect 28130 30438 28142 30490
rect 28142 30438 28172 30490
rect 28196 30438 28206 30490
rect 28206 30438 28252 30490
rect 27956 30436 28012 30438
rect 28036 30436 28092 30438
rect 28116 30436 28172 30438
rect 28196 30436 28252 30438
rect 27956 29402 28012 29404
rect 28036 29402 28092 29404
rect 28116 29402 28172 29404
rect 28196 29402 28252 29404
rect 27956 29350 28002 29402
rect 28002 29350 28012 29402
rect 28036 29350 28066 29402
rect 28066 29350 28078 29402
rect 28078 29350 28092 29402
rect 28116 29350 28130 29402
rect 28130 29350 28142 29402
rect 28142 29350 28172 29402
rect 28196 29350 28206 29402
rect 28206 29350 28252 29402
rect 27956 29348 28012 29350
rect 28036 29348 28092 29350
rect 28116 29348 28172 29350
rect 28196 29348 28252 29350
rect 27956 28314 28012 28316
rect 28036 28314 28092 28316
rect 28116 28314 28172 28316
rect 28196 28314 28252 28316
rect 27956 28262 28002 28314
rect 28002 28262 28012 28314
rect 28036 28262 28066 28314
rect 28066 28262 28078 28314
rect 28078 28262 28092 28314
rect 28116 28262 28130 28314
rect 28130 28262 28142 28314
rect 28142 28262 28172 28314
rect 28196 28262 28206 28314
rect 28206 28262 28252 28314
rect 27956 28260 28012 28262
rect 28036 28260 28092 28262
rect 28116 28260 28172 28262
rect 28196 28260 28252 28262
rect 28906 40840 28962 40896
rect 28998 40568 29054 40624
rect 29182 39752 29238 39808
rect 28906 39616 28962 39672
rect 28814 34584 28870 34640
rect 30102 44240 30158 44296
rect 29642 35264 29698 35320
rect 27956 27226 28012 27228
rect 28036 27226 28092 27228
rect 28116 27226 28172 27228
rect 28196 27226 28252 27228
rect 27956 27174 28002 27226
rect 28002 27174 28012 27226
rect 28036 27174 28066 27226
rect 28066 27174 28078 27226
rect 28078 27174 28092 27226
rect 28116 27174 28130 27226
rect 28130 27174 28142 27226
rect 28142 27174 28172 27226
rect 28196 27174 28206 27226
rect 28206 27174 28252 27226
rect 27956 27172 28012 27174
rect 28036 27172 28092 27174
rect 28116 27172 28172 27174
rect 28196 27172 28252 27174
rect 27956 26138 28012 26140
rect 28036 26138 28092 26140
rect 28116 26138 28172 26140
rect 28196 26138 28252 26140
rect 27956 26086 28002 26138
rect 28002 26086 28012 26138
rect 28036 26086 28066 26138
rect 28066 26086 28078 26138
rect 28078 26086 28092 26138
rect 28116 26086 28130 26138
rect 28130 26086 28142 26138
rect 28142 26086 28172 26138
rect 28196 26086 28206 26138
rect 28206 26086 28252 26138
rect 27956 26084 28012 26086
rect 28036 26084 28092 26086
rect 28116 26084 28172 26086
rect 28196 26084 28252 26086
rect 27956 25050 28012 25052
rect 28036 25050 28092 25052
rect 28116 25050 28172 25052
rect 28196 25050 28252 25052
rect 27956 24998 28002 25050
rect 28002 24998 28012 25050
rect 28036 24998 28066 25050
rect 28066 24998 28078 25050
rect 28078 24998 28092 25050
rect 28116 24998 28130 25050
rect 28130 24998 28142 25050
rect 28142 24998 28172 25050
rect 28196 24998 28206 25050
rect 28206 24998 28252 25050
rect 27956 24996 28012 24998
rect 28036 24996 28092 24998
rect 28116 24996 28172 24998
rect 28196 24996 28252 24998
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 28906 31884 28962 31920
rect 28906 31864 28908 31884
rect 28908 31864 28960 31884
rect 28960 31864 28962 31884
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 30378 38256 30434 38312
rect 30010 33516 30066 33552
rect 30010 33496 30012 33516
rect 30012 33496 30064 33516
rect 30064 33496 30066 33516
rect 30286 32836 30342 32872
rect 30286 32816 30288 32836
rect 30288 32816 30340 32836
rect 30340 32816 30342 32836
rect 31206 42336 31262 42392
rect 31206 40976 31262 41032
rect 31574 43288 31630 43344
rect 31206 38936 31262 38992
rect 30930 37324 30986 37360
rect 30930 37304 30932 37324
rect 30932 37304 30984 37324
rect 30984 37304 30986 37324
rect 31206 37168 31262 37224
rect 31298 32816 31354 32872
rect 32126 48184 32182 48240
rect 32956 53882 33012 53884
rect 33036 53882 33092 53884
rect 33116 53882 33172 53884
rect 33196 53882 33252 53884
rect 32956 53830 33002 53882
rect 33002 53830 33012 53882
rect 33036 53830 33066 53882
rect 33066 53830 33078 53882
rect 33078 53830 33092 53882
rect 33116 53830 33130 53882
rect 33130 53830 33142 53882
rect 33142 53830 33172 53882
rect 33196 53830 33206 53882
rect 33206 53830 33252 53882
rect 32956 53828 33012 53830
rect 33036 53828 33092 53830
rect 33116 53828 33172 53830
rect 33196 53828 33252 53830
rect 32956 52794 33012 52796
rect 33036 52794 33092 52796
rect 33116 52794 33172 52796
rect 33196 52794 33252 52796
rect 32956 52742 33002 52794
rect 33002 52742 33012 52794
rect 33036 52742 33066 52794
rect 33066 52742 33078 52794
rect 33078 52742 33092 52794
rect 33116 52742 33130 52794
rect 33130 52742 33142 52794
rect 33142 52742 33172 52794
rect 33196 52742 33206 52794
rect 33206 52742 33252 52794
rect 32956 52740 33012 52742
rect 33036 52740 33092 52742
rect 33116 52740 33172 52742
rect 33196 52740 33252 52742
rect 32956 51706 33012 51708
rect 33036 51706 33092 51708
rect 33116 51706 33172 51708
rect 33196 51706 33252 51708
rect 32956 51654 33002 51706
rect 33002 51654 33012 51706
rect 33036 51654 33066 51706
rect 33066 51654 33078 51706
rect 33078 51654 33092 51706
rect 33116 51654 33130 51706
rect 33130 51654 33142 51706
rect 33142 51654 33172 51706
rect 33196 51654 33206 51706
rect 33206 51654 33252 51706
rect 32956 51652 33012 51654
rect 33036 51652 33092 51654
rect 33116 51652 33172 51654
rect 33196 51652 33252 51654
rect 32956 50618 33012 50620
rect 33036 50618 33092 50620
rect 33116 50618 33172 50620
rect 33196 50618 33252 50620
rect 32956 50566 33002 50618
rect 33002 50566 33012 50618
rect 33036 50566 33066 50618
rect 33066 50566 33078 50618
rect 33078 50566 33092 50618
rect 33116 50566 33130 50618
rect 33130 50566 33142 50618
rect 33142 50566 33172 50618
rect 33196 50566 33206 50618
rect 33206 50566 33252 50618
rect 32956 50564 33012 50566
rect 33036 50564 33092 50566
rect 33116 50564 33172 50566
rect 33196 50564 33252 50566
rect 32770 48048 32826 48104
rect 32956 49530 33012 49532
rect 33036 49530 33092 49532
rect 33116 49530 33172 49532
rect 33196 49530 33252 49532
rect 32956 49478 33002 49530
rect 33002 49478 33012 49530
rect 33036 49478 33066 49530
rect 33066 49478 33078 49530
rect 33078 49478 33092 49530
rect 33116 49478 33130 49530
rect 33130 49478 33142 49530
rect 33142 49478 33172 49530
rect 33196 49478 33206 49530
rect 33206 49478 33252 49530
rect 32956 49476 33012 49478
rect 33036 49476 33092 49478
rect 33116 49476 33172 49478
rect 33196 49476 33252 49478
rect 32956 48442 33012 48444
rect 33036 48442 33092 48444
rect 33116 48442 33172 48444
rect 33196 48442 33252 48444
rect 32956 48390 33002 48442
rect 33002 48390 33012 48442
rect 33036 48390 33066 48442
rect 33066 48390 33078 48442
rect 33078 48390 33092 48442
rect 33116 48390 33130 48442
rect 33130 48390 33142 48442
rect 33142 48390 33172 48442
rect 33196 48390 33206 48442
rect 33206 48390 33252 48442
rect 32956 48388 33012 48390
rect 33036 48388 33092 48390
rect 33116 48388 33172 48390
rect 33196 48388 33252 48390
rect 32956 47354 33012 47356
rect 33036 47354 33092 47356
rect 33116 47354 33172 47356
rect 33196 47354 33252 47356
rect 32956 47302 33002 47354
rect 33002 47302 33012 47354
rect 33036 47302 33066 47354
rect 33066 47302 33078 47354
rect 33078 47302 33092 47354
rect 33116 47302 33130 47354
rect 33130 47302 33142 47354
rect 33142 47302 33172 47354
rect 33196 47302 33206 47354
rect 33206 47302 33252 47354
rect 32956 47300 33012 47302
rect 33036 47300 33092 47302
rect 33116 47300 33172 47302
rect 33196 47300 33252 47302
rect 32956 46266 33012 46268
rect 33036 46266 33092 46268
rect 33116 46266 33172 46268
rect 33196 46266 33252 46268
rect 32956 46214 33002 46266
rect 33002 46214 33012 46266
rect 33036 46214 33066 46266
rect 33066 46214 33078 46266
rect 33078 46214 33092 46266
rect 33116 46214 33130 46266
rect 33130 46214 33142 46266
rect 33142 46214 33172 46266
rect 33196 46214 33206 46266
rect 33206 46214 33252 46266
rect 32956 46212 33012 46214
rect 33036 46212 33092 46214
rect 33116 46212 33172 46214
rect 33196 46212 33252 46214
rect 31758 39636 31814 39672
rect 31758 39616 31760 39636
rect 31760 39616 31812 39636
rect 31812 39616 31814 39636
rect 31942 39072 31998 39128
rect 31758 37032 31814 37088
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 30378 14320 30434 14376
rect 32126 41248 32182 41304
rect 32956 45178 33012 45180
rect 33036 45178 33092 45180
rect 33116 45178 33172 45180
rect 33196 45178 33252 45180
rect 32956 45126 33002 45178
rect 33002 45126 33012 45178
rect 33036 45126 33066 45178
rect 33066 45126 33078 45178
rect 33078 45126 33092 45178
rect 33116 45126 33130 45178
rect 33130 45126 33142 45178
rect 33142 45126 33172 45178
rect 33196 45126 33206 45178
rect 33206 45126 33252 45178
rect 32956 45124 33012 45126
rect 33036 45124 33092 45126
rect 33116 45124 33172 45126
rect 33196 45124 33252 45126
rect 33138 44940 33194 44976
rect 33138 44920 33140 44940
rect 33140 44920 33192 44940
rect 33192 44920 33194 44940
rect 32956 44090 33012 44092
rect 33036 44090 33092 44092
rect 33116 44090 33172 44092
rect 33196 44090 33252 44092
rect 32956 44038 33002 44090
rect 33002 44038 33012 44090
rect 33036 44038 33066 44090
rect 33066 44038 33078 44090
rect 33078 44038 33092 44090
rect 33116 44038 33130 44090
rect 33130 44038 33142 44090
rect 33142 44038 33172 44090
rect 33196 44038 33206 44090
rect 33206 44038 33252 44090
rect 32956 44036 33012 44038
rect 33036 44036 33092 44038
rect 33116 44036 33172 44038
rect 33196 44036 33252 44038
rect 32956 43002 33012 43004
rect 33036 43002 33092 43004
rect 33116 43002 33172 43004
rect 33196 43002 33252 43004
rect 32956 42950 33002 43002
rect 33002 42950 33012 43002
rect 33036 42950 33066 43002
rect 33066 42950 33078 43002
rect 33078 42950 33092 43002
rect 33116 42950 33130 43002
rect 33130 42950 33142 43002
rect 33142 42950 33172 43002
rect 33196 42950 33206 43002
rect 33206 42950 33252 43002
rect 32956 42948 33012 42950
rect 33036 42948 33092 42950
rect 33116 42948 33172 42950
rect 33196 42948 33252 42950
rect 32494 41248 32550 41304
rect 32494 40976 32550 41032
rect 32218 39072 32274 39128
rect 32494 39752 32550 39808
rect 32956 41914 33012 41916
rect 33036 41914 33092 41916
rect 33116 41914 33172 41916
rect 33196 41914 33252 41916
rect 32956 41862 33002 41914
rect 33002 41862 33012 41914
rect 33036 41862 33066 41914
rect 33066 41862 33078 41914
rect 33078 41862 33092 41914
rect 33116 41862 33130 41914
rect 33130 41862 33142 41914
rect 33142 41862 33172 41914
rect 33196 41862 33206 41914
rect 33206 41862 33252 41914
rect 32956 41860 33012 41862
rect 33036 41860 33092 41862
rect 33116 41860 33172 41862
rect 33196 41860 33252 41862
rect 37956 54426 38012 54428
rect 38036 54426 38092 54428
rect 38116 54426 38172 54428
rect 38196 54426 38252 54428
rect 37956 54374 38002 54426
rect 38002 54374 38012 54426
rect 38036 54374 38066 54426
rect 38066 54374 38078 54426
rect 38078 54374 38092 54426
rect 38116 54374 38130 54426
rect 38130 54374 38142 54426
rect 38142 54374 38172 54426
rect 38196 54374 38206 54426
rect 38206 54374 38252 54426
rect 37956 54372 38012 54374
rect 38036 54372 38092 54374
rect 38116 54372 38172 54374
rect 38196 54372 38252 54374
rect 33782 48184 33838 48240
rect 33506 44104 33562 44160
rect 32956 40826 33012 40828
rect 33036 40826 33092 40828
rect 33116 40826 33172 40828
rect 33196 40826 33252 40828
rect 32956 40774 33002 40826
rect 33002 40774 33012 40826
rect 33036 40774 33066 40826
rect 33066 40774 33078 40826
rect 33078 40774 33092 40826
rect 33116 40774 33130 40826
rect 33130 40774 33142 40826
rect 33142 40774 33172 40826
rect 33196 40774 33206 40826
rect 33206 40774 33252 40826
rect 32956 40772 33012 40774
rect 33036 40772 33092 40774
rect 33116 40772 33172 40774
rect 33196 40772 33252 40774
rect 33414 40024 33470 40080
rect 32770 39616 32826 39672
rect 32402 34060 32458 34096
rect 32402 34040 32404 34060
rect 32404 34040 32456 34060
rect 32456 34040 32458 34060
rect 32956 39738 33012 39740
rect 33036 39738 33092 39740
rect 33116 39738 33172 39740
rect 33196 39738 33252 39740
rect 32956 39686 33002 39738
rect 33002 39686 33012 39738
rect 33036 39686 33066 39738
rect 33066 39686 33078 39738
rect 33078 39686 33092 39738
rect 33116 39686 33130 39738
rect 33130 39686 33142 39738
rect 33142 39686 33172 39738
rect 33196 39686 33206 39738
rect 33206 39686 33252 39738
rect 32956 39684 33012 39686
rect 33036 39684 33092 39686
rect 33116 39684 33172 39686
rect 33196 39684 33252 39686
rect 32956 38650 33012 38652
rect 33036 38650 33092 38652
rect 33116 38650 33172 38652
rect 33196 38650 33252 38652
rect 32956 38598 33002 38650
rect 33002 38598 33012 38650
rect 33036 38598 33066 38650
rect 33066 38598 33078 38650
rect 33078 38598 33092 38650
rect 33116 38598 33130 38650
rect 33130 38598 33142 38650
rect 33142 38598 33172 38650
rect 33196 38598 33206 38650
rect 33206 38598 33252 38650
rect 32956 38596 33012 38598
rect 33036 38596 33092 38598
rect 33116 38596 33172 38598
rect 33196 38596 33252 38598
rect 32956 37562 33012 37564
rect 33036 37562 33092 37564
rect 33116 37562 33172 37564
rect 33196 37562 33252 37564
rect 32956 37510 33002 37562
rect 33002 37510 33012 37562
rect 33036 37510 33066 37562
rect 33066 37510 33078 37562
rect 33078 37510 33092 37562
rect 33116 37510 33130 37562
rect 33130 37510 33142 37562
rect 33142 37510 33172 37562
rect 33196 37510 33206 37562
rect 33206 37510 33252 37562
rect 32956 37508 33012 37510
rect 33036 37508 33092 37510
rect 33116 37508 33172 37510
rect 33196 37508 33252 37510
rect 32956 36474 33012 36476
rect 33036 36474 33092 36476
rect 33116 36474 33172 36476
rect 33196 36474 33252 36476
rect 32956 36422 33002 36474
rect 33002 36422 33012 36474
rect 33036 36422 33066 36474
rect 33066 36422 33078 36474
rect 33078 36422 33092 36474
rect 33116 36422 33130 36474
rect 33130 36422 33142 36474
rect 33142 36422 33172 36474
rect 33196 36422 33206 36474
rect 33206 36422 33252 36474
rect 32956 36420 33012 36422
rect 33036 36420 33092 36422
rect 33116 36420 33172 36422
rect 33196 36420 33252 36422
rect 32956 35386 33012 35388
rect 33036 35386 33092 35388
rect 33116 35386 33172 35388
rect 33196 35386 33252 35388
rect 32956 35334 33002 35386
rect 33002 35334 33012 35386
rect 33036 35334 33066 35386
rect 33066 35334 33078 35386
rect 33078 35334 33092 35386
rect 33116 35334 33130 35386
rect 33130 35334 33142 35386
rect 33142 35334 33172 35386
rect 33196 35334 33206 35386
rect 33206 35334 33252 35386
rect 32956 35332 33012 35334
rect 33036 35332 33092 35334
rect 33116 35332 33172 35334
rect 33196 35332 33252 35334
rect 32494 33496 32550 33552
rect 32956 34298 33012 34300
rect 33036 34298 33092 34300
rect 33116 34298 33172 34300
rect 33196 34298 33252 34300
rect 32956 34246 33002 34298
rect 33002 34246 33012 34298
rect 33036 34246 33066 34298
rect 33066 34246 33078 34298
rect 33078 34246 33092 34298
rect 33116 34246 33130 34298
rect 33130 34246 33142 34298
rect 33142 34246 33172 34298
rect 33196 34246 33206 34298
rect 33206 34246 33252 34298
rect 32956 34244 33012 34246
rect 33036 34244 33092 34246
rect 33116 34244 33172 34246
rect 33196 34244 33252 34246
rect 32956 33210 33012 33212
rect 33036 33210 33092 33212
rect 33116 33210 33172 33212
rect 33196 33210 33252 33212
rect 32956 33158 33002 33210
rect 33002 33158 33012 33210
rect 33036 33158 33066 33210
rect 33066 33158 33078 33210
rect 33078 33158 33092 33210
rect 33116 33158 33130 33210
rect 33130 33158 33142 33210
rect 33142 33158 33172 33210
rect 33196 33158 33206 33210
rect 33206 33158 33252 33210
rect 32956 33156 33012 33158
rect 33036 33156 33092 33158
rect 33116 33156 33172 33158
rect 33196 33156 33252 33158
rect 32956 32122 33012 32124
rect 33036 32122 33092 32124
rect 33116 32122 33172 32124
rect 33196 32122 33252 32124
rect 32956 32070 33002 32122
rect 33002 32070 33012 32122
rect 33036 32070 33066 32122
rect 33066 32070 33078 32122
rect 33078 32070 33092 32122
rect 33116 32070 33130 32122
rect 33130 32070 33142 32122
rect 33142 32070 33172 32122
rect 33196 32070 33206 32122
rect 33206 32070 33252 32122
rect 32956 32068 33012 32070
rect 33036 32068 33092 32070
rect 33116 32068 33172 32070
rect 33196 32068 33252 32070
rect 32956 31034 33012 31036
rect 33036 31034 33092 31036
rect 33116 31034 33172 31036
rect 33196 31034 33252 31036
rect 32956 30982 33002 31034
rect 33002 30982 33012 31034
rect 33036 30982 33066 31034
rect 33066 30982 33078 31034
rect 33078 30982 33092 31034
rect 33116 30982 33130 31034
rect 33130 30982 33142 31034
rect 33142 30982 33172 31034
rect 33196 30982 33206 31034
rect 33206 30982 33252 31034
rect 32956 30980 33012 30982
rect 33036 30980 33092 30982
rect 33116 30980 33172 30982
rect 33196 30980 33252 30982
rect 32956 29946 33012 29948
rect 33036 29946 33092 29948
rect 33116 29946 33172 29948
rect 33196 29946 33252 29948
rect 32956 29894 33002 29946
rect 33002 29894 33012 29946
rect 33036 29894 33066 29946
rect 33066 29894 33078 29946
rect 33078 29894 33092 29946
rect 33116 29894 33130 29946
rect 33130 29894 33142 29946
rect 33142 29894 33172 29946
rect 33196 29894 33206 29946
rect 33206 29894 33252 29946
rect 32956 29892 33012 29894
rect 33036 29892 33092 29894
rect 33116 29892 33172 29894
rect 33196 29892 33252 29894
rect 32956 28858 33012 28860
rect 33036 28858 33092 28860
rect 33116 28858 33172 28860
rect 33196 28858 33252 28860
rect 32956 28806 33002 28858
rect 33002 28806 33012 28858
rect 33036 28806 33066 28858
rect 33066 28806 33078 28858
rect 33078 28806 33092 28858
rect 33116 28806 33130 28858
rect 33130 28806 33142 28858
rect 33142 28806 33172 28858
rect 33196 28806 33206 28858
rect 33206 28806 33252 28858
rect 32956 28804 33012 28806
rect 33036 28804 33092 28806
rect 33116 28804 33172 28806
rect 33196 28804 33252 28806
rect 32956 27770 33012 27772
rect 33036 27770 33092 27772
rect 33116 27770 33172 27772
rect 33196 27770 33252 27772
rect 32956 27718 33002 27770
rect 33002 27718 33012 27770
rect 33036 27718 33066 27770
rect 33066 27718 33078 27770
rect 33078 27718 33092 27770
rect 33116 27718 33130 27770
rect 33130 27718 33142 27770
rect 33142 27718 33172 27770
rect 33196 27718 33206 27770
rect 33206 27718 33252 27770
rect 32956 27716 33012 27718
rect 33036 27716 33092 27718
rect 33116 27716 33172 27718
rect 33196 27716 33252 27718
rect 32956 26682 33012 26684
rect 33036 26682 33092 26684
rect 33116 26682 33172 26684
rect 33196 26682 33252 26684
rect 32956 26630 33002 26682
rect 33002 26630 33012 26682
rect 33036 26630 33066 26682
rect 33066 26630 33078 26682
rect 33078 26630 33092 26682
rect 33116 26630 33130 26682
rect 33130 26630 33142 26682
rect 33142 26630 33172 26682
rect 33196 26630 33206 26682
rect 33206 26630 33252 26682
rect 32956 26628 33012 26630
rect 33036 26628 33092 26630
rect 33116 26628 33172 26630
rect 33196 26628 33252 26630
rect 32956 25594 33012 25596
rect 33036 25594 33092 25596
rect 33116 25594 33172 25596
rect 33196 25594 33252 25596
rect 32956 25542 33002 25594
rect 33002 25542 33012 25594
rect 33036 25542 33066 25594
rect 33066 25542 33078 25594
rect 33078 25542 33092 25594
rect 33116 25542 33130 25594
rect 33130 25542 33142 25594
rect 33142 25542 33172 25594
rect 33196 25542 33206 25594
rect 33206 25542 33252 25594
rect 32956 25540 33012 25542
rect 33036 25540 33092 25542
rect 33116 25540 33172 25542
rect 33196 25540 33252 25542
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 34518 48184 34574 48240
rect 33874 40060 33876 40080
rect 33876 40060 33928 40080
rect 33928 40060 33930 40080
rect 33874 40024 33930 40060
rect 33966 39244 33968 39264
rect 33968 39244 34020 39264
rect 34020 39244 34022 39264
rect 33966 39208 34022 39244
rect 34794 46824 34850 46880
rect 34886 43852 34942 43888
rect 34886 43832 34888 43852
rect 34888 43832 34940 43852
rect 34940 43832 34942 43852
rect 36358 48068 36414 48104
rect 36358 48048 36360 48068
rect 36360 48048 36412 48068
rect 36412 48048 36414 48068
rect 35162 44104 35218 44160
rect 34242 37304 34298 37360
rect 34150 34040 34206 34096
rect 33414 24792 33470 24848
rect 34518 31864 34574 31920
rect 36726 48068 36782 48104
rect 36726 48048 36728 48068
rect 36728 48048 36780 48068
rect 36780 48048 36782 48068
rect 36450 44920 36506 44976
rect 36266 42336 36322 42392
rect 35990 37304 36046 37360
rect 37094 48048 37150 48104
rect 37278 48184 37334 48240
rect 37956 53338 38012 53340
rect 38036 53338 38092 53340
rect 38116 53338 38172 53340
rect 38196 53338 38252 53340
rect 37956 53286 38002 53338
rect 38002 53286 38012 53338
rect 38036 53286 38066 53338
rect 38066 53286 38078 53338
rect 38078 53286 38092 53338
rect 38116 53286 38130 53338
rect 38130 53286 38142 53338
rect 38142 53286 38172 53338
rect 38196 53286 38206 53338
rect 38206 53286 38252 53338
rect 37956 53284 38012 53286
rect 38036 53284 38092 53286
rect 38116 53284 38172 53286
rect 38196 53284 38252 53286
rect 37956 52250 38012 52252
rect 38036 52250 38092 52252
rect 38116 52250 38172 52252
rect 38196 52250 38252 52252
rect 37956 52198 38002 52250
rect 38002 52198 38012 52250
rect 38036 52198 38066 52250
rect 38066 52198 38078 52250
rect 38078 52198 38092 52250
rect 38116 52198 38130 52250
rect 38130 52198 38142 52250
rect 38142 52198 38172 52250
rect 38196 52198 38206 52250
rect 38206 52198 38252 52250
rect 37956 52196 38012 52198
rect 38036 52196 38092 52198
rect 38116 52196 38172 52198
rect 38196 52196 38252 52198
rect 37956 51162 38012 51164
rect 38036 51162 38092 51164
rect 38116 51162 38172 51164
rect 38196 51162 38252 51164
rect 37956 51110 38002 51162
rect 38002 51110 38012 51162
rect 38036 51110 38066 51162
rect 38066 51110 38078 51162
rect 38078 51110 38092 51162
rect 38116 51110 38130 51162
rect 38130 51110 38142 51162
rect 38142 51110 38172 51162
rect 38196 51110 38206 51162
rect 38206 51110 38252 51162
rect 37956 51108 38012 51110
rect 38036 51108 38092 51110
rect 38116 51108 38172 51110
rect 38196 51108 38252 51110
rect 37956 50074 38012 50076
rect 38036 50074 38092 50076
rect 38116 50074 38172 50076
rect 38196 50074 38252 50076
rect 37956 50022 38002 50074
rect 38002 50022 38012 50074
rect 38036 50022 38066 50074
rect 38066 50022 38078 50074
rect 38078 50022 38092 50074
rect 38116 50022 38130 50074
rect 38130 50022 38142 50074
rect 38142 50022 38172 50074
rect 38196 50022 38206 50074
rect 38206 50022 38252 50074
rect 37956 50020 38012 50022
rect 38036 50020 38092 50022
rect 38116 50020 38172 50022
rect 38196 50020 38252 50022
rect 37956 48986 38012 48988
rect 38036 48986 38092 48988
rect 38116 48986 38172 48988
rect 38196 48986 38252 48988
rect 37956 48934 38002 48986
rect 38002 48934 38012 48986
rect 38036 48934 38066 48986
rect 38066 48934 38078 48986
rect 38078 48934 38092 48986
rect 38116 48934 38130 48986
rect 38130 48934 38142 48986
rect 38142 48934 38172 48986
rect 38196 48934 38206 48986
rect 38206 48934 38252 48986
rect 37956 48932 38012 48934
rect 38036 48932 38092 48934
rect 38116 48932 38172 48934
rect 38196 48932 38252 48934
rect 37956 47898 38012 47900
rect 38036 47898 38092 47900
rect 38116 47898 38172 47900
rect 38196 47898 38252 47900
rect 37956 47846 38002 47898
rect 38002 47846 38012 47898
rect 38036 47846 38066 47898
rect 38066 47846 38078 47898
rect 38078 47846 38092 47898
rect 38116 47846 38130 47898
rect 38130 47846 38142 47898
rect 38142 47846 38172 47898
rect 38196 47846 38206 47898
rect 38206 47846 38252 47898
rect 37956 47844 38012 47846
rect 38036 47844 38092 47846
rect 38116 47844 38172 47846
rect 38196 47844 38252 47846
rect 37278 43852 37334 43888
rect 37278 43832 37280 43852
rect 37280 43832 37332 43852
rect 37332 43832 37334 43852
rect 36542 37848 36598 37904
rect 37956 46810 38012 46812
rect 38036 46810 38092 46812
rect 38116 46810 38172 46812
rect 38196 46810 38252 46812
rect 37956 46758 38002 46810
rect 38002 46758 38012 46810
rect 38036 46758 38066 46810
rect 38066 46758 38078 46810
rect 38078 46758 38092 46810
rect 38116 46758 38130 46810
rect 38130 46758 38142 46810
rect 38142 46758 38172 46810
rect 38196 46758 38206 46810
rect 38206 46758 38252 46810
rect 37956 46756 38012 46758
rect 38036 46756 38092 46758
rect 38116 46756 38172 46758
rect 38196 46756 38252 46758
rect 37956 45722 38012 45724
rect 38036 45722 38092 45724
rect 38116 45722 38172 45724
rect 38196 45722 38252 45724
rect 37956 45670 38002 45722
rect 38002 45670 38012 45722
rect 38036 45670 38066 45722
rect 38066 45670 38078 45722
rect 38078 45670 38092 45722
rect 38116 45670 38130 45722
rect 38130 45670 38142 45722
rect 38142 45670 38172 45722
rect 38196 45670 38206 45722
rect 38206 45670 38252 45722
rect 37956 45668 38012 45670
rect 38036 45668 38092 45670
rect 38116 45668 38172 45670
rect 38196 45668 38252 45670
rect 37554 43288 37610 43344
rect 37956 44634 38012 44636
rect 38036 44634 38092 44636
rect 38116 44634 38172 44636
rect 38196 44634 38252 44636
rect 37956 44582 38002 44634
rect 38002 44582 38012 44634
rect 38036 44582 38066 44634
rect 38066 44582 38078 44634
rect 38078 44582 38092 44634
rect 38116 44582 38130 44634
rect 38130 44582 38142 44634
rect 38142 44582 38172 44634
rect 38196 44582 38206 44634
rect 38206 44582 38252 44634
rect 37956 44580 38012 44582
rect 38036 44580 38092 44582
rect 38116 44580 38172 44582
rect 38196 44580 38252 44582
rect 42956 53882 43012 53884
rect 43036 53882 43092 53884
rect 43116 53882 43172 53884
rect 43196 53882 43252 53884
rect 42956 53830 43002 53882
rect 43002 53830 43012 53882
rect 43036 53830 43066 53882
rect 43066 53830 43078 53882
rect 43078 53830 43092 53882
rect 43116 53830 43130 53882
rect 43130 53830 43142 53882
rect 43142 53830 43172 53882
rect 43196 53830 43206 53882
rect 43206 53830 43252 53882
rect 42956 53828 43012 53830
rect 43036 53828 43092 53830
rect 43116 53828 43172 53830
rect 43196 53828 43252 53830
rect 42956 52794 43012 52796
rect 43036 52794 43092 52796
rect 43116 52794 43172 52796
rect 43196 52794 43252 52796
rect 42956 52742 43002 52794
rect 43002 52742 43012 52794
rect 43036 52742 43066 52794
rect 43066 52742 43078 52794
rect 43078 52742 43092 52794
rect 43116 52742 43130 52794
rect 43130 52742 43142 52794
rect 43142 52742 43172 52794
rect 43196 52742 43206 52794
rect 43206 52742 43252 52794
rect 42956 52740 43012 52742
rect 43036 52740 43092 52742
rect 43116 52740 43172 52742
rect 43196 52740 43252 52742
rect 42956 51706 43012 51708
rect 43036 51706 43092 51708
rect 43116 51706 43172 51708
rect 43196 51706 43252 51708
rect 42956 51654 43002 51706
rect 43002 51654 43012 51706
rect 43036 51654 43066 51706
rect 43066 51654 43078 51706
rect 43078 51654 43092 51706
rect 43116 51654 43130 51706
rect 43130 51654 43142 51706
rect 43142 51654 43172 51706
rect 43196 51654 43206 51706
rect 43206 51654 43252 51706
rect 42956 51652 43012 51654
rect 43036 51652 43092 51654
rect 43116 51652 43172 51654
rect 43196 51652 43252 51654
rect 47766 54576 47822 54632
rect 47956 54426 48012 54428
rect 48036 54426 48092 54428
rect 48116 54426 48172 54428
rect 48196 54426 48252 54428
rect 47956 54374 48002 54426
rect 48002 54374 48012 54426
rect 48036 54374 48066 54426
rect 48066 54374 48078 54426
rect 48078 54374 48092 54426
rect 48116 54374 48130 54426
rect 48130 54374 48142 54426
rect 48142 54374 48172 54426
rect 48196 54374 48206 54426
rect 48206 54374 48252 54426
rect 47956 54372 48012 54374
rect 48036 54372 48092 54374
rect 48116 54372 48172 54374
rect 48196 54372 48252 54374
rect 48318 53760 48374 53816
rect 47956 53338 48012 53340
rect 48036 53338 48092 53340
rect 48116 53338 48172 53340
rect 48196 53338 48252 53340
rect 47956 53286 48002 53338
rect 48002 53286 48012 53338
rect 48036 53286 48066 53338
rect 48066 53286 48078 53338
rect 48078 53286 48092 53338
rect 48116 53286 48130 53338
rect 48130 53286 48142 53338
rect 48142 53286 48172 53338
rect 48196 53286 48206 53338
rect 48206 53286 48252 53338
rect 47956 53284 48012 53286
rect 48036 53284 48092 53286
rect 48116 53284 48172 53286
rect 48196 53284 48252 53286
rect 48502 52980 48504 53000
rect 48504 52980 48556 53000
rect 48556 52980 48558 53000
rect 48502 52944 48558 52980
rect 42956 50618 43012 50620
rect 43036 50618 43092 50620
rect 43116 50618 43172 50620
rect 43196 50618 43252 50620
rect 42956 50566 43002 50618
rect 43002 50566 43012 50618
rect 43036 50566 43066 50618
rect 43066 50566 43078 50618
rect 43078 50566 43092 50618
rect 43116 50566 43130 50618
rect 43130 50566 43142 50618
rect 43142 50566 43172 50618
rect 43196 50566 43206 50618
rect 43206 50566 43252 50618
rect 42956 50564 43012 50566
rect 43036 50564 43092 50566
rect 43116 50564 43172 50566
rect 43196 50564 43252 50566
rect 42956 49530 43012 49532
rect 43036 49530 43092 49532
rect 43116 49530 43172 49532
rect 43196 49530 43252 49532
rect 42956 49478 43002 49530
rect 43002 49478 43012 49530
rect 43036 49478 43066 49530
rect 43066 49478 43078 49530
rect 43078 49478 43092 49530
rect 43116 49478 43130 49530
rect 43130 49478 43142 49530
rect 43142 49478 43172 49530
rect 43196 49478 43206 49530
rect 43206 49478 43252 49530
rect 42956 49476 43012 49478
rect 43036 49476 43092 49478
rect 43116 49476 43172 49478
rect 43196 49476 43252 49478
rect 42956 48442 43012 48444
rect 43036 48442 43092 48444
rect 43116 48442 43172 48444
rect 43196 48442 43252 48444
rect 42956 48390 43002 48442
rect 43002 48390 43012 48442
rect 43036 48390 43066 48442
rect 43066 48390 43078 48442
rect 43078 48390 43092 48442
rect 43116 48390 43130 48442
rect 43130 48390 43142 48442
rect 43142 48390 43172 48442
rect 43196 48390 43206 48442
rect 43206 48390 43252 48442
rect 42956 48388 43012 48390
rect 43036 48388 43092 48390
rect 43116 48388 43172 48390
rect 43196 48388 43252 48390
rect 38014 44104 38070 44160
rect 37956 43546 38012 43548
rect 38036 43546 38092 43548
rect 38116 43546 38172 43548
rect 38196 43546 38252 43548
rect 37956 43494 38002 43546
rect 38002 43494 38012 43546
rect 38036 43494 38066 43546
rect 38066 43494 38078 43546
rect 38078 43494 38092 43546
rect 38116 43494 38130 43546
rect 38130 43494 38142 43546
rect 38142 43494 38172 43546
rect 38196 43494 38206 43546
rect 38206 43494 38252 43546
rect 37956 43492 38012 43494
rect 38036 43492 38092 43494
rect 38116 43492 38172 43494
rect 38196 43492 38252 43494
rect 37646 40588 37702 40624
rect 37646 40568 37648 40588
rect 37648 40568 37700 40588
rect 37700 40568 37702 40588
rect 37646 39480 37702 39536
rect 37462 39364 37518 39400
rect 37462 39344 37464 39364
rect 37464 39344 37516 39364
rect 37516 39344 37518 39364
rect 37956 42458 38012 42460
rect 38036 42458 38092 42460
rect 38116 42458 38172 42460
rect 38196 42458 38252 42460
rect 37956 42406 38002 42458
rect 38002 42406 38012 42458
rect 38036 42406 38066 42458
rect 38066 42406 38078 42458
rect 38078 42406 38092 42458
rect 38116 42406 38130 42458
rect 38130 42406 38142 42458
rect 38142 42406 38172 42458
rect 38196 42406 38206 42458
rect 38206 42406 38252 42458
rect 37956 42404 38012 42406
rect 38036 42404 38092 42406
rect 38116 42404 38172 42406
rect 38196 42404 38252 42406
rect 37956 41370 38012 41372
rect 38036 41370 38092 41372
rect 38116 41370 38172 41372
rect 38196 41370 38252 41372
rect 37956 41318 38002 41370
rect 38002 41318 38012 41370
rect 38036 41318 38066 41370
rect 38066 41318 38078 41370
rect 38078 41318 38092 41370
rect 38116 41318 38130 41370
rect 38130 41318 38142 41370
rect 38142 41318 38172 41370
rect 38196 41318 38206 41370
rect 38206 41318 38252 41370
rect 37956 41316 38012 41318
rect 38036 41316 38092 41318
rect 38116 41316 38172 41318
rect 38196 41316 38252 41318
rect 37956 40282 38012 40284
rect 38036 40282 38092 40284
rect 38116 40282 38172 40284
rect 38196 40282 38252 40284
rect 37956 40230 38002 40282
rect 38002 40230 38012 40282
rect 38036 40230 38066 40282
rect 38066 40230 38078 40282
rect 38078 40230 38092 40282
rect 38116 40230 38130 40282
rect 38130 40230 38142 40282
rect 38142 40230 38172 40282
rect 38196 40230 38206 40282
rect 38206 40230 38252 40282
rect 37956 40228 38012 40230
rect 38036 40228 38092 40230
rect 38116 40228 38172 40230
rect 38196 40228 38252 40230
rect 37956 39194 38012 39196
rect 38036 39194 38092 39196
rect 38116 39194 38172 39196
rect 38196 39194 38252 39196
rect 37956 39142 38002 39194
rect 38002 39142 38012 39194
rect 38036 39142 38066 39194
rect 38066 39142 38078 39194
rect 38078 39142 38092 39194
rect 38116 39142 38130 39194
rect 38130 39142 38142 39194
rect 38142 39142 38172 39194
rect 38196 39142 38206 39194
rect 38206 39142 38252 39194
rect 37956 39140 38012 39142
rect 38036 39140 38092 39142
rect 38116 39140 38172 39142
rect 38196 39140 38252 39142
rect 38106 38956 38162 38992
rect 38106 38936 38108 38956
rect 38108 38936 38160 38956
rect 38160 38936 38162 38956
rect 38474 38256 38530 38312
rect 37956 38106 38012 38108
rect 38036 38106 38092 38108
rect 38116 38106 38172 38108
rect 38196 38106 38252 38108
rect 37956 38054 38002 38106
rect 38002 38054 38012 38106
rect 38036 38054 38066 38106
rect 38066 38054 38078 38106
rect 38078 38054 38092 38106
rect 38116 38054 38130 38106
rect 38130 38054 38142 38106
rect 38142 38054 38172 38106
rect 38196 38054 38206 38106
rect 38206 38054 38252 38106
rect 37956 38052 38012 38054
rect 38036 38052 38092 38054
rect 38116 38052 38172 38054
rect 38196 38052 38252 38054
rect 37646 37068 37648 37088
rect 37648 37068 37700 37088
rect 37700 37068 37702 37088
rect 37646 37032 37702 37068
rect 37956 37018 38012 37020
rect 38036 37018 38092 37020
rect 38116 37018 38172 37020
rect 38196 37018 38252 37020
rect 37956 36966 38002 37018
rect 38002 36966 38012 37018
rect 38036 36966 38066 37018
rect 38066 36966 38078 37018
rect 38078 36966 38092 37018
rect 38116 36966 38130 37018
rect 38130 36966 38142 37018
rect 38142 36966 38172 37018
rect 38196 36966 38206 37018
rect 38206 36966 38252 37018
rect 37956 36964 38012 36966
rect 38036 36964 38092 36966
rect 38116 36964 38172 36966
rect 38196 36964 38252 36966
rect 37956 35930 38012 35932
rect 38036 35930 38092 35932
rect 38116 35930 38172 35932
rect 38196 35930 38252 35932
rect 37956 35878 38002 35930
rect 38002 35878 38012 35930
rect 38036 35878 38066 35930
rect 38066 35878 38078 35930
rect 38078 35878 38092 35930
rect 38116 35878 38130 35930
rect 38130 35878 38142 35930
rect 38142 35878 38172 35930
rect 38196 35878 38206 35930
rect 38206 35878 38252 35930
rect 37956 35876 38012 35878
rect 38036 35876 38092 35878
rect 38116 35876 38172 35878
rect 38196 35876 38252 35878
rect 37956 34842 38012 34844
rect 38036 34842 38092 34844
rect 38116 34842 38172 34844
rect 38196 34842 38252 34844
rect 37956 34790 38002 34842
rect 38002 34790 38012 34842
rect 38036 34790 38066 34842
rect 38066 34790 38078 34842
rect 38078 34790 38092 34842
rect 38116 34790 38130 34842
rect 38130 34790 38142 34842
rect 38142 34790 38172 34842
rect 38196 34790 38206 34842
rect 38206 34790 38252 34842
rect 37956 34788 38012 34790
rect 38036 34788 38092 34790
rect 38116 34788 38172 34790
rect 38196 34788 38252 34790
rect 37956 33754 38012 33756
rect 38036 33754 38092 33756
rect 38116 33754 38172 33756
rect 38196 33754 38252 33756
rect 37956 33702 38002 33754
rect 38002 33702 38012 33754
rect 38036 33702 38066 33754
rect 38066 33702 38078 33754
rect 38078 33702 38092 33754
rect 38116 33702 38130 33754
rect 38130 33702 38142 33754
rect 38142 33702 38172 33754
rect 38196 33702 38206 33754
rect 38206 33702 38252 33754
rect 37956 33700 38012 33702
rect 38036 33700 38092 33702
rect 38116 33700 38172 33702
rect 38196 33700 38252 33702
rect 37956 32666 38012 32668
rect 38036 32666 38092 32668
rect 38116 32666 38172 32668
rect 38196 32666 38252 32668
rect 37956 32614 38002 32666
rect 38002 32614 38012 32666
rect 38036 32614 38066 32666
rect 38066 32614 38078 32666
rect 38078 32614 38092 32666
rect 38116 32614 38130 32666
rect 38130 32614 38142 32666
rect 38142 32614 38172 32666
rect 38196 32614 38206 32666
rect 38206 32614 38252 32666
rect 37956 32612 38012 32614
rect 38036 32612 38092 32614
rect 38116 32612 38172 32614
rect 38196 32612 38252 32614
rect 37956 31578 38012 31580
rect 38036 31578 38092 31580
rect 38116 31578 38172 31580
rect 38196 31578 38252 31580
rect 37956 31526 38002 31578
rect 38002 31526 38012 31578
rect 38036 31526 38066 31578
rect 38066 31526 38078 31578
rect 38078 31526 38092 31578
rect 38116 31526 38130 31578
rect 38130 31526 38142 31578
rect 38142 31526 38172 31578
rect 38196 31526 38206 31578
rect 38206 31526 38252 31578
rect 37956 31524 38012 31526
rect 38036 31524 38092 31526
rect 38116 31524 38172 31526
rect 38196 31524 38252 31526
rect 37956 30490 38012 30492
rect 38036 30490 38092 30492
rect 38116 30490 38172 30492
rect 38196 30490 38252 30492
rect 37956 30438 38002 30490
rect 38002 30438 38012 30490
rect 38036 30438 38066 30490
rect 38066 30438 38078 30490
rect 38078 30438 38092 30490
rect 38116 30438 38130 30490
rect 38130 30438 38142 30490
rect 38142 30438 38172 30490
rect 38196 30438 38206 30490
rect 38206 30438 38252 30490
rect 37956 30436 38012 30438
rect 38036 30436 38092 30438
rect 38116 30436 38172 30438
rect 38196 30436 38252 30438
rect 37956 29402 38012 29404
rect 38036 29402 38092 29404
rect 38116 29402 38172 29404
rect 38196 29402 38252 29404
rect 37956 29350 38002 29402
rect 38002 29350 38012 29402
rect 38036 29350 38066 29402
rect 38066 29350 38078 29402
rect 38078 29350 38092 29402
rect 38116 29350 38130 29402
rect 38130 29350 38142 29402
rect 38142 29350 38172 29402
rect 38196 29350 38206 29402
rect 38206 29350 38252 29402
rect 37956 29348 38012 29350
rect 38036 29348 38092 29350
rect 38116 29348 38172 29350
rect 38196 29348 38252 29350
rect 37956 28314 38012 28316
rect 38036 28314 38092 28316
rect 38116 28314 38172 28316
rect 38196 28314 38252 28316
rect 37956 28262 38002 28314
rect 38002 28262 38012 28314
rect 38036 28262 38066 28314
rect 38066 28262 38078 28314
rect 38078 28262 38092 28314
rect 38116 28262 38130 28314
rect 38130 28262 38142 28314
rect 38142 28262 38172 28314
rect 38196 28262 38206 28314
rect 38206 28262 38252 28314
rect 37956 28260 38012 28262
rect 38036 28260 38092 28262
rect 38116 28260 38172 28262
rect 38196 28260 38252 28262
rect 37956 27226 38012 27228
rect 38036 27226 38092 27228
rect 38116 27226 38172 27228
rect 38196 27226 38252 27228
rect 37956 27174 38002 27226
rect 38002 27174 38012 27226
rect 38036 27174 38066 27226
rect 38066 27174 38078 27226
rect 38078 27174 38092 27226
rect 38116 27174 38130 27226
rect 38130 27174 38142 27226
rect 38142 27174 38172 27226
rect 38196 27174 38206 27226
rect 38206 27174 38252 27226
rect 37956 27172 38012 27174
rect 38036 27172 38092 27174
rect 38116 27172 38172 27174
rect 38196 27172 38252 27174
rect 37956 26138 38012 26140
rect 38036 26138 38092 26140
rect 38116 26138 38172 26140
rect 38196 26138 38252 26140
rect 37956 26086 38002 26138
rect 38002 26086 38012 26138
rect 38036 26086 38066 26138
rect 38066 26086 38078 26138
rect 38078 26086 38092 26138
rect 38116 26086 38130 26138
rect 38130 26086 38142 26138
rect 38142 26086 38172 26138
rect 38196 26086 38206 26138
rect 38206 26086 38252 26138
rect 37956 26084 38012 26086
rect 38036 26084 38092 26086
rect 38116 26084 38172 26086
rect 38196 26084 38252 26086
rect 37956 25050 38012 25052
rect 38036 25050 38092 25052
rect 38116 25050 38172 25052
rect 38196 25050 38252 25052
rect 37956 24998 38002 25050
rect 38002 24998 38012 25050
rect 38036 24998 38066 25050
rect 38066 24998 38078 25050
rect 38078 24998 38092 25050
rect 38116 24998 38130 25050
rect 38130 24998 38142 25050
rect 38142 24998 38172 25050
rect 38196 24998 38206 25050
rect 38206 24998 38252 25050
rect 37956 24996 38012 24998
rect 38036 24996 38092 24998
rect 38116 24996 38172 24998
rect 38196 24996 38252 24998
rect 42956 47354 43012 47356
rect 43036 47354 43092 47356
rect 43116 47354 43172 47356
rect 43196 47354 43252 47356
rect 42956 47302 43002 47354
rect 43002 47302 43012 47354
rect 43036 47302 43066 47354
rect 43066 47302 43078 47354
rect 43078 47302 43092 47354
rect 43116 47302 43130 47354
rect 43130 47302 43142 47354
rect 43142 47302 43172 47354
rect 43196 47302 43206 47354
rect 43206 47302 43252 47354
rect 42956 47300 43012 47302
rect 43036 47300 43092 47302
rect 43116 47300 43172 47302
rect 43196 47300 43252 47302
rect 42956 46266 43012 46268
rect 43036 46266 43092 46268
rect 43116 46266 43172 46268
rect 43196 46266 43252 46268
rect 42956 46214 43002 46266
rect 43002 46214 43012 46266
rect 43036 46214 43066 46266
rect 43066 46214 43078 46266
rect 43078 46214 43092 46266
rect 43116 46214 43130 46266
rect 43130 46214 43142 46266
rect 43142 46214 43172 46266
rect 43196 46214 43206 46266
rect 43206 46214 43252 46266
rect 42956 46212 43012 46214
rect 43036 46212 43092 46214
rect 43116 46212 43172 46214
rect 43196 46212 43252 46214
rect 42956 45178 43012 45180
rect 43036 45178 43092 45180
rect 43116 45178 43172 45180
rect 43196 45178 43252 45180
rect 42956 45126 43002 45178
rect 43002 45126 43012 45178
rect 43036 45126 43066 45178
rect 43066 45126 43078 45178
rect 43078 45126 43092 45178
rect 43116 45126 43130 45178
rect 43130 45126 43142 45178
rect 43142 45126 43172 45178
rect 43196 45126 43206 45178
rect 43206 45126 43252 45178
rect 42956 45124 43012 45126
rect 43036 45124 43092 45126
rect 43116 45124 43172 45126
rect 43196 45124 43252 45126
rect 47956 52250 48012 52252
rect 48036 52250 48092 52252
rect 48116 52250 48172 52252
rect 48196 52250 48252 52252
rect 47956 52198 48002 52250
rect 48002 52198 48012 52250
rect 48036 52198 48066 52250
rect 48066 52198 48078 52250
rect 48078 52198 48092 52250
rect 48116 52198 48130 52250
rect 48130 52198 48142 52250
rect 48142 52198 48172 52250
rect 48196 52198 48206 52250
rect 48206 52198 48252 52250
rect 47956 52196 48012 52198
rect 48036 52196 48092 52198
rect 48116 52196 48172 52198
rect 48196 52196 48252 52198
rect 48502 52128 48558 52184
rect 48502 51348 48504 51368
rect 48504 51348 48556 51368
rect 48556 51348 48558 51368
rect 48502 51312 48558 51348
rect 47956 51162 48012 51164
rect 48036 51162 48092 51164
rect 48116 51162 48172 51164
rect 48196 51162 48252 51164
rect 47956 51110 48002 51162
rect 48002 51110 48012 51162
rect 48036 51110 48066 51162
rect 48066 51110 48078 51162
rect 48078 51110 48092 51162
rect 48116 51110 48130 51162
rect 48130 51110 48142 51162
rect 48142 51110 48172 51162
rect 48196 51110 48206 51162
rect 48206 51110 48252 51162
rect 47956 51108 48012 51110
rect 48036 51108 48092 51110
rect 48116 51108 48172 51110
rect 48196 51108 48252 51110
rect 47956 50074 48012 50076
rect 48036 50074 48092 50076
rect 48116 50074 48172 50076
rect 48196 50074 48252 50076
rect 47956 50022 48002 50074
rect 48002 50022 48012 50074
rect 48036 50022 48066 50074
rect 48066 50022 48078 50074
rect 48078 50022 48092 50074
rect 48116 50022 48130 50074
rect 48130 50022 48142 50074
rect 48142 50022 48172 50074
rect 48196 50022 48206 50074
rect 48206 50022 48252 50074
rect 47956 50020 48012 50022
rect 48036 50020 48092 50022
rect 48116 50020 48172 50022
rect 48196 50020 48252 50022
rect 47956 48986 48012 48988
rect 48036 48986 48092 48988
rect 48116 48986 48172 48988
rect 48196 48986 48252 48988
rect 47956 48934 48002 48986
rect 48002 48934 48012 48986
rect 48036 48934 48066 48986
rect 48066 48934 48078 48986
rect 48078 48934 48092 48986
rect 48116 48934 48130 48986
rect 48130 48934 48142 48986
rect 48142 48934 48172 48986
rect 48196 48934 48206 48986
rect 48206 48934 48252 48986
rect 47956 48932 48012 48934
rect 48036 48932 48092 48934
rect 48116 48932 48172 48934
rect 48196 48932 48252 48934
rect 47956 47898 48012 47900
rect 48036 47898 48092 47900
rect 48116 47898 48172 47900
rect 48196 47898 48252 47900
rect 47956 47846 48002 47898
rect 48002 47846 48012 47898
rect 48036 47846 48066 47898
rect 48066 47846 48078 47898
rect 48078 47846 48092 47898
rect 48116 47846 48130 47898
rect 48130 47846 48142 47898
rect 48142 47846 48172 47898
rect 48196 47846 48206 47898
rect 48206 47846 48252 47898
rect 47956 47844 48012 47846
rect 48036 47844 48092 47846
rect 48116 47844 48172 47846
rect 48196 47844 48252 47846
rect 49330 50496 49386 50552
rect 49330 49680 49386 49736
rect 49054 48864 49110 48920
rect 49330 48084 49332 48104
rect 49332 48084 49384 48104
rect 49384 48084 49386 48104
rect 49330 48048 49386 48084
rect 49330 47232 49386 47288
rect 47956 46810 48012 46812
rect 48036 46810 48092 46812
rect 48116 46810 48172 46812
rect 48196 46810 48252 46812
rect 47956 46758 48002 46810
rect 48002 46758 48012 46810
rect 48036 46758 48066 46810
rect 48066 46758 48078 46810
rect 48078 46758 48092 46810
rect 48116 46758 48130 46810
rect 48130 46758 48142 46810
rect 48142 46758 48172 46810
rect 48196 46758 48206 46810
rect 48206 46758 48252 46810
rect 47956 46756 48012 46758
rect 48036 46756 48092 46758
rect 48116 46756 48172 46758
rect 48196 46756 48252 46758
rect 49054 46416 49110 46472
rect 47956 45722 48012 45724
rect 48036 45722 48092 45724
rect 48116 45722 48172 45724
rect 48196 45722 48252 45724
rect 47956 45670 48002 45722
rect 48002 45670 48012 45722
rect 48036 45670 48066 45722
rect 48066 45670 48078 45722
rect 48078 45670 48092 45722
rect 48116 45670 48130 45722
rect 48130 45670 48142 45722
rect 48142 45670 48172 45722
rect 48196 45670 48206 45722
rect 48206 45670 48252 45722
rect 47956 45668 48012 45670
rect 48036 45668 48092 45670
rect 48116 45668 48172 45670
rect 48196 45668 48252 45670
rect 39670 39888 39726 39944
rect 42956 44090 43012 44092
rect 43036 44090 43092 44092
rect 43116 44090 43172 44092
rect 43196 44090 43252 44092
rect 42956 44038 43002 44090
rect 43002 44038 43012 44090
rect 43036 44038 43066 44090
rect 43066 44038 43078 44090
rect 43078 44038 43092 44090
rect 43116 44038 43130 44090
rect 43130 44038 43142 44090
rect 43142 44038 43172 44090
rect 43196 44038 43206 44090
rect 43206 44038 43252 44090
rect 42956 44036 43012 44038
rect 43036 44036 43092 44038
rect 43116 44036 43172 44038
rect 43196 44036 43252 44038
rect 42956 43002 43012 43004
rect 43036 43002 43092 43004
rect 43116 43002 43172 43004
rect 43196 43002 43252 43004
rect 42956 42950 43002 43002
rect 43002 42950 43012 43002
rect 43036 42950 43066 43002
rect 43066 42950 43078 43002
rect 43078 42950 43092 43002
rect 43116 42950 43130 43002
rect 43130 42950 43142 43002
rect 43142 42950 43172 43002
rect 43196 42950 43206 43002
rect 43206 42950 43252 43002
rect 42956 42948 43012 42950
rect 43036 42948 43092 42950
rect 43116 42948 43172 42950
rect 43196 42948 43252 42950
rect 42956 41914 43012 41916
rect 43036 41914 43092 41916
rect 43116 41914 43172 41916
rect 43196 41914 43252 41916
rect 42956 41862 43002 41914
rect 43002 41862 43012 41914
rect 43036 41862 43066 41914
rect 43066 41862 43078 41914
rect 43078 41862 43092 41914
rect 43116 41862 43130 41914
rect 43130 41862 43142 41914
rect 43142 41862 43172 41914
rect 43196 41862 43206 41914
rect 43206 41862 43252 41914
rect 42956 41860 43012 41862
rect 43036 41860 43092 41862
rect 43116 41860 43172 41862
rect 43196 41860 43252 41862
rect 42956 40826 43012 40828
rect 43036 40826 43092 40828
rect 43116 40826 43172 40828
rect 43196 40826 43252 40828
rect 42956 40774 43002 40826
rect 43002 40774 43012 40826
rect 43036 40774 43066 40826
rect 43066 40774 43078 40826
rect 43078 40774 43092 40826
rect 43116 40774 43130 40826
rect 43130 40774 43142 40826
rect 43142 40774 43172 40826
rect 43196 40774 43206 40826
rect 43206 40774 43252 40826
rect 42956 40772 43012 40774
rect 43036 40772 43092 40774
rect 43116 40772 43172 40774
rect 43196 40772 43252 40774
rect 49054 45600 49110 45656
rect 49054 44820 49056 44840
rect 49056 44820 49108 44840
rect 49108 44820 49110 44840
rect 49054 44784 49110 44820
rect 47956 44634 48012 44636
rect 48036 44634 48092 44636
rect 48116 44634 48172 44636
rect 48196 44634 48252 44636
rect 47956 44582 48002 44634
rect 48002 44582 48012 44634
rect 48036 44582 48066 44634
rect 48066 44582 48078 44634
rect 48078 44582 48092 44634
rect 48116 44582 48130 44634
rect 48130 44582 48142 44634
rect 48142 44582 48172 44634
rect 48196 44582 48206 44634
rect 48206 44582 48252 44634
rect 47956 44580 48012 44582
rect 48036 44580 48092 44582
rect 48116 44580 48172 44582
rect 48196 44580 48252 44582
rect 49330 43968 49386 44024
rect 47956 43546 48012 43548
rect 48036 43546 48092 43548
rect 48116 43546 48172 43548
rect 48196 43546 48252 43548
rect 47956 43494 48002 43546
rect 48002 43494 48012 43546
rect 48036 43494 48066 43546
rect 48066 43494 48078 43546
rect 48078 43494 48092 43546
rect 48116 43494 48130 43546
rect 48130 43494 48142 43546
rect 48142 43494 48172 43546
rect 48196 43494 48206 43546
rect 48206 43494 48252 43546
rect 47956 43492 48012 43494
rect 48036 43492 48092 43494
rect 48116 43492 48172 43494
rect 48196 43492 48252 43494
rect 49146 43152 49202 43208
rect 47956 42458 48012 42460
rect 48036 42458 48092 42460
rect 48116 42458 48172 42460
rect 48196 42458 48252 42460
rect 47956 42406 48002 42458
rect 48002 42406 48012 42458
rect 48036 42406 48066 42458
rect 48066 42406 48078 42458
rect 48078 42406 48092 42458
rect 48116 42406 48130 42458
rect 48130 42406 48142 42458
rect 48142 42406 48172 42458
rect 48196 42406 48206 42458
rect 48206 42406 48252 42458
rect 47956 42404 48012 42406
rect 48036 42404 48092 42406
rect 48116 42404 48172 42406
rect 48196 42404 48252 42406
rect 49054 42336 49110 42392
rect 49054 41556 49056 41576
rect 49056 41556 49108 41576
rect 49108 41556 49110 41576
rect 49054 41520 49110 41556
rect 47956 41370 48012 41372
rect 48036 41370 48092 41372
rect 48116 41370 48172 41372
rect 48196 41370 48252 41372
rect 47956 41318 48002 41370
rect 48002 41318 48012 41370
rect 48036 41318 48066 41370
rect 48066 41318 48078 41370
rect 48078 41318 48092 41370
rect 48116 41318 48130 41370
rect 48130 41318 48142 41370
rect 48142 41318 48172 41370
rect 48196 41318 48206 41370
rect 48206 41318 48252 41370
rect 47956 41316 48012 41318
rect 48036 41316 48092 41318
rect 48116 41316 48172 41318
rect 48196 41316 48252 41318
rect 47956 40282 48012 40284
rect 48036 40282 48092 40284
rect 48116 40282 48172 40284
rect 48196 40282 48252 40284
rect 47956 40230 48002 40282
rect 48002 40230 48012 40282
rect 48036 40230 48066 40282
rect 48066 40230 48078 40282
rect 48078 40230 48092 40282
rect 48116 40230 48130 40282
rect 48130 40230 48142 40282
rect 48142 40230 48172 40282
rect 48196 40230 48206 40282
rect 48206 40230 48252 40282
rect 47956 40228 48012 40230
rect 48036 40228 48092 40230
rect 48116 40228 48172 40230
rect 48196 40228 48252 40230
rect 49054 39888 49110 39944
rect 42956 39738 43012 39740
rect 43036 39738 43092 39740
rect 43116 39738 43172 39740
rect 43196 39738 43252 39740
rect 42956 39686 43002 39738
rect 43002 39686 43012 39738
rect 43036 39686 43066 39738
rect 43066 39686 43078 39738
rect 43078 39686 43092 39738
rect 43116 39686 43130 39738
rect 43130 39686 43142 39738
rect 43142 39686 43172 39738
rect 43196 39686 43206 39738
rect 43206 39686 43252 39738
rect 42956 39684 43012 39686
rect 43036 39684 43092 39686
rect 43116 39684 43172 39686
rect 43196 39684 43252 39686
rect 40130 38800 40186 38856
rect 49330 40704 49386 40760
rect 47956 39194 48012 39196
rect 48036 39194 48092 39196
rect 48116 39194 48172 39196
rect 48196 39194 48252 39196
rect 47956 39142 48002 39194
rect 48002 39142 48012 39194
rect 48036 39142 48066 39194
rect 48066 39142 48078 39194
rect 48078 39142 48092 39194
rect 48116 39142 48130 39194
rect 48130 39142 48142 39194
rect 48142 39142 48172 39194
rect 48196 39142 48206 39194
rect 48206 39142 48252 39194
rect 47956 39140 48012 39142
rect 48036 39140 48092 39142
rect 48116 39140 48172 39142
rect 48196 39140 48252 39142
rect 49146 39072 49202 39128
rect 42956 38650 43012 38652
rect 43036 38650 43092 38652
rect 43116 38650 43172 38652
rect 43196 38650 43252 38652
rect 42956 38598 43002 38650
rect 43002 38598 43012 38650
rect 43036 38598 43066 38650
rect 43066 38598 43078 38650
rect 43078 38598 43092 38650
rect 43116 38598 43130 38650
rect 43130 38598 43142 38650
rect 43142 38598 43172 38650
rect 43196 38598 43206 38650
rect 43206 38598 43252 38650
rect 42956 38596 43012 38598
rect 43036 38596 43092 38598
rect 43116 38596 43172 38598
rect 43196 38596 43252 38598
rect 49146 38276 49202 38312
rect 49146 38256 49148 38276
rect 49148 38256 49200 38276
rect 49200 38256 49202 38276
rect 47956 38106 48012 38108
rect 48036 38106 48092 38108
rect 48116 38106 48172 38108
rect 48196 38106 48252 38108
rect 47956 38054 48002 38106
rect 48002 38054 48012 38106
rect 48036 38054 48066 38106
rect 48066 38054 48078 38106
rect 48078 38054 48092 38106
rect 48116 38054 48130 38106
rect 48130 38054 48142 38106
rect 48142 38054 48172 38106
rect 48196 38054 48206 38106
rect 48206 38054 48252 38106
rect 47956 38052 48012 38054
rect 48036 38052 48092 38054
rect 48116 38052 48172 38054
rect 48196 38052 48252 38054
rect 42956 37562 43012 37564
rect 43036 37562 43092 37564
rect 43116 37562 43172 37564
rect 43196 37562 43252 37564
rect 42956 37510 43002 37562
rect 43002 37510 43012 37562
rect 43036 37510 43066 37562
rect 43066 37510 43078 37562
rect 43078 37510 43092 37562
rect 43116 37510 43130 37562
rect 43130 37510 43142 37562
rect 43142 37510 43172 37562
rect 43196 37510 43206 37562
rect 43206 37510 43252 37562
rect 42956 37508 43012 37510
rect 43036 37508 43092 37510
rect 43116 37508 43172 37510
rect 43196 37508 43252 37510
rect 49330 37440 49386 37496
rect 47956 37018 48012 37020
rect 48036 37018 48092 37020
rect 48116 37018 48172 37020
rect 48196 37018 48252 37020
rect 47956 36966 48002 37018
rect 48002 36966 48012 37018
rect 48036 36966 48066 37018
rect 48066 36966 48078 37018
rect 48078 36966 48092 37018
rect 48116 36966 48130 37018
rect 48130 36966 48142 37018
rect 48142 36966 48172 37018
rect 48196 36966 48206 37018
rect 48206 36966 48252 37018
rect 47956 36964 48012 36966
rect 48036 36964 48092 36966
rect 48116 36964 48172 36966
rect 48196 36964 48252 36966
rect 42956 36474 43012 36476
rect 43036 36474 43092 36476
rect 43116 36474 43172 36476
rect 43196 36474 43252 36476
rect 42956 36422 43002 36474
rect 43002 36422 43012 36474
rect 43036 36422 43066 36474
rect 43066 36422 43078 36474
rect 43078 36422 43092 36474
rect 43116 36422 43130 36474
rect 43130 36422 43142 36474
rect 43142 36422 43172 36474
rect 43196 36422 43206 36474
rect 43206 36422 43252 36474
rect 42956 36420 43012 36422
rect 43036 36420 43092 36422
rect 43116 36420 43172 36422
rect 43196 36420 43252 36422
rect 42956 35386 43012 35388
rect 43036 35386 43092 35388
rect 43116 35386 43172 35388
rect 43196 35386 43252 35388
rect 42956 35334 43002 35386
rect 43002 35334 43012 35386
rect 43036 35334 43066 35386
rect 43066 35334 43078 35386
rect 43078 35334 43092 35386
rect 43116 35334 43130 35386
rect 43130 35334 43142 35386
rect 43142 35334 43172 35386
rect 43196 35334 43206 35386
rect 43206 35334 43252 35386
rect 42956 35332 43012 35334
rect 43036 35332 43092 35334
rect 43116 35332 43172 35334
rect 43196 35332 43252 35334
rect 48318 36644 48374 36680
rect 48318 36624 48320 36644
rect 48320 36624 48372 36644
rect 48372 36624 48374 36644
rect 49054 36624 49110 36680
rect 47956 35930 48012 35932
rect 48036 35930 48092 35932
rect 48116 35930 48172 35932
rect 48196 35930 48252 35932
rect 47956 35878 48002 35930
rect 48002 35878 48012 35930
rect 48036 35878 48066 35930
rect 48066 35878 48078 35930
rect 48078 35878 48092 35930
rect 48116 35878 48130 35930
rect 48130 35878 48142 35930
rect 48142 35878 48172 35930
rect 48196 35878 48206 35930
rect 48206 35878 48252 35930
rect 47956 35876 48012 35878
rect 48036 35876 48092 35878
rect 48116 35876 48172 35878
rect 48196 35876 48252 35878
rect 48410 35808 48466 35864
rect 48318 34992 48374 35048
rect 49054 35028 49056 35048
rect 49056 35028 49108 35048
rect 49108 35028 49110 35048
rect 49054 34992 49110 35028
rect 47956 34842 48012 34844
rect 48036 34842 48092 34844
rect 48116 34842 48172 34844
rect 48196 34842 48252 34844
rect 47956 34790 48002 34842
rect 48002 34790 48012 34842
rect 48036 34790 48066 34842
rect 48066 34790 48078 34842
rect 48078 34790 48092 34842
rect 48116 34790 48130 34842
rect 48130 34790 48142 34842
rect 48142 34790 48172 34842
rect 48196 34790 48206 34842
rect 48206 34790 48252 34842
rect 47956 34788 48012 34790
rect 48036 34788 48092 34790
rect 48116 34788 48172 34790
rect 48196 34788 48252 34790
rect 42956 34298 43012 34300
rect 43036 34298 43092 34300
rect 43116 34298 43172 34300
rect 43196 34298 43252 34300
rect 42956 34246 43002 34298
rect 43002 34246 43012 34298
rect 43036 34246 43066 34298
rect 43066 34246 43078 34298
rect 43078 34246 43092 34298
rect 43116 34246 43130 34298
rect 43130 34246 43142 34298
rect 43142 34246 43172 34298
rect 43196 34246 43206 34298
rect 43206 34246 43252 34298
rect 42956 34244 43012 34246
rect 43036 34244 43092 34246
rect 43116 34244 43172 34246
rect 43196 34244 43252 34246
rect 42956 33210 43012 33212
rect 43036 33210 43092 33212
rect 43116 33210 43172 33212
rect 43196 33210 43252 33212
rect 42956 33158 43002 33210
rect 43002 33158 43012 33210
rect 43036 33158 43066 33210
rect 43066 33158 43078 33210
rect 43078 33158 43092 33210
rect 43116 33158 43130 33210
rect 43130 33158 43142 33210
rect 43142 33158 43172 33210
rect 43196 33158 43206 33210
rect 43206 33158 43252 33210
rect 42956 33156 43012 33158
rect 43036 33156 43092 33158
rect 43116 33156 43172 33158
rect 43196 33156 43252 33158
rect 42956 32122 43012 32124
rect 43036 32122 43092 32124
rect 43116 32122 43172 32124
rect 43196 32122 43252 32124
rect 42956 32070 43002 32122
rect 43002 32070 43012 32122
rect 43036 32070 43066 32122
rect 43066 32070 43078 32122
rect 43078 32070 43092 32122
rect 43116 32070 43130 32122
rect 43130 32070 43142 32122
rect 43142 32070 43172 32122
rect 43196 32070 43206 32122
rect 43206 32070 43252 32122
rect 42956 32068 43012 32070
rect 43036 32068 43092 32070
rect 43116 32068 43172 32070
rect 43196 32068 43252 32070
rect 42956 31034 43012 31036
rect 43036 31034 43092 31036
rect 43116 31034 43172 31036
rect 43196 31034 43252 31036
rect 42956 30982 43002 31034
rect 43002 30982 43012 31034
rect 43036 30982 43066 31034
rect 43066 30982 43078 31034
rect 43078 30982 43092 31034
rect 43116 30982 43130 31034
rect 43130 30982 43142 31034
rect 43142 30982 43172 31034
rect 43196 30982 43206 31034
rect 43206 30982 43252 31034
rect 42956 30980 43012 30982
rect 43036 30980 43092 30982
rect 43116 30980 43172 30982
rect 43196 30980 43252 30982
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 42956 29946 43012 29948
rect 43036 29946 43092 29948
rect 43116 29946 43172 29948
rect 43196 29946 43252 29948
rect 42956 29894 43002 29946
rect 43002 29894 43012 29946
rect 43036 29894 43066 29946
rect 43066 29894 43078 29946
rect 43078 29894 43092 29946
rect 43116 29894 43130 29946
rect 43130 29894 43142 29946
rect 43142 29894 43172 29946
rect 43196 29894 43206 29946
rect 43206 29894 43252 29946
rect 42956 29892 43012 29894
rect 43036 29892 43092 29894
rect 43116 29892 43172 29894
rect 43196 29892 43252 29894
rect 42956 28858 43012 28860
rect 43036 28858 43092 28860
rect 43116 28858 43172 28860
rect 43196 28858 43252 28860
rect 42956 28806 43002 28858
rect 43002 28806 43012 28858
rect 43036 28806 43066 28858
rect 43066 28806 43078 28858
rect 43078 28806 43092 28858
rect 43116 28806 43130 28858
rect 43130 28806 43142 28858
rect 43142 28806 43172 28858
rect 43196 28806 43206 28858
rect 43206 28806 43252 28858
rect 42956 28804 43012 28806
rect 43036 28804 43092 28806
rect 43116 28804 43172 28806
rect 43196 28804 43252 28806
rect 42956 27770 43012 27772
rect 43036 27770 43092 27772
rect 43116 27770 43172 27772
rect 43196 27770 43252 27772
rect 42956 27718 43002 27770
rect 43002 27718 43012 27770
rect 43036 27718 43066 27770
rect 43066 27718 43078 27770
rect 43078 27718 43092 27770
rect 43116 27718 43130 27770
rect 43130 27718 43142 27770
rect 43142 27718 43172 27770
rect 43196 27718 43206 27770
rect 43206 27718 43252 27770
rect 42956 27716 43012 27718
rect 43036 27716 43092 27718
rect 43116 27716 43172 27718
rect 43196 27716 43252 27718
rect 42956 26682 43012 26684
rect 43036 26682 43092 26684
rect 43116 26682 43172 26684
rect 43196 26682 43252 26684
rect 42956 26630 43002 26682
rect 43002 26630 43012 26682
rect 43036 26630 43066 26682
rect 43066 26630 43078 26682
rect 43078 26630 43092 26682
rect 43116 26630 43130 26682
rect 43130 26630 43142 26682
rect 43142 26630 43172 26682
rect 43196 26630 43206 26682
rect 43206 26630 43252 26682
rect 42956 26628 43012 26630
rect 43036 26628 43092 26630
rect 43116 26628 43172 26630
rect 43196 26628 43252 26630
rect 42956 25594 43012 25596
rect 43036 25594 43092 25596
rect 43116 25594 43172 25596
rect 43196 25594 43252 25596
rect 42956 25542 43002 25594
rect 43002 25542 43012 25594
rect 43036 25542 43066 25594
rect 43066 25542 43078 25594
rect 43078 25542 43092 25594
rect 43116 25542 43130 25594
rect 43130 25542 43142 25594
rect 43142 25542 43172 25594
rect 43196 25542 43206 25594
rect 43206 25542 43252 25594
rect 42956 25540 43012 25542
rect 43036 25540 43092 25542
rect 43116 25540 43172 25542
rect 43196 25540 43252 25542
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 49330 34176 49386 34232
rect 47956 33754 48012 33756
rect 48036 33754 48092 33756
rect 48116 33754 48172 33756
rect 48196 33754 48252 33756
rect 47956 33702 48002 33754
rect 48002 33702 48012 33754
rect 48036 33702 48066 33754
rect 48066 33702 48078 33754
rect 48078 33702 48092 33754
rect 48116 33702 48130 33754
rect 48130 33702 48142 33754
rect 48142 33702 48172 33754
rect 48196 33702 48206 33754
rect 48206 33702 48252 33754
rect 47956 33700 48012 33702
rect 48036 33700 48092 33702
rect 48116 33700 48172 33702
rect 48196 33700 48252 33702
rect 49146 33360 49202 33416
rect 47956 32666 48012 32668
rect 48036 32666 48092 32668
rect 48116 32666 48172 32668
rect 48196 32666 48252 32668
rect 47956 32614 48002 32666
rect 48002 32614 48012 32666
rect 48036 32614 48066 32666
rect 48066 32614 48078 32666
rect 48078 32614 48092 32666
rect 48116 32614 48130 32666
rect 48130 32614 48142 32666
rect 48142 32614 48172 32666
rect 48196 32614 48206 32666
rect 48206 32614 48252 32666
rect 47956 32612 48012 32614
rect 48036 32612 48092 32614
rect 48116 32612 48172 32614
rect 48196 32612 48252 32614
rect 49054 32544 49110 32600
rect 49054 31764 49056 31784
rect 49056 31764 49108 31784
rect 49108 31764 49110 31784
rect 49054 31728 49110 31764
rect 47956 31578 48012 31580
rect 48036 31578 48092 31580
rect 48116 31578 48172 31580
rect 48196 31578 48252 31580
rect 47956 31526 48002 31578
rect 48002 31526 48012 31578
rect 48036 31526 48066 31578
rect 48066 31526 48078 31578
rect 48078 31526 48092 31578
rect 48116 31526 48130 31578
rect 48130 31526 48142 31578
rect 48142 31526 48172 31578
rect 48196 31526 48206 31578
rect 48206 31526 48252 31578
rect 47956 31524 48012 31526
rect 48036 31524 48092 31526
rect 48116 31524 48172 31526
rect 48196 31524 48252 31526
rect 49330 30912 49386 30968
rect 47956 30490 48012 30492
rect 48036 30490 48092 30492
rect 48116 30490 48172 30492
rect 48196 30490 48252 30492
rect 47956 30438 48002 30490
rect 48002 30438 48012 30490
rect 48036 30438 48066 30490
rect 48066 30438 48078 30490
rect 48078 30438 48092 30490
rect 48116 30438 48130 30490
rect 48130 30438 48142 30490
rect 48142 30438 48172 30490
rect 48196 30438 48206 30490
rect 48206 30438 48252 30490
rect 47956 30436 48012 30438
rect 48036 30436 48092 30438
rect 48116 30436 48172 30438
rect 48196 30436 48252 30438
rect 49054 30096 49110 30152
rect 47956 29402 48012 29404
rect 48036 29402 48092 29404
rect 48116 29402 48172 29404
rect 48196 29402 48252 29404
rect 47956 29350 48002 29402
rect 48002 29350 48012 29402
rect 48036 29350 48066 29402
rect 48066 29350 48078 29402
rect 48078 29350 48092 29402
rect 48116 29350 48130 29402
rect 48130 29350 48142 29402
rect 48142 29350 48172 29402
rect 48196 29350 48206 29402
rect 48206 29350 48252 29402
rect 47956 29348 48012 29350
rect 48036 29348 48092 29350
rect 48116 29348 48172 29350
rect 48196 29348 48252 29350
rect 49146 29280 49202 29336
rect 49054 28500 49056 28520
rect 49056 28500 49108 28520
rect 49108 28500 49110 28520
rect 49054 28464 49110 28500
rect 47956 28314 48012 28316
rect 48036 28314 48092 28316
rect 48116 28314 48172 28316
rect 48196 28314 48252 28316
rect 47956 28262 48002 28314
rect 48002 28262 48012 28314
rect 48036 28262 48066 28314
rect 48066 28262 48078 28314
rect 48078 28262 48092 28314
rect 48116 28262 48130 28314
rect 48130 28262 48142 28314
rect 48142 28262 48172 28314
rect 48196 28262 48206 28314
rect 48206 28262 48252 28314
rect 47956 28260 48012 28262
rect 48036 28260 48092 28262
rect 48116 28260 48172 28262
rect 48196 28260 48252 28262
rect 49330 27648 49386 27704
rect 47956 27226 48012 27228
rect 48036 27226 48092 27228
rect 48116 27226 48172 27228
rect 48196 27226 48252 27228
rect 47956 27174 48002 27226
rect 48002 27174 48012 27226
rect 48036 27174 48066 27226
rect 48066 27174 48078 27226
rect 48078 27174 48092 27226
rect 48116 27174 48130 27226
rect 48130 27174 48142 27226
rect 48142 27174 48172 27226
rect 48196 27174 48206 27226
rect 48206 27174 48252 27226
rect 47956 27172 48012 27174
rect 48036 27172 48092 27174
rect 48116 27172 48172 27174
rect 48196 27172 48252 27174
rect 49146 26868 49148 26888
rect 49148 26868 49200 26888
rect 49200 26868 49202 26888
rect 49146 26832 49202 26868
rect 47956 26138 48012 26140
rect 48036 26138 48092 26140
rect 48116 26138 48172 26140
rect 48196 26138 48252 26140
rect 47956 26086 48002 26138
rect 48002 26086 48012 26138
rect 48036 26086 48066 26138
rect 48066 26086 48078 26138
rect 48078 26086 48092 26138
rect 48116 26086 48130 26138
rect 48130 26086 48142 26138
rect 48142 26086 48172 26138
rect 48196 26086 48206 26138
rect 48206 26086 48252 26138
rect 47956 26084 48012 26086
rect 48036 26084 48092 26086
rect 48116 26084 48172 26086
rect 48196 26084 48252 26086
rect 48410 26016 48466 26072
rect 49146 25236 49148 25256
rect 49148 25236 49200 25256
rect 49200 25236 49202 25256
rect 49146 25200 49202 25236
rect 47956 25050 48012 25052
rect 48036 25050 48092 25052
rect 48116 25050 48172 25052
rect 48196 25050 48252 25052
rect 47956 24998 48002 25050
rect 48002 24998 48012 25050
rect 48036 24998 48066 25050
rect 48066 24998 48078 25050
rect 48078 24998 48092 25050
rect 48116 24998 48130 25050
rect 48130 24998 48142 25050
rect 48142 24998 48172 25050
rect 48196 24998 48206 25050
rect 48206 24998 48252 25050
rect 47956 24996 48012 24998
rect 48036 24996 48092 24998
rect 48116 24996 48172 24998
rect 48196 24996 48252 24998
rect 49146 24384 49202 24440
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 49146 23604 49148 23624
rect 49148 23604 49200 23624
rect 49200 23604 49202 23624
rect 49146 23568 49202 23604
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 49146 22752 49202 22808
rect 49146 21972 49148 21992
rect 49148 21972 49200 21992
rect 49200 21972 49202 21992
rect 49146 21936 49202 21972
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 49146 21120 49202 21176
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 49146 20340 49148 20360
rect 49148 20340 49200 20360
rect 49200 20340 49202 20360
rect 49146 20304 49202 20340
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 49146 19488 49202 19544
rect 49146 18708 49148 18728
rect 49148 18708 49200 18728
rect 49200 18708 49202 18728
rect 49146 18672 49202 18708
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 49146 17856 49202 17912
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49146 17076 49148 17096
rect 49148 17076 49200 17096
rect 49200 17076 49202 17096
rect 49146 17040 49202 17076
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 49146 16224 49202 16280
rect 49146 15444 49148 15464
rect 49148 15444 49200 15464
rect 49200 15444 49202 15464
rect 49146 15408 49202 15444
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 49146 14592 49202 14648
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 49146 13812 49148 13832
rect 49148 13812 49200 13832
rect 49200 13812 49202 13832
rect 49146 13776 49202 13812
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 49146 12960 49202 13016
rect 49146 12180 49148 12200
rect 49148 12180 49200 12200
rect 49200 12180 49202 12200
rect 49146 12144 49202 12180
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 49146 11328 49202 11384
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49146 10548 49148 10568
rect 49148 10548 49200 10568
rect 49200 10548 49202 10568
rect 49146 10512 49202 10548
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 49146 9696 49202 9752
rect 49146 8916 49148 8936
rect 49148 8916 49200 8936
rect 49200 8916 49202 8936
rect 49146 8880 49202 8916
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 49146 8064 49202 8120
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7284 49148 7304
rect 49148 7284 49200 7304
rect 49200 7284 49202 7304
rect 49146 7248 49202 7284
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 49146 6432 49202 6488
rect 49146 5652 49148 5672
rect 49148 5652 49200 5672
rect 49200 5652 49202 5672
rect 49146 5616 49202 5652
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 49146 4800 49202 4856
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 4020 49148 4040
rect 49148 4020 49200 4040
rect 49200 4020 49202 4040
rect 49146 3984 49202 4020
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
rect 49146 3168 49202 3224
rect 49146 2372 49202 2408
rect 49146 2352 49148 2372
rect 49148 2352 49200 2372
rect 49200 2352 49202 2372
<< metal3 >>
rect 0 54634 800 54664
rect 3417 54634 3483 54637
rect 0 54632 3483 54634
rect 0 54576 3422 54632
rect 3478 54576 3483 54632
rect 0 54574 3483 54576
rect 0 54544 800 54574
rect 3417 54571 3483 54574
rect 47761 54634 47827 54637
rect 50200 54634 51000 54664
rect 47761 54632 51000 54634
rect 47761 54576 47766 54632
rect 47822 54576 51000 54632
rect 47761 54574 51000 54576
rect 47761 54571 47827 54574
rect 50200 54544 51000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 27946 54432 28262 54433
rect 27946 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28262 54432
rect 27946 54367 28262 54368
rect 37946 54432 38262 54433
rect 37946 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38262 54432
rect 37946 54367 38262 54368
rect 47946 54432 48262 54433
rect 47946 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48262 54432
rect 47946 54367 48262 54368
rect 2946 53888 3262 53889
rect 0 53818 800 53848
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 32946 53888 33262 53889
rect 32946 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33262 53888
rect 32946 53823 33262 53824
rect 42946 53888 43262 53889
rect 42946 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43262 53888
rect 42946 53823 43262 53824
rect 48313 53818 48379 53821
rect 50200 53818 51000 53848
rect 0 53758 1778 53818
rect 0 53728 800 53758
rect 1718 53682 1778 53758
rect 48313 53816 51000 53818
rect 48313 53760 48318 53816
rect 48374 53760 51000 53816
rect 48313 53758 51000 53760
rect 48313 53755 48379 53758
rect 50200 53728 51000 53758
rect 3325 53682 3391 53685
rect 1718 53680 3391 53682
rect 1718 53624 3330 53680
rect 3386 53624 3391 53680
rect 1718 53622 3391 53624
rect 3325 53619 3391 53622
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 27946 53344 28262 53345
rect 27946 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28262 53344
rect 27946 53279 28262 53280
rect 37946 53344 38262 53345
rect 37946 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38262 53344
rect 37946 53279 38262 53280
rect 47946 53344 48262 53345
rect 47946 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48262 53344
rect 47946 53279 48262 53280
rect 0 53002 800 53032
rect 3601 53002 3667 53005
rect 0 53000 3667 53002
rect 0 52944 3606 53000
rect 3662 52944 3667 53000
rect 0 52942 3667 52944
rect 0 52912 800 52942
rect 3601 52939 3667 52942
rect 48497 53002 48563 53005
rect 50200 53002 51000 53032
rect 48497 53000 51000 53002
rect 48497 52944 48502 53000
rect 48558 52944 51000 53000
rect 48497 52942 51000 52944
rect 48497 52939 48563 52942
rect 50200 52912 51000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 32946 52800 33262 52801
rect 32946 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33262 52800
rect 32946 52735 33262 52736
rect 42946 52800 43262 52801
rect 42946 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43262 52800
rect 42946 52735 43262 52736
rect 7946 52256 8262 52257
rect 0 52186 800 52216
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 27946 52256 28262 52257
rect 27946 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28262 52256
rect 27946 52191 28262 52192
rect 37946 52256 38262 52257
rect 37946 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38262 52256
rect 37946 52191 38262 52192
rect 47946 52256 48262 52257
rect 47946 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48262 52256
rect 47946 52191 48262 52192
rect 48497 52186 48563 52189
rect 50200 52186 51000 52216
rect 0 52126 6930 52186
rect 0 52096 800 52126
rect 6870 52050 6930 52126
rect 48497 52184 51000 52186
rect 48497 52128 48502 52184
rect 48558 52128 51000 52184
rect 48497 52126 51000 52128
rect 48497 52123 48563 52126
rect 50200 52096 51000 52126
rect 21214 52050 21220 52052
rect 6870 51990 21220 52050
rect 21214 51988 21220 51990
rect 21284 51988 21290 52052
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 32946 51712 33262 51713
rect 32946 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33262 51712
rect 32946 51647 33262 51648
rect 42946 51712 43262 51713
rect 42946 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43262 51712
rect 42946 51647 43262 51648
rect 0 51370 800 51400
rect 1301 51370 1367 51373
rect 0 51368 1367 51370
rect 0 51312 1306 51368
rect 1362 51312 1367 51368
rect 0 51310 1367 51312
rect 0 51280 800 51310
rect 1301 51307 1367 51310
rect 48497 51370 48563 51373
rect 50200 51370 51000 51400
rect 48497 51368 51000 51370
rect 48497 51312 48502 51368
rect 48558 51312 51000 51368
rect 48497 51310 51000 51312
rect 48497 51307 48563 51310
rect 50200 51280 51000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 27946 51168 28262 51169
rect 27946 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28262 51168
rect 27946 51103 28262 51104
rect 37946 51168 38262 51169
rect 37946 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38262 51168
rect 37946 51103 38262 51104
rect 47946 51168 48262 51169
rect 47946 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48262 51168
rect 47946 51103 48262 51104
rect 2946 50624 3262 50625
rect 0 50554 800 50584
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 32946 50624 33262 50625
rect 32946 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33262 50624
rect 32946 50559 33262 50560
rect 42946 50624 43262 50625
rect 42946 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43262 50624
rect 42946 50559 43262 50560
rect 1301 50554 1367 50557
rect 0 50552 1367 50554
rect 0 50496 1306 50552
rect 1362 50496 1367 50552
rect 0 50494 1367 50496
rect 0 50464 800 50494
rect 1301 50491 1367 50494
rect 49325 50554 49391 50557
rect 50200 50554 51000 50584
rect 49325 50552 51000 50554
rect 49325 50496 49330 50552
rect 49386 50496 51000 50552
rect 49325 50494 51000 50496
rect 49325 50491 49391 50494
rect 50200 50464 51000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 27946 50080 28262 50081
rect 27946 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28262 50080
rect 27946 50015 28262 50016
rect 37946 50080 38262 50081
rect 37946 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38262 50080
rect 37946 50015 38262 50016
rect 47946 50080 48262 50081
rect 47946 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48262 50080
rect 47946 50015 48262 50016
rect 0 49738 800 49768
rect 1301 49738 1367 49741
rect 0 49736 1367 49738
rect 0 49680 1306 49736
rect 1362 49680 1367 49736
rect 0 49678 1367 49680
rect 0 49648 800 49678
rect 1301 49675 1367 49678
rect 49325 49738 49391 49741
rect 50200 49738 51000 49768
rect 49325 49736 51000 49738
rect 49325 49680 49330 49736
rect 49386 49680 51000 49736
rect 49325 49678 51000 49680
rect 49325 49675 49391 49678
rect 50200 49648 51000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 32946 49536 33262 49537
rect 32946 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33262 49536
rect 32946 49471 33262 49472
rect 42946 49536 43262 49537
rect 42946 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43262 49536
rect 42946 49471 43262 49472
rect 7946 48992 8262 48993
rect 0 48922 800 48952
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 27946 48992 28262 48993
rect 27946 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28262 48992
rect 27946 48927 28262 48928
rect 37946 48992 38262 48993
rect 37946 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38262 48992
rect 37946 48927 38262 48928
rect 47946 48992 48262 48993
rect 47946 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48262 48992
rect 47946 48927 48262 48928
rect 1301 48922 1367 48925
rect 0 48920 1367 48922
rect 0 48864 1306 48920
rect 1362 48864 1367 48920
rect 0 48862 1367 48864
rect 0 48832 800 48862
rect 1301 48859 1367 48862
rect 49049 48922 49115 48925
rect 50200 48922 51000 48952
rect 49049 48920 51000 48922
rect 49049 48864 49054 48920
rect 49110 48864 51000 48920
rect 49049 48862 51000 48864
rect 49049 48859 49115 48862
rect 50200 48832 51000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 32946 48448 33262 48449
rect 32946 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33262 48448
rect 32946 48383 33262 48384
rect 42946 48448 43262 48449
rect 42946 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43262 48448
rect 42946 48383 43262 48384
rect 32121 48242 32187 48245
rect 33777 48242 33843 48245
rect 32121 48240 33843 48242
rect 32121 48184 32126 48240
rect 32182 48184 33782 48240
rect 33838 48184 33843 48240
rect 32121 48182 33843 48184
rect 32121 48179 32187 48182
rect 33777 48179 33843 48182
rect 34513 48242 34579 48245
rect 37273 48242 37339 48245
rect 34513 48240 37339 48242
rect 34513 48184 34518 48240
rect 34574 48184 37278 48240
rect 37334 48184 37339 48240
rect 34513 48182 37339 48184
rect 34513 48179 34579 48182
rect 37273 48179 37339 48182
rect 0 48106 800 48136
rect 1301 48106 1367 48109
rect 0 48104 1367 48106
rect 0 48048 1306 48104
rect 1362 48048 1367 48104
rect 0 48046 1367 48048
rect 0 48016 800 48046
rect 1301 48043 1367 48046
rect 32765 48106 32831 48109
rect 36353 48106 36419 48109
rect 32765 48104 36419 48106
rect 32765 48048 32770 48104
rect 32826 48048 36358 48104
rect 36414 48048 36419 48104
rect 32765 48046 36419 48048
rect 32765 48043 32831 48046
rect 36353 48043 36419 48046
rect 36721 48106 36787 48109
rect 37089 48106 37155 48109
rect 36721 48104 37155 48106
rect 36721 48048 36726 48104
rect 36782 48048 37094 48104
rect 37150 48048 37155 48104
rect 36721 48046 37155 48048
rect 36721 48043 36787 48046
rect 37089 48043 37155 48046
rect 49325 48106 49391 48109
rect 50200 48106 51000 48136
rect 49325 48104 51000 48106
rect 49325 48048 49330 48104
rect 49386 48048 51000 48104
rect 49325 48046 51000 48048
rect 49325 48043 49391 48046
rect 50200 48016 51000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 27946 47904 28262 47905
rect 27946 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28262 47904
rect 27946 47839 28262 47840
rect 37946 47904 38262 47905
rect 37946 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38262 47904
rect 37946 47839 38262 47840
rect 47946 47904 48262 47905
rect 47946 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48262 47904
rect 47946 47839 48262 47840
rect 2946 47360 3262 47361
rect 0 47290 800 47320
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 32946 47360 33262 47361
rect 32946 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33262 47360
rect 32946 47295 33262 47296
rect 42946 47360 43262 47361
rect 42946 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43262 47360
rect 42946 47295 43262 47296
rect 1301 47290 1367 47293
rect 0 47288 1367 47290
rect 0 47232 1306 47288
rect 1362 47232 1367 47288
rect 0 47230 1367 47232
rect 0 47200 800 47230
rect 1301 47227 1367 47230
rect 49325 47290 49391 47293
rect 50200 47290 51000 47320
rect 49325 47288 51000 47290
rect 49325 47232 49330 47288
rect 49386 47232 51000 47288
rect 49325 47230 51000 47232
rect 49325 47227 49391 47230
rect 50200 47200 51000 47230
rect 26877 47154 26943 47157
rect 27613 47154 27679 47157
rect 26877 47152 27679 47154
rect 26877 47096 26882 47152
rect 26938 47096 27618 47152
rect 27674 47096 27679 47152
rect 26877 47094 27679 47096
rect 26877 47091 26943 47094
rect 27613 47091 27679 47094
rect 24894 46956 24900 47020
rect 24964 47018 24970 47020
rect 25313 47018 25379 47021
rect 28809 47020 28875 47021
rect 24964 47016 25379 47018
rect 24964 46960 25318 47016
rect 25374 46960 25379 47016
rect 24964 46958 25379 46960
rect 24964 46956 24970 46958
rect 25313 46955 25379 46958
rect 28758 46956 28764 47020
rect 28828 47018 28875 47020
rect 28828 47016 28920 47018
rect 28870 46960 28920 47016
rect 28828 46958 28920 46960
rect 28828 46956 28875 46958
rect 28809 46955 28875 46956
rect 28533 46882 28599 46885
rect 34789 46882 34855 46885
rect 28533 46880 34855 46882
rect 28533 46824 28538 46880
rect 28594 46824 34794 46880
rect 34850 46824 34855 46880
rect 28533 46822 34855 46824
rect 28533 46819 28599 46822
rect 34789 46819 34855 46822
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 27946 46816 28262 46817
rect 27946 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28262 46816
rect 27946 46751 28262 46752
rect 37946 46816 38262 46817
rect 37946 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38262 46816
rect 37946 46751 38262 46752
rect 47946 46816 48262 46817
rect 47946 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48262 46816
rect 47946 46751 48262 46752
rect 26233 46746 26299 46749
rect 27613 46746 27679 46749
rect 26233 46744 27679 46746
rect 26233 46688 26238 46744
rect 26294 46688 27618 46744
rect 27674 46688 27679 46744
rect 26233 46686 27679 46688
rect 26233 46683 26299 46686
rect 27613 46683 27679 46686
rect 0 46474 800 46504
rect 1301 46474 1367 46477
rect 0 46472 1367 46474
rect 0 46416 1306 46472
rect 1362 46416 1367 46472
rect 0 46414 1367 46416
rect 0 46384 800 46414
rect 1301 46411 1367 46414
rect 49049 46474 49115 46477
rect 50200 46474 51000 46504
rect 49049 46472 51000 46474
rect 49049 46416 49054 46472
rect 49110 46416 51000 46472
rect 49049 46414 51000 46416
rect 49049 46411 49115 46414
rect 50200 46384 51000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 32946 46272 33262 46273
rect 32946 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33262 46272
rect 32946 46207 33262 46208
rect 42946 46272 43262 46273
rect 42946 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43262 46272
rect 42946 46207 43262 46208
rect 27337 46066 27403 46069
rect 29269 46066 29335 46069
rect 27337 46064 29335 46066
rect 27337 46008 27342 46064
rect 27398 46008 29274 46064
rect 29330 46008 29335 46064
rect 27337 46006 29335 46008
rect 27337 46003 27403 46006
rect 29269 46003 29335 46006
rect 13629 45930 13695 45933
rect 25262 45930 25268 45932
rect 13629 45928 25268 45930
rect 13629 45872 13634 45928
rect 13690 45872 25268 45928
rect 13629 45870 25268 45872
rect 13629 45867 13695 45870
rect 25262 45868 25268 45870
rect 25332 45930 25338 45932
rect 27889 45930 27955 45933
rect 25332 45928 27955 45930
rect 25332 45872 27894 45928
rect 27950 45872 27955 45928
rect 25332 45870 27955 45872
rect 25332 45868 25338 45870
rect 27889 45867 27955 45870
rect 7946 45728 8262 45729
rect 0 45658 800 45688
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 27946 45728 28262 45729
rect 27946 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28262 45728
rect 27946 45663 28262 45664
rect 37946 45728 38262 45729
rect 37946 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38262 45728
rect 37946 45663 38262 45664
rect 47946 45728 48262 45729
rect 47946 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48262 45728
rect 47946 45663 48262 45664
rect 1301 45658 1367 45661
rect 0 45656 1367 45658
rect 0 45600 1306 45656
rect 1362 45600 1367 45656
rect 0 45598 1367 45600
rect 0 45568 800 45598
rect 1301 45595 1367 45598
rect 49049 45658 49115 45661
rect 50200 45658 51000 45688
rect 49049 45656 51000 45658
rect 49049 45600 49054 45656
rect 49110 45600 51000 45656
rect 49049 45598 51000 45600
rect 49049 45595 49115 45598
rect 50200 45568 51000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 32946 45184 33262 45185
rect 32946 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33262 45184
rect 32946 45119 33262 45120
rect 42946 45184 43262 45185
rect 42946 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43262 45184
rect 42946 45119 43262 45120
rect 33133 44978 33199 44981
rect 36445 44978 36511 44981
rect 33133 44976 36511 44978
rect 33133 44920 33138 44976
rect 33194 44920 36450 44976
rect 36506 44920 36511 44976
rect 33133 44918 36511 44920
rect 33133 44915 33199 44918
rect 36445 44915 36511 44918
rect 0 44842 800 44872
rect 1301 44842 1367 44845
rect 0 44840 1367 44842
rect 0 44784 1306 44840
rect 1362 44784 1367 44840
rect 0 44782 1367 44784
rect 0 44752 800 44782
rect 1301 44779 1367 44782
rect 49049 44842 49115 44845
rect 50200 44842 51000 44872
rect 49049 44840 51000 44842
rect 49049 44784 49054 44840
rect 49110 44784 51000 44840
rect 49049 44782 51000 44784
rect 49049 44779 49115 44782
rect 50200 44752 51000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 27946 44640 28262 44641
rect 27946 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28262 44640
rect 27946 44575 28262 44576
rect 37946 44640 38262 44641
rect 37946 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38262 44640
rect 37946 44575 38262 44576
rect 47946 44640 48262 44641
rect 47946 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48262 44640
rect 47946 44575 48262 44576
rect 3509 44434 3575 44437
rect 22369 44434 22435 44437
rect 3509 44432 22435 44434
rect 3509 44376 3514 44432
rect 3570 44376 22374 44432
rect 22430 44376 22435 44432
rect 3509 44374 22435 44376
rect 3509 44371 3575 44374
rect 22369 44371 22435 44374
rect 23841 44298 23907 44301
rect 22050 44296 23907 44298
rect 22050 44240 23846 44296
rect 23902 44240 23907 44296
rect 22050 44238 23907 44240
rect 13445 44162 13511 44165
rect 22050 44162 22110 44238
rect 23841 44235 23907 44238
rect 28390 44236 28396 44300
rect 28460 44298 28466 44300
rect 28533 44298 28599 44301
rect 28460 44296 28599 44298
rect 28460 44240 28538 44296
rect 28594 44240 28599 44296
rect 28460 44238 28599 44240
rect 28460 44236 28466 44238
rect 28533 44235 28599 44238
rect 30097 44298 30163 44301
rect 30230 44298 30236 44300
rect 30097 44296 30236 44298
rect 30097 44240 30102 44296
rect 30158 44240 30236 44296
rect 30097 44238 30236 44240
rect 30097 44235 30163 44238
rect 30230 44236 30236 44238
rect 30300 44236 30306 44300
rect 13445 44160 22110 44162
rect 13445 44104 13450 44160
rect 13506 44104 22110 44160
rect 13445 44102 22110 44104
rect 33501 44162 33567 44165
rect 35157 44162 35223 44165
rect 38009 44162 38075 44165
rect 33501 44160 38075 44162
rect 33501 44104 33506 44160
rect 33562 44104 35162 44160
rect 35218 44104 38014 44160
rect 38070 44104 38075 44160
rect 33501 44102 38075 44104
rect 13445 44099 13511 44102
rect 33501 44099 33567 44102
rect 35157 44099 35223 44102
rect 38009 44099 38075 44102
rect 2946 44096 3262 44097
rect 0 44026 800 44056
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 32946 44096 33262 44097
rect 32946 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33262 44096
rect 32946 44031 33262 44032
rect 42946 44096 43262 44097
rect 42946 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43262 44096
rect 42946 44031 43262 44032
rect 2037 44026 2103 44029
rect 0 44024 2103 44026
rect 0 43968 2042 44024
rect 2098 43968 2103 44024
rect 0 43966 2103 43968
rect 0 43936 800 43966
rect 2037 43963 2103 43966
rect 49325 44026 49391 44029
rect 50200 44026 51000 44056
rect 49325 44024 51000 44026
rect 49325 43968 49330 44024
rect 49386 43968 51000 44024
rect 49325 43966 51000 43968
rect 49325 43963 49391 43966
rect 50200 43936 51000 43966
rect 34881 43890 34947 43893
rect 37273 43890 37339 43893
rect 34881 43888 37339 43890
rect 34881 43832 34886 43888
rect 34942 43832 37278 43888
rect 37334 43832 37339 43888
rect 34881 43830 37339 43832
rect 34881 43827 34947 43830
rect 37273 43827 37339 43830
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 27946 43552 28262 43553
rect 27946 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28262 43552
rect 27946 43487 28262 43488
rect 37946 43552 38262 43553
rect 37946 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38262 43552
rect 37946 43487 38262 43488
rect 47946 43552 48262 43553
rect 47946 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48262 43552
rect 47946 43487 48262 43488
rect 31569 43346 31635 43349
rect 37549 43346 37615 43349
rect 31569 43344 37615 43346
rect 31569 43288 31574 43344
rect 31630 43288 37554 43344
rect 37610 43288 37615 43344
rect 31569 43286 37615 43288
rect 31569 43283 31635 43286
rect 37549 43283 37615 43286
rect 0 43210 800 43240
rect 1301 43210 1367 43213
rect 0 43208 1367 43210
rect 0 43152 1306 43208
rect 1362 43152 1367 43208
rect 0 43150 1367 43152
rect 0 43120 800 43150
rect 1301 43147 1367 43150
rect 21909 43210 21975 43213
rect 26693 43210 26759 43213
rect 21909 43208 26759 43210
rect 21909 43152 21914 43208
rect 21970 43152 26698 43208
rect 26754 43152 26759 43208
rect 21909 43150 26759 43152
rect 21909 43147 21975 43150
rect 26693 43147 26759 43150
rect 49141 43210 49207 43213
rect 50200 43210 51000 43240
rect 49141 43208 51000 43210
rect 49141 43152 49146 43208
rect 49202 43152 51000 43208
rect 49141 43150 51000 43152
rect 49141 43147 49207 43150
rect 50200 43120 51000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 32946 43008 33262 43009
rect 32946 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33262 43008
rect 32946 42943 33262 42944
rect 42946 43008 43262 43009
rect 42946 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43262 43008
rect 42946 42943 43262 42944
rect 7946 42464 8262 42465
rect 0 42394 800 42424
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 27946 42464 28262 42465
rect 27946 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28262 42464
rect 27946 42399 28262 42400
rect 37946 42464 38262 42465
rect 37946 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38262 42464
rect 37946 42399 38262 42400
rect 47946 42464 48262 42465
rect 47946 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48262 42464
rect 47946 42399 48262 42400
rect 1301 42394 1367 42397
rect 0 42392 1367 42394
rect 0 42336 1306 42392
rect 1362 42336 1367 42392
rect 0 42334 1367 42336
rect 0 42304 800 42334
rect 1301 42331 1367 42334
rect 31201 42394 31267 42397
rect 36261 42394 36327 42397
rect 31201 42392 36327 42394
rect 31201 42336 31206 42392
rect 31262 42336 36266 42392
rect 36322 42336 36327 42392
rect 31201 42334 36327 42336
rect 31201 42331 31267 42334
rect 36261 42331 36327 42334
rect 49049 42394 49115 42397
rect 50200 42394 51000 42424
rect 49049 42392 51000 42394
rect 49049 42336 49054 42392
rect 49110 42336 51000 42392
rect 49049 42334 51000 42336
rect 49049 42331 49115 42334
rect 50200 42304 51000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 32946 41920 33262 41921
rect 32946 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33262 41920
rect 32946 41855 33262 41856
rect 42946 41920 43262 41921
rect 42946 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43262 41920
rect 42946 41855 43262 41856
rect 0 41578 800 41608
rect 1301 41578 1367 41581
rect 0 41576 1367 41578
rect 0 41520 1306 41576
rect 1362 41520 1367 41576
rect 0 41518 1367 41520
rect 0 41488 800 41518
rect 1301 41515 1367 41518
rect 20345 41578 20411 41581
rect 26601 41578 26667 41581
rect 20345 41576 26667 41578
rect 20345 41520 20350 41576
rect 20406 41520 26606 41576
rect 26662 41520 26667 41576
rect 20345 41518 26667 41520
rect 20345 41515 20411 41518
rect 26601 41515 26667 41518
rect 49049 41578 49115 41581
rect 50200 41578 51000 41608
rect 49049 41576 51000 41578
rect 49049 41520 49054 41576
rect 49110 41520 51000 41576
rect 49049 41518 51000 41520
rect 49049 41515 49115 41518
rect 50200 41488 51000 41518
rect 20897 41442 20963 41445
rect 21173 41442 21239 41445
rect 20897 41440 21239 41442
rect 20897 41384 20902 41440
rect 20958 41384 21178 41440
rect 21234 41384 21239 41440
rect 20897 41382 21239 41384
rect 20897 41379 20963 41382
rect 21173 41379 21239 41382
rect 24853 41442 24919 41445
rect 25313 41442 25379 41445
rect 24853 41440 25379 41442
rect 24853 41384 24858 41440
rect 24914 41384 25318 41440
rect 25374 41384 25379 41440
rect 24853 41382 25379 41384
rect 24853 41379 24919 41382
rect 25313 41379 25379 41382
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 27946 41376 28262 41377
rect 27946 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28262 41376
rect 27946 41311 28262 41312
rect 37946 41376 38262 41377
rect 37946 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38262 41376
rect 37946 41311 38262 41312
rect 47946 41376 48262 41377
rect 47946 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48262 41376
rect 47946 41311 48262 41312
rect 25221 41308 25287 41309
rect 25221 41306 25268 41308
rect 25176 41304 25268 41306
rect 25176 41248 25226 41304
rect 25176 41246 25268 41248
rect 25221 41244 25268 41246
rect 25332 41244 25338 41308
rect 32121 41306 32187 41309
rect 32489 41306 32555 41309
rect 32121 41304 32555 41306
rect 32121 41248 32126 41304
rect 32182 41248 32494 41304
rect 32550 41248 32555 41304
rect 32121 41246 32555 41248
rect 25221 41243 25287 41244
rect 32121 41243 32187 41246
rect 32489 41243 32555 41246
rect 31201 41034 31267 41037
rect 32489 41034 32555 41037
rect 31201 41032 32555 41034
rect 31201 40976 31206 41032
rect 31262 40976 32494 41032
rect 32550 40976 32555 41032
rect 31201 40974 32555 40976
rect 31201 40971 31267 40974
rect 32489 40971 32555 40974
rect 28625 40898 28691 40901
rect 28901 40898 28967 40901
rect 28625 40896 28967 40898
rect 28625 40840 28630 40896
rect 28686 40840 28906 40896
rect 28962 40840 28967 40896
rect 28625 40838 28967 40840
rect 28625 40835 28691 40838
rect 28901 40835 28967 40838
rect 2946 40832 3262 40833
rect 0 40762 800 40792
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 32946 40832 33262 40833
rect 32946 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33262 40832
rect 32946 40767 33262 40768
rect 42946 40832 43262 40833
rect 42946 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43262 40832
rect 42946 40767 43262 40768
rect 1301 40762 1367 40765
rect 0 40760 1367 40762
rect 0 40704 1306 40760
rect 1362 40704 1367 40760
rect 0 40702 1367 40704
rect 0 40672 800 40702
rect 1301 40699 1367 40702
rect 28533 40760 28599 40765
rect 28533 40704 28538 40760
rect 28594 40704 28599 40760
rect 28533 40699 28599 40704
rect 49325 40762 49391 40765
rect 50200 40762 51000 40792
rect 49325 40760 51000 40762
rect 49325 40704 49330 40760
rect 49386 40704 51000 40760
rect 49325 40702 51000 40704
rect 49325 40699 49391 40702
rect 20069 40626 20135 40629
rect 20437 40626 20503 40629
rect 22553 40626 22619 40629
rect 20069 40624 22619 40626
rect 20069 40568 20074 40624
rect 20130 40568 20442 40624
rect 20498 40568 22558 40624
rect 22614 40568 22619 40624
rect 20069 40566 22619 40568
rect 20069 40563 20135 40566
rect 20437 40563 20503 40566
rect 22553 40563 22619 40566
rect 28536 40493 28596 40699
rect 50200 40672 51000 40702
rect 28993 40626 29059 40629
rect 37641 40626 37707 40629
rect 28993 40624 37707 40626
rect 28993 40568 28998 40624
rect 29054 40568 37646 40624
rect 37702 40568 37707 40624
rect 28993 40566 37707 40568
rect 28993 40563 29059 40566
rect 37641 40563 37707 40566
rect 13629 40490 13695 40493
rect 19149 40490 19215 40493
rect 26233 40490 26299 40493
rect 13629 40488 26299 40490
rect 13629 40432 13634 40488
rect 13690 40432 19154 40488
rect 19210 40432 26238 40488
rect 26294 40432 26299 40488
rect 13629 40430 26299 40432
rect 13629 40427 13695 40430
rect 19149 40427 19215 40430
rect 26233 40427 26299 40430
rect 28533 40488 28599 40493
rect 28533 40432 28538 40488
rect 28594 40432 28599 40488
rect 28533 40427 28599 40432
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 27946 40288 28262 40289
rect 27946 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28262 40288
rect 27946 40223 28262 40224
rect 37946 40288 38262 40289
rect 37946 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38262 40288
rect 37946 40223 38262 40224
rect 47946 40288 48262 40289
rect 47946 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48262 40288
rect 47946 40223 48262 40224
rect 21214 40156 21220 40220
rect 21284 40218 21290 40220
rect 22829 40218 22895 40221
rect 21284 40216 22895 40218
rect 21284 40160 22834 40216
rect 22890 40160 22895 40216
rect 21284 40158 22895 40160
rect 21284 40156 21290 40158
rect 22829 40155 22895 40158
rect 33409 40082 33475 40085
rect 33869 40082 33935 40085
rect 33409 40080 33935 40082
rect 33409 40024 33414 40080
rect 33470 40024 33874 40080
rect 33930 40024 33935 40080
rect 33409 40022 33935 40024
rect 33409 40019 33475 40022
rect 33869 40019 33935 40022
rect 0 39946 800 39976
rect 2037 39946 2103 39949
rect 0 39944 2103 39946
rect 0 39888 2042 39944
rect 2098 39888 2103 39944
rect 0 39886 2103 39888
rect 0 39856 800 39886
rect 2037 39883 2103 39886
rect 18413 39946 18479 39949
rect 18965 39946 19031 39949
rect 24894 39946 24900 39948
rect 18413 39944 24900 39946
rect 18413 39888 18418 39944
rect 18474 39888 18970 39944
rect 19026 39888 24900 39944
rect 18413 39886 24900 39888
rect 18413 39883 18479 39886
rect 18965 39883 19031 39886
rect 24894 39884 24900 39886
rect 24964 39884 24970 39948
rect 27337 39946 27403 39949
rect 39665 39946 39731 39949
rect 27337 39944 39731 39946
rect 27337 39888 27342 39944
rect 27398 39888 39670 39944
rect 39726 39888 39731 39944
rect 27337 39886 39731 39888
rect 27337 39883 27403 39886
rect 39665 39883 39731 39886
rect 49049 39946 49115 39949
rect 50200 39946 51000 39976
rect 49049 39944 51000 39946
rect 49049 39888 49054 39944
rect 49110 39888 51000 39944
rect 49049 39886 51000 39888
rect 49049 39883 49115 39886
rect 50200 39856 51000 39886
rect 26325 39810 26391 39813
rect 29177 39810 29243 39813
rect 32489 39810 32555 39813
rect 26325 39808 29010 39810
rect 26325 39752 26330 39808
rect 26386 39752 29010 39808
rect 26325 39750 29010 39752
rect 26325 39747 26391 39750
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 28950 39677 29010 39750
rect 29177 39808 32555 39810
rect 29177 39752 29182 39808
rect 29238 39752 32494 39808
rect 32550 39752 32555 39808
rect 29177 39750 32555 39752
rect 29177 39747 29243 39750
rect 32489 39747 32555 39750
rect 32946 39744 33262 39745
rect 32946 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33262 39744
rect 32946 39679 33262 39680
rect 42946 39744 43262 39745
rect 42946 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43262 39744
rect 42946 39679 43262 39680
rect 28901 39672 29010 39677
rect 28901 39616 28906 39672
rect 28962 39616 29010 39672
rect 28901 39614 29010 39616
rect 31753 39674 31819 39677
rect 32765 39674 32831 39677
rect 31753 39672 32831 39674
rect 31753 39616 31758 39672
rect 31814 39616 32770 39672
rect 32826 39616 32831 39672
rect 31753 39614 32831 39616
rect 28901 39611 28967 39614
rect 31753 39611 31819 39614
rect 32765 39611 32831 39614
rect 19057 39538 19123 39541
rect 23013 39538 23079 39541
rect 19057 39536 23079 39538
rect 19057 39480 19062 39536
rect 19118 39480 23018 39536
rect 23074 39480 23079 39536
rect 19057 39478 23079 39480
rect 19057 39475 19123 39478
rect 23013 39475 23079 39478
rect 24393 39538 24459 39541
rect 28758 39538 28764 39540
rect 24393 39536 28764 39538
rect 24393 39480 24398 39536
rect 24454 39480 28764 39536
rect 24393 39478 28764 39480
rect 24393 39475 24459 39478
rect 28758 39476 28764 39478
rect 28828 39538 28834 39540
rect 37641 39538 37707 39541
rect 28828 39536 37707 39538
rect 28828 39480 37646 39536
rect 37702 39480 37707 39536
rect 28828 39478 37707 39480
rect 28828 39476 28834 39478
rect 37641 39475 37707 39478
rect 24894 39340 24900 39404
rect 24964 39402 24970 39404
rect 37457 39402 37523 39405
rect 24964 39400 37523 39402
rect 24964 39344 37462 39400
rect 37518 39344 37523 39400
rect 24964 39342 37523 39344
rect 24964 39340 24970 39342
rect 37457 39339 37523 39342
rect 18597 39266 18663 39269
rect 27429 39266 27495 39269
rect 18597 39264 27495 39266
rect 18597 39208 18602 39264
rect 18658 39208 27434 39264
rect 27490 39208 27495 39264
rect 18597 39206 27495 39208
rect 18597 39203 18663 39206
rect 27429 39203 27495 39206
rect 33961 39266 34027 39269
rect 34094 39266 34100 39268
rect 33961 39264 34100 39266
rect 33961 39208 33966 39264
rect 34022 39208 34100 39264
rect 33961 39206 34100 39208
rect 33961 39203 34027 39206
rect 34094 39204 34100 39206
rect 34164 39204 34170 39268
rect 7946 39200 8262 39201
rect 0 39130 800 39160
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 27946 39200 28262 39201
rect 27946 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28262 39200
rect 27946 39135 28262 39136
rect 37946 39200 38262 39201
rect 37946 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38262 39200
rect 37946 39135 38262 39136
rect 47946 39200 48262 39201
rect 47946 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48262 39200
rect 47946 39135 48262 39136
rect 1301 39130 1367 39133
rect 0 39128 1367 39130
rect 0 39072 1306 39128
rect 1362 39072 1367 39128
rect 0 39070 1367 39072
rect 0 39040 800 39070
rect 1301 39067 1367 39070
rect 16113 39130 16179 39133
rect 17769 39130 17835 39133
rect 16113 39128 17835 39130
rect 16113 39072 16118 39128
rect 16174 39072 17774 39128
rect 17830 39072 17835 39128
rect 16113 39070 17835 39072
rect 16113 39067 16179 39070
rect 17769 39067 17835 39070
rect 18413 39130 18479 39133
rect 27337 39130 27403 39133
rect 18413 39128 27403 39130
rect 18413 39072 18418 39128
rect 18474 39072 27342 39128
rect 27398 39072 27403 39128
rect 18413 39070 27403 39072
rect 18413 39067 18479 39070
rect 27337 39067 27403 39070
rect 31937 39130 32003 39133
rect 32213 39130 32279 39133
rect 31937 39128 32279 39130
rect 31937 39072 31942 39128
rect 31998 39072 32218 39128
rect 32274 39072 32279 39128
rect 31937 39070 32279 39072
rect 31937 39067 32003 39070
rect 32213 39067 32279 39070
rect 49141 39130 49207 39133
rect 50200 39130 51000 39160
rect 49141 39128 51000 39130
rect 49141 39072 49146 39128
rect 49202 39072 51000 39128
rect 49141 39070 51000 39072
rect 49141 39067 49207 39070
rect 50200 39040 51000 39070
rect 22737 38994 22803 38997
rect 23381 38994 23447 38997
rect 22737 38992 23447 38994
rect 22737 38936 22742 38992
rect 22798 38936 23386 38992
rect 23442 38936 23447 38992
rect 22737 38934 23447 38936
rect 22737 38931 22803 38934
rect 23381 38931 23447 38934
rect 26182 38932 26188 38996
rect 26252 38994 26258 38996
rect 26325 38994 26391 38997
rect 26252 38992 26391 38994
rect 26252 38936 26330 38992
rect 26386 38936 26391 38992
rect 26252 38934 26391 38936
rect 26252 38932 26258 38934
rect 26325 38931 26391 38934
rect 31201 38994 31267 38997
rect 38101 38994 38167 38997
rect 31201 38992 38167 38994
rect 31201 38936 31206 38992
rect 31262 38936 38106 38992
rect 38162 38936 38167 38992
rect 31201 38934 38167 38936
rect 31201 38931 31267 38934
rect 38101 38931 38167 38934
rect 22921 38858 22987 38861
rect 24577 38858 24643 38861
rect 24710 38858 24716 38860
rect 22050 38856 24716 38858
rect 22050 38800 22926 38856
rect 22982 38800 24582 38856
rect 24638 38800 24716 38856
rect 22050 38798 24716 38800
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 19701 38586 19767 38589
rect 21725 38586 21791 38589
rect 19701 38584 21791 38586
rect 19701 38528 19706 38584
rect 19762 38528 21730 38584
rect 21786 38528 21791 38584
rect 19701 38526 21791 38528
rect 19701 38523 19767 38526
rect 21725 38523 21791 38526
rect 19977 38450 20043 38453
rect 22050 38450 22110 38798
rect 22921 38795 22987 38798
rect 24577 38795 24643 38798
rect 24710 38796 24716 38798
rect 24780 38796 24786 38860
rect 27429 38858 27495 38861
rect 40125 38858 40191 38861
rect 27429 38856 40191 38858
rect 27429 38800 27434 38856
rect 27490 38800 40130 38856
rect 40186 38800 40191 38856
rect 27429 38798 40191 38800
rect 27429 38795 27495 38798
rect 40125 38795 40191 38798
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 32946 38656 33262 38657
rect 32946 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33262 38656
rect 32946 38591 33262 38592
rect 42946 38656 43262 38657
rect 42946 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43262 38656
rect 42946 38591 43262 38592
rect 19977 38448 22110 38450
rect 19977 38392 19982 38448
rect 20038 38392 22110 38448
rect 19977 38390 22110 38392
rect 19977 38387 20043 38390
rect 0 38314 800 38344
rect 1301 38314 1367 38317
rect 0 38312 1367 38314
rect 0 38256 1306 38312
rect 1362 38256 1367 38312
rect 0 38254 1367 38256
rect 0 38224 800 38254
rect 1301 38251 1367 38254
rect 20069 38314 20135 38317
rect 25681 38314 25747 38317
rect 20069 38312 25747 38314
rect 20069 38256 20074 38312
rect 20130 38256 25686 38312
rect 25742 38256 25747 38312
rect 20069 38254 25747 38256
rect 20069 38251 20135 38254
rect 25681 38251 25747 38254
rect 30373 38314 30439 38317
rect 38469 38314 38535 38317
rect 30373 38312 38535 38314
rect 30373 38256 30378 38312
rect 30434 38256 38474 38312
rect 38530 38256 38535 38312
rect 30373 38254 38535 38256
rect 30373 38251 30439 38254
rect 38469 38251 38535 38254
rect 49141 38314 49207 38317
rect 50200 38314 51000 38344
rect 49141 38312 51000 38314
rect 49141 38256 49146 38312
rect 49202 38256 51000 38312
rect 49141 38254 51000 38256
rect 49141 38251 49207 38254
rect 50200 38224 51000 38254
rect 14549 38178 14615 38181
rect 17401 38178 17467 38181
rect 14549 38176 17467 38178
rect 14549 38120 14554 38176
rect 14610 38120 17406 38176
rect 17462 38120 17467 38176
rect 14549 38118 17467 38120
rect 14549 38115 14615 38118
rect 17401 38115 17467 38118
rect 19425 38178 19491 38181
rect 25405 38178 25471 38181
rect 19425 38176 25471 38178
rect 19425 38120 19430 38176
rect 19486 38120 25410 38176
rect 25466 38120 25471 38176
rect 19425 38118 25471 38120
rect 19425 38115 19491 38118
rect 25405 38115 25471 38118
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 27946 38112 28262 38113
rect 27946 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28262 38112
rect 27946 38047 28262 38048
rect 37946 38112 38262 38113
rect 37946 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38262 38112
rect 37946 38047 38262 38048
rect 47946 38112 48262 38113
rect 47946 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48262 38112
rect 47946 38047 48262 38048
rect 23381 37906 23447 37909
rect 24393 37906 24459 37909
rect 23381 37904 24459 37906
rect 23381 37848 23386 37904
rect 23442 37848 24398 37904
rect 24454 37848 24459 37904
rect 23381 37846 24459 37848
rect 23381 37843 23447 37846
rect 24393 37843 24459 37846
rect 24761 37906 24827 37909
rect 25865 37906 25931 37909
rect 36537 37906 36603 37909
rect 24761 37904 36603 37906
rect 24761 37848 24766 37904
rect 24822 37848 25870 37904
rect 25926 37848 36542 37904
rect 36598 37848 36603 37904
rect 24761 37846 36603 37848
rect 24761 37843 24827 37846
rect 25865 37843 25931 37846
rect 36537 37843 36603 37846
rect 16297 37770 16363 37773
rect 27337 37770 27403 37773
rect 16297 37768 27403 37770
rect 16297 37712 16302 37768
rect 16358 37712 27342 37768
rect 27398 37712 27403 37768
rect 16297 37710 27403 37712
rect 16297 37707 16363 37710
rect 27337 37707 27403 37710
rect 28257 37770 28323 37773
rect 28390 37770 28396 37772
rect 28257 37768 28396 37770
rect 28257 37712 28262 37768
rect 28318 37712 28396 37768
rect 28257 37710 28396 37712
rect 28257 37707 28323 37710
rect 28390 37708 28396 37710
rect 28460 37708 28466 37772
rect 2946 37568 3262 37569
rect 0 37498 800 37528
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 32946 37568 33262 37569
rect 32946 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33262 37568
rect 32946 37503 33262 37504
rect 42946 37568 43262 37569
rect 42946 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43262 37568
rect 42946 37503 43262 37504
rect 1301 37498 1367 37501
rect 0 37496 1367 37498
rect 0 37440 1306 37496
rect 1362 37440 1367 37496
rect 0 37438 1367 37440
rect 0 37408 800 37438
rect 1301 37435 1367 37438
rect 49325 37498 49391 37501
rect 50200 37498 51000 37528
rect 49325 37496 51000 37498
rect 49325 37440 49330 37496
rect 49386 37440 51000 37496
rect 49325 37438 51000 37440
rect 49325 37435 49391 37438
rect 50200 37408 51000 37438
rect 30925 37362 30991 37365
rect 34237 37362 34303 37365
rect 35985 37362 36051 37365
rect 30925 37360 36051 37362
rect 30925 37304 30930 37360
rect 30986 37304 34242 37360
rect 34298 37304 35990 37360
rect 36046 37304 36051 37360
rect 30925 37302 36051 37304
rect 30925 37299 30991 37302
rect 34237 37299 34303 37302
rect 35985 37299 36051 37302
rect 17309 37226 17375 37229
rect 18781 37226 18847 37229
rect 31201 37226 31267 37229
rect 17309 37224 18847 37226
rect 17309 37168 17314 37224
rect 17370 37168 18786 37224
rect 18842 37168 18847 37224
rect 17309 37166 18847 37168
rect 17309 37163 17375 37166
rect 18781 37163 18847 37166
rect 19290 37224 31267 37226
rect 19290 37168 31206 37224
rect 31262 37168 31267 37224
rect 19290 37166 31267 37168
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 16757 36818 16823 36821
rect 18873 36818 18939 36821
rect 16757 36816 18939 36818
rect 16757 36760 16762 36816
rect 16818 36760 18878 36816
rect 18934 36760 18939 36816
rect 16757 36758 18939 36760
rect 16757 36755 16823 36758
rect 18873 36755 18939 36758
rect 19057 36818 19123 36821
rect 19290 36818 19350 37166
rect 31201 37163 31267 37166
rect 31753 37090 31819 37093
rect 37641 37090 37707 37093
rect 31753 37088 37707 37090
rect 31753 37032 31758 37088
rect 31814 37032 37646 37088
rect 37702 37032 37707 37088
rect 31753 37030 37707 37032
rect 31753 37027 31819 37030
rect 37641 37027 37707 37030
rect 27946 37024 28262 37025
rect 27946 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28262 37024
rect 27946 36959 28262 36960
rect 37946 37024 38262 37025
rect 37946 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38262 37024
rect 37946 36959 38262 36960
rect 47946 37024 48262 37025
rect 47946 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48262 37024
rect 47946 36959 48262 36960
rect 20253 36954 20319 36957
rect 25221 36954 25287 36957
rect 20253 36952 25287 36954
rect 20253 36896 20258 36952
rect 20314 36896 25226 36952
rect 25282 36896 25287 36952
rect 20253 36894 25287 36896
rect 20253 36891 20319 36894
rect 25221 36891 25287 36894
rect 19057 36816 19350 36818
rect 19057 36760 19062 36816
rect 19118 36760 19350 36816
rect 19057 36758 19350 36760
rect 19057 36755 19123 36758
rect 0 36682 800 36712
rect 1301 36682 1367 36685
rect 0 36680 1367 36682
rect 0 36624 1306 36680
rect 1362 36624 1367 36680
rect 0 36622 1367 36624
rect 0 36592 800 36622
rect 1301 36619 1367 36622
rect 11973 36682 12039 36685
rect 20897 36682 20963 36685
rect 26182 36682 26188 36684
rect 11973 36680 26188 36682
rect 11973 36624 11978 36680
rect 12034 36624 20902 36680
rect 20958 36624 26188 36680
rect 11973 36622 26188 36624
rect 11973 36619 12039 36622
rect 20897 36619 20963 36622
rect 26182 36620 26188 36622
rect 26252 36682 26258 36684
rect 48313 36682 48379 36685
rect 26252 36680 48379 36682
rect 26252 36624 48318 36680
rect 48374 36624 48379 36680
rect 26252 36622 48379 36624
rect 26252 36620 26258 36622
rect 48313 36619 48379 36622
rect 49049 36682 49115 36685
rect 50200 36682 51000 36712
rect 49049 36680 51000 36682
rect 49049 36624 49054 36680
rect 49110 36624 51000 36680
rect 49049 36622 51000 36624
rect 49049 36619 49115 36622
rect 50200 36592 51000 36622
rect 17493 36546 17559 36549
rect 19241 36546 19307 36549
rect 17493 36544 19307 36546
rect 17493 36488 17498 36544
rect 17554 36488 19246 36544
rect 19302 36488 19307 36544
rect 17493 36486 19307 36488
rect 17493 36483 17559 36486
rect 19241 36483 19307 36486
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 32946 36480 33262 36481
rect 32946 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33262 36480
rect 32946 36415 33262 36416
rect 42946 36480 43262 36481
rect 42946 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43262 36480
rect 42946 36415 43262 36416
rect 15101 36410 15167 36413
rect 15929 36410 15995 36413
rect 16941 36410 17007 36413
rect 15101 36408 17007 36410
rect 15101 36352 15106 36408
rect 15162 36352 15934 36408
rect 15990 36352 16946 36408
rect 17002 36352 17007 36408
rect 15101 36350 17007 36352
rect 15101 36347 15167 36350
rect 15929 36347 15995 36350
rect 16941 36347 17007 36350
rect 16849 36274 16915 36277
rect 18689 36274 18755 36277
rect 16849 36272 18755 36274
rect 16849 36216 16854 36272
rect 16910 36216 18694 36272
rect 18750 36216 18755 36272
rect 16849 36214 18755 36216
rect 16849 36211 16915 36214
rect 18689 36211 18755 36214
rect 15101 36138 15167 36141
rect 19609 36138 19675 36141
rect 26049 36138 26115 36141
rect 15101 36136 26115 36138
rect 15101 36080 15106 36136
rect 15162 36080 19614 36136
rect 19670 36080 26054 36136
rect 26110 36080 26115 36136
rect 15101 36078 26115 36080
rect 15101 36075 15167 36078
rect 19609 36075 19675 36078
rect 26049 36075 26115 36078
rect 28165 36138 28231 36141
rect 28625 36138 28691 36141
rect 28165 36136 28691 36138
rect 28165 36080 28170 36136
rect 28226 36080 28630 36136
rect 28686 36080 28691 36136
rect 28165 36078 28691 36080
rect 28165 36075 28231 36078
rect 28625 36075 28691 36078
rect 11053 36002 11119 36005
rect 17309 36002 17375 36005
rect 11053 36000 17375 36002
rect 11053 35944 11058 36000
rect 11114 35944 17314 36000
rect 17370 35944 17375 36000
rect 11053 35942 17375 35944
rect 11053 35939 11119 35942
rect 17309 35939 17375 35942
rect 23841 36002 23907 36005
rect 24393 36002 24459 36005
rect 25497 36002 25563 36005
rect 25681 36002 25747 36005
rect 23841 36000 25747 36002
rect 23841 35944 23846 36000
rect 23902 35944 24398 36000
rect 24454 35944 25502 36000
rect 25558 35944 25686 36000
rect 25742 35944 25747 36000
rect 23841 35942 25747 35944
rect 23841 35939 23907 35942
rect 24393 35939 24459 35942
rect 25497 35939 25563 35942
rect 25681 35939 25747 35942
rect 7946 35936 8262 35937
rect 0 35866 800 35896
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 27946 35936 28262 35937
rect 27946 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28262 35936
rect 27946 35871 28262 35872
rect 37946 35936 38262 35937
rect 37946 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38262 35936
rect 37946 35871 38262 35872
rect 47946 35936 48262 35937
rect 47946 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48262 35936
rect 47946 35871 48262 35872
rect 2773 35866 2839 35869
rect 0 35864 2839 35866
rect 0 35808 2778 35864
rect 2834 35808 2839 35864
rect 0 35806 2839 35808
rect 0 35776 800 35806
rect 2773 35803 2839 35806
rect 48405 35866 48471 35869
rect 50200 35866 51000 35896
rect 48405 35864 51000 35866
rect 48405 35808 48410 35864
rect 48466 35808 51000 35864
rect 48405 35806 51000 35808
rect 48405 35803 48471 35806
rect 50200 35776 51000 35806
rect 14641 35730 14707 35733
rect 14917 35730 14983 35733
rect 16021 35730 16087 35733
rect 14641 35728 16087 35730
rect 14641 35672 14646 35728
rect 14702 35672 14922 35728
rect 14978 35672 16026 35728
rect 16082 35672 16087 35728
rect 14641 35670 16087 35672
rect 14641 35667 14707 35670
rect 14917 35667 14983 35670
rect 16021 35667 16087 35670
rect 19793 35594 19859 35597
rect 23381 35594 23447 35597
rect 19793 35592 23447 35594
rect 19793 35536 19798 35592
rect 19854 35536 23386 35592
rect 23442 35536 23447 35592
rect 19793 35534 23447 35536
rect 19793 35531 19859 35534
rect 23381 35531 23447 35534
rect 23381 35458 23447 35461
rect 26325 35458 26391 35461
rect 23381 35456 26391 35458
rect 23381 35400 23386 35456
rect 23442 35400 26330 35456
rect 26386 35400 26391 35456
rect 23381 35398 26391 35400
rect 23381 35395 23447 35398
rect 26325 35395 26391 35398
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 32946 35392 33262 35393
rect 32946 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33262 35392
rect 32946 35327 33262 35328
rect 42946 35392 43262 35393
rect 42946 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43262 35392
rect 42946 35327 43262 35328
rect 27981 35322 28047 35325
rect 29637 35322 29703 35325
rect 30230 35322 30236 35324
rect 27981 35320 30236 35322
rect 27981 35264 27986 35320
rect 28042 35264 29642 35320
rect 29698 35264 30236 35320
rect 27981 35262 30236 35264
rect 27981 35259 28047 35262
rect 29637 35259 29703 35262
rect 30230 35260 30236 35262
rect 30300 35260 30306 35324
rect 10869 35186 10935 35189
rect 14641 35186 14707 35189
rect 26693 35186 26759 35189
rect 10869 35184 31770 35186
rect 10869 35128 10874 35184
rect 10930 35128 14646 35184
rect 14702 35128 26698 35184
rect 26754 35128 31770 35184
rect 10869 35126 31770 35128
rect 10869 35123 10935 35126
rect 14641 35123 14707 35126
rect 26693 35123 26759 35126
rect 0 35050 800 35080
rect 1301 35050 1367 35053
rect 0 35048 1367 35050
rect 0 34992 1306 35048
rect 1362 34992 1367 35048
rect 0 34990 1367 34992
rect 0 34960 800 34990
rect 1301 34987 1367 34990
rect 18229 35050 18295 35053
rect 18454 35050 18460 35052
rect 18229 35048 18460 35050
rect 18229 34992 18234 35048
rect 18290 34992 18460 35048
rect 18229 34990 18460 34992
rect 18229 34987 18295 34990
rect 18454 34988 18460 34990
rect 18524 34988 18530 35052
rect 27981 35050 28047 35053
rect 22050 35048 28047 35050
rect 22050 34992 27986 35048
rect 28042 34992 28047 35048
rect 22050 34990 28047 34992
rect 31710 35050 31770 35126
rect 48313 35050 48379 35053
rect 31710 35048 48379 35050
rect 31710 34992 48318 35048
rect 48374 34992 48379 35048
rect 31710 34990 48379 34992
rect 18689 34914 18755 34917
rect 22050 34914 22110 34990
rect 27981 34987 28047 34990
rect 48313 34987 48379 34990
rect 49049 35050 49115 35053
rect 50200 35050 51000 35080
rect 49049 35048 51000 35050
rect 49049 34992 49054 35048
rect 49110 34992 51000 35048
rect 49049 34990 51000 34992
rect 49049 34987 49115 34990
rect 50200 34960 51000 34990
rect 18689 34912 22110 34914
rect 18689 34856 18694 34912
rect 18750 34856 22110 34912
rect 18689 34854 22110 34856
rect 18689 34851 18755 34854
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 27946 34848 28262 34849
rect 27946 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28262 34848
rect 27946 34783 28262 34784
rect 37946 34848 38262 34849
rect 37946 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38262 34848
rect 37946 34783 38262 34784
rect 47946 34848 48262 34849
rect 47946 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48262 34848
rect 47946 34783 48262 34784
rect 22686 34716 22692 34780
rect 22756 34778 22762 34780
rect 23381 34778 23447 34781
rect 22756 34776 23447 34778
rect 22756 34720 23386 34776
rect 23442 34720 23447 34776
rect 22756 34718 23447 34720
rect 22756 34716 22762 34718
rect 23381 34715 23447 34718
rect 23197 34642 23263 34645
rect 27337 34642 27403 34645
rect 28809 34642 28875 34645
rect 23197 34640 28875 34642
rect 23197 34584 23202 34640
rect 23258 34584 27342 34640
rect 27398 34584 28814 34640
rect 28870 34584 28875 34640
rect 23197 34582 28875 34584
rect 23197 34579 23263 34582
rect 27337 34579 27403 34582
rect 28809 34579 28875 34582
rect 2946 34304 3262 34305
rect 0 34234 800 34264
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 32946 34304 33262 34305
rect 32946 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33262 34304
rect 32946 34239 33262 34240
rect 42946 34304 43262 34305
rect 42946 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43262 34304
rect 42946 34239 43262 34240
rect 2037 34234 2103 34237
rect 0 34232 2103 34234
rect 0 34176 2042 34232
rect 2098 34176 2103 34232
rect 0 34174 2103 34176
rect 0 34144 800 34174
rect 2037 34171 2103 34174
rect 18229 34234 18295 34237
rect 18965 34234 19031 34237
rect 18229 34232 19031 34234
rect 18229 34176 18234 34232
rect 18290 34176 18970 34232
rect 19026 34176 19031 34232
rect 18229 34174 19031 34176
rect 18229 34171 18295 34174
rect 18965 34171 19031 34174
rect 49325 34234 49391 34237
rect 50200 34234 51000 34264
rect 49325 34232 51000 34234
rect 49325 34176 49330 34232
rect 49386 34176 51000 34232
rect 49325 34174 51000 34176
rect 49325 34171 49391 34174
rect 50200 34144 51000 34174
rect 32397 34098 32463 34101
rect 34145 34098 34211 34101
rect 32397 34096 34211 34098
rect 32397 34040 32402 34096
rect 32458 34040 34150 34096
rect 34206 34040 34211 34096
rect 32397 34038 34211 34040
rect 32397 34035 32463 34038
rect 34145 34035 34211 34038
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 27946 33760 28262 33761
rect 27946 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28262 33760
rect 27946 33695 28262 33696
rect 37946 33760 38262 33761
rect 37946 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38262 33760
rect 37946 33695 38262 33696
rect 47946 33760 48262 33761
rect 47946 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48262 33760
rect 47946 33695 48262 33696
rect 30005 33554 30071 33557
rect 32489 33554 32555 33557
rect 30005 33552 32555 33554
rect 30005 33496 30010 33552
rect 30066 33496 32494 33552
rect 32550 33496 32555 33552
rect 30005 33494 32555 33496
rect 30005 33491 30071 33494
rect 32489 33491 32555 33494
rect 0 33418 800 33448
rect 1301 33418 1367 33421
rect 0 33416 1367 33418
rect 0 33360 1306 33416
rect 1362 33360 1367 33416
rect 0 33358 1367 33360
rect 0 33328 800 33358
rect 1301 33355 1367 33358
rect 49141 33418 49207 33421
rect 50200 33418 51000 33448
rect 49141 33416 51000 33418
rect 49141 33360 49146 33416
rect 49202 33360 51000 33416
rect 49141 33358 51000 33360
rect 49141 33355 49207 33358
rect 50200 33328 51000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 32946 33216 33262 33217
rect 32946 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33262 33216
rect 32946 33151 33262 33152
rect 42946 33216 43262 33217
rect 42946 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43262 33216
rect 42946 33151 43262 33152
rect 22645 33146 22711 33149
rect 22645 33144 22754 33146
rect 22645 33088 22650 33144
rect 22706 33088 22754 33144
rect 22645 33083 22754 33088
rect 22369 33010 22435 33013
rect 22694 33010 22754 33083
rect 22921 33010 22987 33013
rect 22369 33008 22987 33010
rect 22369 32952 22374 33008
rect 22430 32952 22926 33008
rect 22982 32952 22987 33008
rect 22369 32950 22987 32952
rect 22369 32947 22435 32950
rect 22921 32947 22987 32950
rect 30281 32874 30347 32877
rect 31293 32874 31359 32877
rect 30281 32872 31359 32874
rect 30281 32816 30286 32872
rect 30342 32816 31298 32872
rect 31354 32816 31359 32872
rect 30281 32814 31359 32816
rect 30281 32811 30347 32814
rect 31293 32811 31359 32814
rect 7946 32672 8262 32673
rect 0 32602 800 32632
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 27946 32672 28262 32673
rect 27946 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28262 32672
rect 27946 32607 28262 32608
rect 37946 32672 38262 32673
rect 37946 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38262 32672
rect 37946 32607 38262 32608
rect 47946 32672 48262 32673
rect 47946 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48262 32672
rect 47946 32607 48262 32608
rect 1301 32602 1367 32605
rect 0 32600 1367 32602
rect 0 32544 1306 32600
rect 1362 32544 1367 32600
rect 0 32542 1367 32544
rect 0 32512 800 32542
rect 1301 32539 1367 32542
rect 49049 32602 49115 32605
rect 50200 32602 51000 32632
rect 49049 32600 51000 32602
rect 49049 32544 49054 32600
rect 49110 32544 51000 32600
rect 49049 32542 51000 32544
rect 49049 32539 49115 32542
rect 50200 32512 51000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 32946 32128 33262 32129
rect 32946 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33262 32128
rect 32946 32063 33262 32064
rect 42946 32128 43262 32129
rect 42946 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43262 32128
rect 42946 32063 43262 32064
rect 28901 31922 28967 31925
rect 34513 31922 34579 31925
rect 28901 31920 34579 31922
rect 28901 31864 28906 31920
rect 28962 31864 34518 31920
rect 34574 31864 34579 31920
rect 28901 31862 34579 31864
rect 28901 31859 28967 31862
rect 34513 31859 34579 31862
rect 0 31786 800 31816
rect 1301 31786 1367 31789
rect 0 31784 1367 31786
rect 0 31728 1306 31784
rect 1362 31728 1367 31784
rect 0 31726 1367 31728
rect 0 31696 800 31726
rect 1301 31723 1367 31726
rect 20713 31786 20779 31789
rect 21357 31786 21423 31789
rect 20713 31784 21423 31786
rect 20713 31728 20718 31784
rect 20774 31728 21362 31784
rect 21418 31728 21423 31784
rect 20713 31726 21423 31728
rect 20713 31723 20779 31726
rect 21357 31723 21423 31726
rect 49049 31786 49115 31789
rect 50200 31786 51000 31816
rect 49049 31784 51000 31786
rect 49049 31728 49054 31784
rect 49110 31728 51000 31784
rect 49049 31726 51000 31728
rect 49049 31723 49115 31726
rect 50200 31696 51000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 27946 31584 28262 31585
rect 27946 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28262 31584
rect 27946 31519 28262 31520
rect 37946 31584 38262 31585
rect 37946 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38262 31584
rect 37946 31519 38262 31520
rect 47946 31584 48262 31585
rect 47946 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48262 31584
rect 47946 31519 48262 31520
rect 2946 31040 3262 31041
rect 0 30970 800 31000
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 32946 31040 33262 31041
rect 32946 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33262 31040
rect 32946 30975 33262 30976
rect 42946 31040 43262 31041
rect 42946 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43262 31040
rect 42946 30975 43262 30976
rect 1301 30970 1367 30973
rect 0 30968 1367 30970
rect 0 30912 1306 30968
rect 1362 30912 1367 30968
rect 0 30910 1367 30912
rect 0 30880 800 30910
rect 1301 30907 1367 30910
rect 49325 30970 49391 30973
rect 50200 30970 51000 31000
rect 49325 30968 51000 30970
rect 49325 30912 49330 30968
rect 49386 30912 51000 30968
rect 49325 30910 51000 30912
rect 49325 30907 49391 30910
rect 50200 30880 51000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 27946 30496 28262 30497
rect 27946 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28262 30496
rect 27946 30431 28262 30432
rect 37946 30496 38262 30497
rect 37946 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38262 30496
rect 37946 30431 38262 30432
rect 47946 30496 48262 30497
rect 47946 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48262 30496
rect 47946 30431 48262 30432
rect 0 30154 800 30184
rect 1301 30154 1367 30157
rect 0 30152 1367 30154
rect 0 30096 1306 30152
rect 1362 30096 1367 30152
rect 0 30094 1367 30096
rect 0 30064 800 30094
rect 1301 30091 1367 30094
rect 49049 30154 49115 30157
rect 50200 30154 51000 30184
rect 49049 30152 51000 30154
rect 49049 30096 49054 30152
rect 49110 30096 51000 30152
rect 49049 30094 51000 30096
rect 49049 30091 49115 30094
rect 50200 30064 51000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 32946 29952 33262 29953
rect 32946 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33262 29952
rect 32946 29887 33262 29888
rect 42946 29952 43262 29953
rect 42946 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43262 29952
rect 42946 29887 43262 29888
rect 7946 29408 8262 29409
rect 0 29338 800 29368
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 27946 29408 28262 29409
rect 27946 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28262 29408
rect 27946 29343 28262 29344
rect 37946 29408 38262 29409
rect 37946 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38262 29408
rect 37946 29343 38262 29344
rect 47946 29408 48262 29409
rect 47946 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48262 29408
rect 47946 29343 48262 29344
rect 1301 29338 1367 29341
rect 0 29336 1367 29338
rect 0 29280 1306 29336
rect 1362 29280 1367 29336
rect 0 29278 1367 29280
rect 0 29248 800 29278
rect 1301 29275 1367 29278
rect 49141 29338 49207 29341
rect 50200 29338 51000 29368
rect 49141 29336 51000 29338
rect 49141 29280 49146 29336
rect 49202 29280 51000 29336
rect 49141 29278 51000 29280
rect 49141 29275 49207 29278
rect 50200 29248 51000 29278
rect 16021 29202 16087 29205
rect 16297 29202 16363 29205
rect 22093 29202 22159 29205
rect 16021 29200 22159 29202
rect 16021 29144 16026 29200
rect 16082 29144 16302 29200
rect 16358 29144 22098 29200
rect 22154 29144 22159 29200
rect 16021 29142 22159 29144
rect 16021 29139 16087 29142
rect 16297 29139 16363 29142
rect 22093 29139 22159 29142
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 32946 28864 33262 28865
rect 32946 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33262 28864
rect 32946 28799 33262 28800
rect 42946 28864 43262 28865
rect 42946 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43262 28864
rect 42946 28799 43262 28800
rect 0 28522 800 28552
rect 1301 28522 1367 28525
rect 0 28520 1367 28522
rect 0 28464 1306 28520
rect 1362 28464 1367 28520
rect 0 28462 1367 28464
rect 0 28432 800 28462
rect 1301 28459 1367 28462
rect 49049 28522 49115 28525
rect 50200 28522 51000 28552
rect 49049 28520 51000 28522
rect 49049 28464 49054 28520
rect 49110 28464 51000 28520
rect 49049 28462 51000 28464
rect 49049 28459 49115 28462
rect 50200 28432 51000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 27946 28320 28262 28321
rect 27946 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28262 28320
rect 27946 28255 28262 28256
rect 37946 28320 38262 28321
rect 37946 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38262 28320
rect 37946 28255 38262 28256
rect 47946 28320 48262 28321
rect 47946 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48262 28320
rect 47946 28255 48262 28256
rect 2946 27776 3262 27777
rect 0 27706 800 27736
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 32946 27776 33262 27777
rect 32946 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33262 27776
rect 32946 27711 33262 27712
rect 42946 27776 43262 27777
rect 42946 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43262 27776
rect 42946 27711 43262 27712
rect 1301 27706 1367 27709
rect 0 27704 1367 27706
rect 0 27648 1306 27704
rect 1362 27648 1367 27704
rect 0 27646 1367 27648
rect 0 27616 800 27646
rect 1301 27643 1367 27646
rect 49325 27706 49391 27709
rect 50200 27706 51000 27736
rect 49325 27704 51000 27706
rect 49325 27648 49330 27704
rect 49386 27648 51000 27704
rect 49325 27646 51000 27648
rect 49325 27643 49391 27646
rect 50200 27616 51000 27646
rect 16941 27570 17007 27573
rect 18454 27570 18460 27572
rect 16941 27568 18460 27570
rect 16941 27512 16946 27568
rect 17002 27512 18460 27568
rect 16941 27510 18460 27512
rect 16941 27507 17007 27510
rect 18454 27508 18460 27510
rect 18524 27508 18530 27572
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 27946 27232 28262 27233
rect 27946 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28262 27232
rect 27946 27167 28262 27168
rect 37946 27232 38262 27233
rect 37946 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38262 27232
rect 37946 27167 38262 27168
rect 47946 27232 48262 27233
rect 47946 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48262 27232
rect 47946 27167 48262 27168
rect 0 26890 800 26920
rect 933 26890 999 26893
rect 0 26888 999 26890
rect 0 26832 938 26888
rect 994 26832 999 26888
rect 0 26830 999 26832
rect 0 26800 800 26830
rect 933 26827 999 26830
rect 49141 26890 49207 26893
rect 50200 26890 51000 26920
rect 49141 26888 51000 26890
rect 49141 26832 49146 26888
rect 49202 26832 51000 26888
rect 49141 26830 51000 26832
rect 49141 26827 49207 26830
rect 50200 26800 51000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 32946 26688 33262 26689
rect 32946 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33262 26688
rect 32946 26623 33262 26624
rect 42946 26688 43262 26689
rect 42946 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43262 26688
rect 42946 26623 43262 26624
rect 7946 26144 8262 26145
rect 0 26074 800 26104
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 27946 26144 28262 26145
rect 27946 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28262 26144
rect 27946 26079 28262 26080
rect 37946 26144 38262 26145
rect 37946 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38262 26144
rect 37946 26079 38262 26080
rect 47946 26144 48262 26145
rect 47946 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48262 26144
rect 47946 26079 48262 26080
rect 1669 26074 1735 26077
rect 0 26072 1735 26074
rect 0 26016 1674 26072
rect 1730 26016 1735 26072
rect 0 26014 1735 26016
rect 0 25984 800 26014
rect 1669 26011 1735 26014
rect 48405 26074 48471 26077
rect 50200 26074 51000 26104
rect 48405 26072 51000 26074
rect 48405 26016 48410 26072
rect 48466 26016 51000 26072
rect 48405 26014 51000 26016
rect 48405 26011 48471 26014
rect 50200 25984 51000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 32946 25600 33262 25601
rect 32946 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33262 25600
rect 32946 25535 33262 25536
rect 42946 25600 43262 25601
rect 42946 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43262 25600
rect 42946 25535 43262 25536
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 49141 25258 49207 25261
rect 50200 25258 51000 25288
rect 49141 25256 51000 25258
rect 49141 25200 49146 25256
rect 49202 25200 51000 25256
rect 49141 25198 51000 25200
rect 49141 25195 49207 25198
rect 50200 25168 51000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 27946 25056 28262 25057
rect 27946 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28262 25056
rect 27946 24991 28262 24992
rect 37946 25056 38262 25057
rect 37946 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38262 25056
rect 37946 24991 38262 24992
rect 47946 25056 48262 25057
rect 47946 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48262 25056
rect 47946 24991 48262 24992
rect 33409 24850 33475 24853
rect 34094 24850 34100 24852
rect 33409 24848 34100 24850
rect 33409 24792 33414 24848
rect 33470 24792 34100 24848
rect 33409 24790 34100 24792
rect 33409 24787 33475 24790
rect 34094 24788 34100 24790
rect 34164 24788 34170 24852
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 933 24442 999 24445
rect 0 24440 999 24442
rect 0 24384 938 24440
rect 994 24384 999 24440
rect 0 24382 999 24384
rect 0 24352 800 24382
rect 933 24379 999 24382
rect 49141 24442 49207 24445
rect 50200 24442 51000 24472
rect 49141 24440 51000 24442
rect 49141 24384 49146 24440
rect 49202 24384 51000 24440
rect 49141 24382 51000 24384
rect 49141 24379 49207 24382
rect 50200 24352 51000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 0 23626 800 23656
rect 933 23626 999 23629
rect 0 23624 999 23626
rect 0 23568 938 23624
rect 994 23568 999 23624
rect 0 23566 999 23568
rect 0 23536 800 23566
rect 933 23563 999 23566
rect 49141 23626 49207 23629
rect 50200 23626 51000 23656
rect 49141 23624 51000 23626
rect 49141 23568 49146 23624
rect 49202 23568 51000 23624
rect 49141 23566 51000 23568
rect 49141 23563 49207 23566
rect 50200 23536 51000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 933 22810 999 22813
rect 0 22808 999 22810
rect 0 22752 938 22808
rect 994 22752 999 22808
rect 0 22750 999 22752
rect 0 22720 800 22750
rect 933 22747 999 22750
rect 49141 22810 49207 22813
rect 50200 22810 51000 22840
rect 49141 22808 51000 22810
rect 49141 22752 49146 22808
rect 49202 22752 51000 22808
rect 49141 22750 51000 22752
rect 49141 22747 49207 22750
rect 50200 22720 51000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 0 21994 800 22024
rect 933 21994 999 21997
rect 0 21992 999 21994
rect 0 21936 938 21992
rect 994 21936 999 21992
rect 0 21934 999 21936
rect 0 21904 800 21934
rect 933 21931 999 21934
rect 49141 21994 49207 21997
rect 50200 21994 51000 22024
rect 49141 21992 51000 21994
rect 49141 21936 49146 21992
rect 49202 21936 51000 21992
rect 49141 21934 51000 21936
rect 49141 21931 49207 21934
rect 50200 21904 51000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 49141 21178 49207 21181
rect 50200 21178 51000 21208
rect 49141 21176 51000 21178
rect 49141 21120 49146 21176
rect 49202 21120 51000 21176
rect 49141 21118 51000 21120
rect 49141 21115 49207 21118
rect 50200 21088 51000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 0 20362 800 20392
rect 933 20362 999 20365
rect 0 20360 999 20362
rect 0 20304 938 20360
rect 994 20304 999 20360
rect 0 20302 999 20304
rect 0 20272 800 20302
rect 933 20299 999 20302
rect 49141 20362 49207 20365
rect 50200 20362 51000 20392
rect 49141 20360 51000 20362
rect 49141 20304 49146 20360
rect 49202 20304 51000 20360
rect 49141 20302 51000 20304
rect 49141 20299 49207 20302
rect 50200 20272 51000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 933 19546 999 19549
rect 0 19544 999 19546
rect 0 19488 938 19544
rect 994 19488 999 19544
rect 0 19486 999 19488
rect 0 19456 800 19486
rect 933 19483 999 19486
rect 49141 19546 49207 19549
rect 50200 19546 51000 19576
rect 49141 19544 51000 19546
rect 49141 19488 49146 19544
rect 49202 19488 51000 19544
rect 49141 19486 51000 19488
rect 49141 19483 49207 19486
rect 50200 19456 51000 19486
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 0 18730 800 18760
rect 933 18730 999 18733
rect 0 18728 999 18730
rect 0 18672 938 18728
rect 994 18672 999 18728
rect 0 18670 999 18672
rect 0 18640 800 18670
rect 933 18667 999 18670
rect 49141 18730 49207 18733
rect 50200 18730 51000 18760
rect 49141 18728 51000 18730
rect 49141 18672 49146 18728
rect 49202 18672 51000 18728
rect 49141 18670 51000 18672
rect 49141 18667 49207 18670
rect 50200 18640 51000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 1577 17914 1643 17917
rect 0 17912 1643 17914
rect 0 17856 1582 17912
rect 1638 17856 1643 17912
rect 0 17854 1643 17856
rect 0 17824 800 17854
rect 1577 17851 1643 17854
rect 49141 17914 49207 17917
rect 50200 17914 51000 17944
rect 49141 17912 51000 17914
rect 49141 17856 49146 17912
rect 49202 17856 51000 17912
rect 49141 17854 51000 17856
rect 49141 17851 49207 17854
rect 50200 17824 51000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 2037 17098 2103 17101
rect 22686 17098 22692 17100
rect 2037 17096 22692 17098
rect 2037 17040 2042 17096
rect 2098 17040 22692 17096
rect 2037 17038 22692 17040
rect 2037 17035 2103 17038
rect 22686 17036 22692 17038
rect 22756 17036 22762 17100
rect 49141 17098 49207 17101
rect 50200 17098 51000 17128
rect 49141 17096 51000 17098
rect 49141 17040 49146 17096
rect 49202 17040 51000 17096
rect 49141 17038 51000 17040
rect 49141 17035 49207 17038
rect 50200 17008 51000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 933 16282 999 16285
rect 0 16280 999 16282
rect 0 16224 938 16280
rect 994 16224 999 16280
rect 0 16222 999 16224
rect 0 16192 800 16222
rect 933 16219 999 16222
rect 49141 16282 49207 16285
rect 50200 16282 51000 16312
rect 49141 16280 51000 16282
rect 49141 16224 49146 16280
rect 49202 16224 51000 16280
rect 49141 16222 51000 16224
rect 49141 16219 49207 16222
rect 50200 16192 51000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 0 15466 800 15496
rect 933 15466 999 15469
rect 0 15464 999 15466
rect 0 15408 938 15464
rect 994 15408 999 15464
rect 0 15406 999 15408
rect 0 15376 800 15406
rect 933 15403 999 15406
rect 49141 15466 49207 15469
rect 50200 15466 51000 15496
rect 49141 15464 51000 15466
rect 49141 15408 49146 15464
rect 49202 15408 51000 15464
rect 49141 15406 51000 15408
rect 49141 15403 49207 15406
rect 50200 15376 51000 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 933 14650 999 14653
rect 0 14648 999 14650
rect 0 14592 938 14648
rect 994 14592 999 14648
rect 0 14590 999 14592
rect 0 14560 800 14590
rect 933 14587 999 14590
rect 49141 14650 49207 14653
rect 50200 14650 51000 14680
rect 49141 14648 51000 14650
rect 49141 14592 49146 14648
rect 49202 14592 51000 14648
rect 49141 14590 51000 14592
rect 49141 14587 49207 14590
rect 50200 14560 51000 14590
rect 24710 14316 24716 14380
rect 24780 14378 24786 14380
rect 30373 14378 30439 14381
rect 24780 14376 30439 14378
rect 24780 14320 30378 14376
rect 30434 14320 30439 14376
rect 24780 14318 30439 14320
rect 24780 14316 24786 14318
rect 30373 14315 30439 14318
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 0 13834 800 13864
rect 933 13834 999 13837
rect 0 13832 999 13834
rect 0 13776 938 13832
rect 994 13776 999 13832
rect 0 13774 999 13776
rect 0 13744 800 13774
rect 933 13771 999 13774
rect 49141 13834 49207 13837
rect 50200 13834 51000 13864
rect 49141 13832 51000 13834
rect 49141 13776 49146 13832
rect 49202 13776 51000 13832
rect 49141 13774 51000 13776
rect 49141 13771 49207 13774
rect 50200 13744 51000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 49141 13018 49207 13021
rect 50200 13018 51000 13048
rect 49141 13016 51000 13018
rect 49141 12960 49146 13016
rect 49202 12960 51000 13016
rect 49141 12958 51000 12960
rect 49141 12955 49207 12958
rect 50200 12928 51000 12958
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 0 12202 800 12232
rect 933 12202 999 12205
rect 0 12200 999 12202
rect 0 12144 938 12200
rect 994 12144 999 12200
rect 0 12142 999 12144
rect 0 12112 800 12142
rect 933 12139 999 12142
rect 49141 12202 49207 12205
rect 50200 12202 51000 12232
rect 49141 12200 51000 12202
rect 49141 12144 49146 12200
rect 49202 12144 51000 12200
rect 49141 12142 51000 12144
rect 49141 12139 49207 12142
rect 50200 12112 51000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 933 11386 999 11389
rect 0 11384 999 11386
rect 0 11328 938 11384
rect 994 11328 999 11384
rect 0 11326 999 11328
rect 0 11296 800 11326
rect 933 11323 999 11326
rect 49141 11386 49207 11389
rect 50200 11386 51000 11416
rect 49141 11384 51000 11386
rect 49141 11328 49146 11384
rect 49202 11328 51000 11384
rect 49141 11326 51000 11328
rect 49141 11323 49207 11326
rect 50200 11296 51000 11326
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 0 10570 800 10600
rect 933 10570 999 10573
rect 0 10568 999 10570
rect 0 10512 938 10568
rect 994 10512 999 10568
rect 0 10510 999 10512
rect 0 10480 800 10510
rect 933 10507 999 10510
rect 49141 10570 49207 10573
rect 50200 10570 51000 10600
rect 49141 10568 51000 10570
rect 49141 10512 49146 10568
rect 49202 10512 51000 10568
rect 49141 10510 51000 10512
rect 49141 10507 49207 10510
rect 50200 10480 51000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 933 9754 999 9757
rect 0 9752 999 9754
rect 0 9696 938 9752
rect 994 9696 999 9752
rect 0 9694 999 9696
rect 0 9664 800 9694
rect 933 9691 999 9694
rect 49141 9754 49207 9757
rect 50200 9754 51000 9784
rect 49141 9752 51000 9754
rect 49141 9696 49146 9752
rect 49202 9696 51000 9752
rect 49141 9694 51000 9696
rect 49141 9691 49207 9694
rect 50200 9664 51000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 49141 8938 49207 8941
rect 50200 8938 51000 8968
rect 49141 8936 51000 8938
rect 49141 8880 49146 8936
rect 49202 8880 51000 8936
rect 49141 8878 51000 8880
rect 49141 8875 49207 8878
rect 50200 8848 51000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 800 8062
rect 1577 8059 1643 8062
rect 49141 8122 49207 8125
rect 50200 8122 51000 8152
rect 49141 8120 51000 8122
rect 49141 8064 49146 8120
rect 49202 8064 51000 8120
rect 49141 8062 51000 8064
rect 49141 8059 49207 8062
rect 50200 8032 51000 8062
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 0 7306 800 7336
rect 933 7306 999 7309
rect 0 7304 999 7306
rect 0 7248 938 7304
rect 994 7248 999 7304
rect 0 7246 999 7248
rect 0 7216 800 7246
rect 933 7243 999 7246
rect 49141 7306 49207 7309
rect 50200 7306 51000 7336
rect 49141 7304 51000 7306
rect 49141 7248 49146 7304
rect 49202 7248 51000 7304
rect 49141 7246 51000 7248
rect 49141 7243 49207 7246
rect 50200 7216 51000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 933 6490 999 6493
rect 0 6488 999 6490
rect 0 6432 938 6488
rect 994 6432 999 6488
rect 0 6430 999 6432
rect 0 6400 800 6430
rect 933 6427 999 6430
rect 49141 6490 49207 6493
rect 50200 6490 51000 6520
rect 49141 6488 51000 6490
rect 49141 6432 49146 6488
rect 49202 6432 51000 6488
rect 49141 6430 51000 6432
rect 49141 6427 49207 6430
rect 50200 6400 51000 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 0 5674 800 5704
rect 933 5674 999 5677
rect 0 5672 999 5674
rect 0 5616 938 5672
rect 994 5616 999 5672
rect 0 5614 999 5616
rect 0 5584 800 5614
rect 933 5611 999 5614
rect 49141 5674 49207 5677
rect 50200 5674 51000 5704
rect 49141 5672 51000 5674
rect 49141 5616 49146 5672
rect 49202 5616 51000 5672
rect 49141 5614 51000 5616
rect 49141 5611 49207 5614
rect 50200 5584 51000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 49141 4858 49207 4861
rect 50200 4858 51000 4888
rect 49141 4856 51000 4858
rect 49141 4800 49146 4856
rect 49202 4800 51000 4856
rect 49141 4798 51000 4800
rect 49141 4795 49207 4798
rect 50200 4768 51000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4042 800 4072
rect 933 4042 999 4045
rect 0 4040 999 4042
rect 0 3984 938 4040
rect 994 3984 999 4040
rect 0 3982 999 3984
rect 0 3952 800 3982
rect 933 3979 999 3982
rect 49141 4042 49207 4045
rect 50200 4042 51000 4072
rect 49141 4040 51000 4042
rect 49141 3984 49146 4040
rect 49202 3984 51000 4040
rect 49141 3982 51000 3984
rect 49141 3979 49207 3982
rect 50200 3952 51000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 933 3226 999 3229
rect 0 3224 999 3226
rect 0 3168 938 3224
rect 994 3168 999 3224
rect 0 3166 999 3168
rect 0 3136 800 3166
rect 933 3163 999 3166
rect 49141 3226 49207 3229
rect 50200 3226 51000 3256
rect 49141 3224 51000 3226
rect 49141 3168 49146 3224
rect 49202 3168 51000 3224
rect 49141 3166 51000 3168
rect 49141 3163 49207 3166
rect 50200 3136 51000 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 49141 2410 49207 2413
rect 50200 2410 51000 2440
rect 49141 2408 51000 2410
rect 49141 2352 49146 2408
rect 49202 2352 51000 2408
rect 49141 2350 51000 2352
rect 49141 2347 49207 2350
rect 50200 2320 51000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 27952 54428 28016 54432
rect 27952 54372 27956 54428
rect 27956 54372 28012 54428
rect 28012 54372 28016 54428
rect 27952 54368 28016 54372
rect 28032 54428 28096 54432
rect 28032 54372 28036 54428
rect 28036 54372 28092 54428
rect 28092 54372 28096 54428
rect 28032 54368 28096 54372
rect 28112 54428 28176 54432
rect 28112 54372 28116 54428
rect 28116 54372 28172 54428
rect 28172 54372 28176 54428
rect 28112 54368 28176 54372
rect 28192 54428 28256 54432
rect 28192 54372 28196 54428
rect 28196 54372 28252 54428
rect 28252 54372 28256 54428
rect 28192 54368 28256 54372
rect 37952 54428 38016 54432
rect 37952 54372 37956 54428
rect 37956 54372 38012 54428
rect 38012 54372 38016 54428
rect 37952 54368 38016 54372
rect 38032 54428 38096 54432
rect 38032 54372 38036 54428
rect 38036 54372 38092 54428
rect 38092 54372 38096 54428
rect 38032 54368 38096 54372
rect 38112 54428 38176 54432
rect 38112 54372 38116 54428
rect 38116 54372 38172 54428
rect 38172 54372 38176 54428
rect 38112 54368 38176 54372
rect 38192 54428 38256 54432
rect 38192 54372 38196 54428
rect 38196 54372 38252 54428
rect 38252 54372 38256 54428
rect 38192 54368 38256 54372
rect 47952 54428 48016 54432
rect 47952 54372 47956 54428
rect 47956 54372 48012 54428
rect 48012 54372 48016 54428
rect 47952 54368 48016 54372
rect 48032 54428 48096 54432
rect 48032 54372 48036 54428
rect 48036 54372 48092 54428
rect 48092 54372 48096 54428
rect 48032 54368 48096 54372
rect 48112 54428 48176 54432
rect 48112 54372 48116 54428
rect 48116 54372 48172 54428
rect 48172 54372 48176 54428
rect 48112 54368 48176 54372
rect 48192 54428 48256 54432
rect 48192 54372 48196 54428
rect 48196 54372 48252 54428
rect 48252 54372 48256 54428
rect 48192 54368 48256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 32952 53884 33016 53888
rect 32952 53828 32956 53884
rect 32956 53828 33012 53884
rect 33012 53828 33016 53884
rect 32952 53824 33016 53828
rect 33032 53884 33096 53888
rect 33032 53828 33036 53884
rect 33036 53828 33092 53884
rect 33092 53828 33096 53884
rect 33032 53824 33096 53828
rect 33112 53884 33176 53888
rect 33112 53828 33116 53884
rect 33116 53828 33172 53884
rect 33172 53828 33176 53884
rect 33112 53824 33176 53828
rect 33192 53884 33256 53888
rect 33192 53828 33196 53884
rect 33196 53828 33252 53884
rect 33252 53828 33256 53884
rect 33192 53824 33256 53828
rect 42952 53884 43016 53888
rect 42952 53828 42956 53884
rect 42956 53828 43012 53884
rect 43012 53828 43016 53884
rect 42952 53824 43016 53828
rect 43032 53884 43096 53888
rect 43032 53828 43036 53884
rect 43036 53828 43092 53884
rect 43092 53828 43096 53884
rect 43032 53824 43096 53828
rect 43112 53884 43176 53888
rect 43112 53828 43116 53884
rect 43116 53828 43172 53884
rect 43172 53828 43176 53884
rect 43112 53824 43176 53828
rect 43192 53884 43256 53888
rect 43192 53828 43196 53884
rect 43196 53828 43252 53884
rect 43252 53828 43256 53884
rect 43192 53824 43256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 27952 53340 28016 53344
rect 27952 53284 27956 53340
rect 27956 53284 28012 53340
rect 28012 53284 28016 53340
rect 27952 53280 28016 53284
rect 28032 53340 28096 53344
rect 28032 53284 28036 53340
rect 28036 53284 28092 53340
rect 28092 53284 28096 53340
rect 28032 53280 28096 53284
rect 28112 53340 28176 53344
rect 28112 53284 28116 53340
rect 28116 53284 28172 53340
rect 28172 53284 28176 53340
rect 28112 53280 28176 53284
rect 28192 53340 28256 53344
rect 28192 53284 28196 53340
rect 28196 53284 28252 53340
rect 28252 53284 28256 53340
rect 28192 53280 28256 53284
rect 37952 53340 38016 53344
rect 37952 53284 37956 53340
rect 37956 53284 38012 53340
rect 38012 53284 38016 53340
rect 37952 53280 38016 53284
rect 38032 53340 38096 53344
rect 38032 53284 38036 53340
rect 38036 53284 38092 53340
rect 38092 53284 38096 53340
rect 38032 53280 38096 53284
rect 38112 53340 38176 53344
rect 38112 53284 38116 53340
rect 38116 53284 38172 53340
rect 38172 53284 38176 53340
rect 38112 53280 38176 53284
rect 38192 53340 38256 53344
rect 38192 53284 38196 53340
rect 38196 53284 38252 53340
rect 38252 53284 38256 53340
rect 38192 53280 38256 53284
rect 47952 53340 48016 53344
rect 47952 53284 47956 53340
rect 47956 53284 48012 53340
rect 48012 53284 48016 53340
rect 47952 53280 48016 53284
rect 48032 53340 48096 53344
rect 48032 53284 48036 53340
rect 48036 53284 48092 53340
rect 48092 53284 48096 53340
rect 48032 53280 48096 53284
rect 48112 53340 48176 53344
rect 48112 53284 48116 53340
rect 48116 53284 48172 53340
rect 48172 53284 48176 53340
rect 48112 53280 48176 53284
rect 48192 53340 48256 53344
rect 48192 53284 48196 53340
rect 48196 53284 48252 53340
rect 48252 53284 48256 53340
rect 48192 53280 48256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 32952 52796 33016 52800
rect 32952 52740 32956 52796
rect 32956 52740 33012 52796
rect 33012 52740 33016 52796
rect 32952 52736 33016 52740
rect 33032 52796 33096 52800
rect 33032 52740 33036 52796
rect 33036 52740 33092 52796
rect 33092 52740 33096 52796
rect 33032 52736 33096 52740
rect 33112 52796 33176 52800
rect 33112 52740 33116 52796
rect 33116 52740 33172 52796
rect 33172 52740 33176 52796
rect 33112 52736 33176 52740
rect 33192 52796 33256 52800
rect 33192 52740 33196 52796
rect 33196 52740 33252 52796
rect 33252 52740 33256 52796
rect 33192 52736 33256 52740
rect 42952 52796 43016 52800
rect 42952 52740 42956 52796
rect 42956 52740 43012 52796
rect 43012 52740 43016 52796
rect 42952 52736 43016 52740
rect 43032 52796 43096 52800
rect 43032 52740 43036 52796
rect 43036 52740 43092 52796
rect 43092 52740 43096 52796
rect 43032 52736 43096 52740
rect 43112 52796 43176 52800
rect 43112 52740 43116 52796
rect 43116 52740 43172 52796
rect 43172 52740 43176 52796
rect 43112 52736 43176 52740
rect 43192 52796 43256 52800
rect 43192 52740 43196 52796
rect 43196 52740 43252 52796
rect 43252 52740 43256 52796
rect 43192 52736 43256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 27952 52252 28016 52256
rect 27952 52196 27956 52252
rect 27956 52196 28012 52252
rect 28012 52196 28016 52252
rect 27952 52192 28016 52196
rect 28032 52252 28096 52256
rect 28032 52196 28036 52252
rect 28036 52196 28092 52252
rect 28092 52196 28096 52252
rect 28032 52192 28096 52196
rect 28112 52252 28176 52256
rect 28112 52196 28116 52252
rect 28116 52196 28172 52252
rect 28172 52196 28176 52252
rect 28112 52192 28176 52196
rect 28192 52252 28256 52256
rect 28192 52196 28196 52252
rect 28196 52196 28252 52252
rect 28252 52196 28256 52252
rect 28192 52192 28256 52196
rect 37952 52252 38016 52256
rect 37952 52196 37956 52252
rect 37956 52196 38012 52252
rect 38012 52196 38016 52252
rect 37952 52192 38016 52196
rect 38032 52252 38096 52256
rect 38032 52196 38036 52252
rect 38036 52196 38092 52252
rect 38092 52196 38096 52252
rect 38032 52192 38096 52196
rect 38112 52252 38176 52256
rect 38112 52196 38116 52252
rect 38116 52196 38172 52252
rect 38172 52196 38176 52252
rect 38112 52192 38176 52196
rect 38192 52252 38256 52256
rect 38192 52196 38196 52252
rect 38196 52196 38252 52252
rect 38252 52196 38256 52252
rect 38192 52192 38256 52196
rect 47952 52252 48016 52256
rect 47952 52196 47956 52252
rect 47956 52196 48012 52252
rect 48012 52196 48016 52252
rect 47952 52192 48016 52196
rect 48032 52252 48096 52256
rect 48032 52196 48036 52252
rect 48036 52196 48092 52252
rect 48092 52196 48096 52252
rect 48032 52192 48096 52196
rect 48112 52252 48176 52256
rect 48112 52196 48116 52252
rect 48116 52196 48172 52252
rect 48172 52196 48176 52252
rect 48112 52192 48176 52196
rect 48192 52252 48256 52256
rect 48192 52196 48196 52252
rect 48196 52196 48252 52252
rect 48252 52196 48256 52252
rect 48192 52192 48256 52196
rect 21220 51988 21284 52052
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 32952 51708 33016 51712
rect 32952 51652 32956 51708
rect 32956 51652 33012 51708
rect 33012 51652 33016 51708
rect 32952 51648 33016 51652
rect 33032 51708 33096 51712
rect 33032 51652 33036 51708
rect 33036 51652 33092 51708
rect 33092 51652 33096 51708
rect 33032 51648 33096 51652
rect 33112 51708 33176 51712
rect 33112 51652 33116 51708
rect 33116 51652 33172 51708
rect 33172 51652 33176 51708
rect 33112 51648 33176 51652
rect 33192 51708 33256 51712
rect 33192 51652 33196 51708
rect 33196 51652 33252 51708
rect 33252 51652 33256 51708
rect 33192 51648 33256 51652
rect 42952 51708 43016 51712
rect 42952 51652 42956 51708
rect 42956 51652 43012 51708
rect 43012 51652 43016 51708
rect 42952 51648 43016 51652
rect 43032 51708 43096 51712
rect 43032 51652 43036 51708
rect 43036 51652 43092 51708
rect 43092 51652 43096 51708
rect 43032 51648 43096 51652
rect 43112 51708 43176 51712
rect 43112 51652 43116 51708
rect 43116 51652 43172 51708
rect 43172 51652 43176 51708
rect 43112 51648 43176 51652
rect 43192 51708 43256 51712
rect 43192 51652 43196 51708
rect 43196 51652 43252 51708
rect 43252 51652 43256 51708
rect 43192 51648 43256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 27952 51164 28016 51168
rect 27952 51108 27956 51164
rect 27956 51108 28012 51164
rect 28012 51108 28016 51164
rect 27952 51104 28016 51108
rect 28032 51164 28096 51168
rect 28032 51108 28036 51164
rect 28036 51108 28092 51164
rect 28092 51108 28096 51164
rect 28032 51104 28096 51108
rect 28112 51164 28176 51168
rect 28112 51108 28116 51164
rect 28116 51108 28172 51164
rect 28172 51108 28176 51164
rect 28112 51104 28176 51108
rect 28192 51164 28256 51168
rect 28192 51108 28196 51164
rect 28196 51108 28252 51164
rect 28252 51108 28256 51164
rect 28192 51104 28256 51108
rect 37952 51164 38016 51168
rect 37952 51108 37956 51164
rect 37956 51108 38012 51164
rect 38012 51108 38016 51164
rect 37952 51104 38016 51108
rect 38032 51164 38096 51168
rect 38032 51108 38036 51164
rect 38036 51108 38092 51164
rect 38092 51108 38096 51164
rect 38032 51104 38096 51108
rect 38112 51164 38176 51168
rect 38112 51108 38116 51164
rect 38116 51108 38172 51164
rect 38172 51108 38176 51164
rect 38112 51104 38176 51108
rect 38192 51164 38256 51168
rect 38192 51108 38196 51164
rect 38196 51108 38252 51164
rect 38252 51108 38256 51164
rect 38192 51104 38256 51108
rect 47952 51164 48016 51168
rect 47952 51108 47956 51164
rect 47956 51108 48012 51164
rect 48012 51108 48016 51164
rect 47952 51104 48016 51108
rect 48032 51164 48096 51168
rect 48032 51108 48036 51164
rect 48036 51108 48092 51164
rect 48092 51108 48096 51164
rect 48032 51104 48096 51108
rect 48112 51164 48176 51168
rect 48112 51108 48116 51164
rect 48116 51108 48172 51164
rect 48172 51108 48176 51164
rect 48112 51104 48176 51108
rect 48192 51164 48256 51168
rect 48192 51108 48196 51164
rect 48196 51108 48252 51164
rect 48252 51108 48256 51164
rect 48192 51104 48256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 32952 50620 33016 50624
rect 32952 50564 32956 50620
rect 32956 50564 33012 50620
rect 33012 50564 33016 50620
rect 32952 50560 33016 50564
rect 33032 50620 33096 50624
rect 33032 50564 33036 50620
rect 33036 50564 33092 50620
rect 33092 50564 33096 50620
rect 33032 50560 33096 50564
rect 33112 50620 33176 50624
rect 33112 50564 33116 50620
rect 33116 50564 33172 50620
rect 33172 50564 33176 50620
rect 33112 50560 33176 50564
rect 33192 50620 33256 50624
rect 33192 50564 33196 50620
rect 33196 50564 33252 50620
rect 33252 50564 33256 50620
rect 33192 50560 33256 50564
rect 42952 50620 43016 50624
rect 42952 50564 42956 50620
rect 42956 50564 43012 50620
rect 43012 50564 43016 50620
rect 42952 50560 43016 50564
rect 43032 50620 43096 50624
rect 43032 50564 43036 50620
rect 43036 50564 43092 50620
rect 43092 50564 43096 50620
rect 43032 50560 43096 50564
rect 43112 50620 43176 50624
rect 43112 50564 43116 50620
rect 43116 50564 43172 50620
rect 43172 50564 43176 50620
rect 43112 50560 43176 50564
rect 43192 50620 43256 50624
rect 43192 50564 43196 50620
rect 43196 50564 43252 50620
rect 43252 50564 43256 50620
rect 43192 50560 43256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 27952 50076 28016 50080
rect 27952 50020 27956 50076
rect 27956 50020 28012 50076
rect 28012 50020 28016 50076
rect 27952 50016 28016 50020
rect 28032 50076 28096 50080
rect 28032 50020 28036 50076
rect 28036 50020 28092 50076
rect 28092 50020 28096 50076
rect 28032 50016 28096 50020
rect 28112 50076 28176 50080
rect 28112 50020 28116 50076
rect 28116 50020 28172 50076
rect 28172 50020 28176 50076
rect 28112 50016 28176 50020
rect 28192 50076 28256 50080
rect 28192 50020 28196 50076
rect 28196 50020 28252 50076
rect 28252 50020 28256 50076
rect 28192 50016 28256 50020
rect 37952 50076 38016 50080
rect 37952 50020 37956 50076
rect 37956 50020 38012 50076
rect 38012 50020 38016 50076
rect 37952 50016 38016 50020
rect 38032 50076 38096 50080
rect 38032 50020 38036 50076
rect 38036 50020 38092 50076
rect 38092 50020 38096 50076
rect 38032 50016 38096 50020
rect 38112 50076 38176 50080
rect 38112 50020 38116 50076
rect 38116 50020 38172 50076
rect 38172 50020 38176 50076
rect 38112 50016 38176 50020
rect 38192 50076 38256 50080
rect 38192 50020 38196 50076
rect 38196 50020 38252 50076
rect 38252 50020 38256 50076
rect 38192 50016 38256 50020
rect 47952 50076 48016 50080
rect 47952 50020 47956 50076
rect 47956 50020 48012 50076
rect 48012 50020 48016 50076
rect 47952 50016 48016 50020
rect 48032 50076 48096 50080
rect 48032 50020 48036 50076
rect 48036 50020 48092 50076
rect 48092 50020 48096 50076
rect 48032 50016 48096 50020
rect 48112 50076 48176 50080
rect 48112 50020 48116 50076
rect 48116 50020 48172 50076
rect 48172 50020 48176 50076
rect 48112 50016 48176 50020
rect 48192 50076 48256 50080
rect 48192 50020 48196 50076
rect 48196 50020 48252 50076
rect 48252 50020 48256 50076
rect 48192 50016 48256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 32952 49532 33016 49536
rect 32952 49476 32956 49532
rect 32956 49476 33012 49532
rect 33012 49476 33016 49532
rect 32952 49472 33016 49476
rect 33032 49532 33096 49536
rect 33032 49476 33036 49532
rect 33036 49476 33092 49532
rect 33092 49476 33096 49532
rect 33032 49472 33096 49476
rect 33112 49532 33176 49536
rect 33112 49476 33116 49532
rect 33116 49476 33172 49532
rect 33172 49476 33176 49532
rect 33112 49472 33176 49476
rect 33192 49532 33256 49536
rect 33192 49476 33196 49532
rect 33196 49476 33252 49532
rect 33252 49476 33256 49532
rect 33192 49472 33256 49476
rect 42952 49532 43016 49536
rect 42952 49476 42956 49532
rect 42956 49476 43012 49532
rect 43012 49476 43016 49532
rect 42952 49472 43016 49476
rect 43032 49532 43096 49536
rect 43032 49476 43036 49532
rect 43036 49476 43092 49532
rect 43092 49476 43096 49532
rect 43032 49472 43096 49476
rect 43112 49532 43176 49536
rect 43112 49476 43116 49532
rect 43116 49476 43172 49532
rect 43172 49476 43176 49532
rect 43112 49472 43176 49476
rect 43192 49532 43256 49536
rect 43192 49476 43196 49532
rect 43196 49476 43252 49532
rect 43252 49476 43256 49532
rect 43192 49472 43256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 27952 48988 28016 48992
rect 27952 48932 27956 48988
rect 27956 48932 28012 48988
rect 28012 48932 28016 48988
rect 27952 48928 28016 48932
rect 28032 48988 28096 48992
rect 28032 48932 28036 48988
rect 28036 48932 28092 48988
rect 28092 48932 28096 48988
rect 28032 48928 28096 48932
rect 28112 48988 28176 48992
rect 28112 48932 28116 48988
rect 28116 48932 28172 48988
rect 28172 48932 28176 48988
rect 28112 48928 28176 48932
rect 28192 48988 28256 48992
rect 28192 48932 28196 48988
rect 28196 48932 28252 48988
rect 28252 48932 28256 48988
rect 28192 48928 28256 48932
rect 37952 48988 38016 48992
rect 37952 48932 37956 48988
rect 37956 48932 38012 48988
rect 38012 48932 38016 48988
rect 37952 48928 38016 48932
rect 38032 48988 38096 48992
rect 38032 48932 38036 48988
rect 38036 48932 38092 48988
rect 38092 48932 38096 48988
rect 38032 48928 38096 48932
rect 38112 48988 38176 48992
rect 38112 48932 38116 48988
rect 38116 48932 38172 48988
rect 38172 48932 38176 48988
rect 38112 48928 38176 48932
rect 38192 48988 38256 48992
rect 38192 48932 38196 48988
rect 38196 48932 38252 48988
rect 38252 48932 38256 48988
rect 38192 48928 38256 48932
rect 47952 48988 48016 48992
rect 47952 48932 47956 48988
rect 47956 48932 48012 48988
rect 48012 48932 48016 48988
rect 47952 48928 48016 48932
rect 48032 48988 48096 48992
rect 48032 48932 48036 48988
rect 48036 48932 48092 48988
rect 48092 48932 48096 48988
rect 48032 48928 48096 48932
rect 48112 48988 48176 48992
rect 48112 48932 48116 48988
rect 48116 48932 48172 48988
rect 48172 48932 48176 48988
rect 48112 48928 48176 48932
rect 48192 48988 48256 48992
rect 48192 48932 48196 48988
rect 48196 48932 48252 48988
rect 48252 48932 48256 48988
rect 48192 48928 48256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 32952 48444 33016 48448
rect 32952 48388 32956 48444
rect 32956 48388 33012 48444
rect 33012 48388 33016 48444
rect 32952 48384 33016 48388
rect 33032 48444 33096 48448
rect 33032 48388 33036 48444
rect 33036 48388 33092 48444
rect 33092 48388 33096 48444
rect 33032 48384 33096 48388
rect 33112 48444 33176 48448
rect 33112 48388 33116 48444
rect 33116 48388 33172 48444
rect 33172 48388 33176 48444
rect 33112 48384 33176 48388
rect 33192 48444 33256 48448
rect 33192 48388 33196 48444
rect 33196 48388 33252 48444
rect 33252 48388 33256 48444
rect 33192 48384 33256 48388
rect 42952 48444 43016 48448
rect 42952 48388 42956 48444
rect 42956 48388 43012 48444
rect 43012 48388 43016 48444
rect 42952 48384 43016 48388
rect 43032 48444 43096 48448
rect 43032 48388 43036 48444
rect 43036 48388 43092 48444
rect 43092 48388 43096 48444
rect 43032 48384 43096 48388
rect 43112 48444 43176 48448
rect 43112 48388 43116 48444
rect 43116 48388 43172 48444
rect 43172 48388 43176 48444
rect 43112 48384 43176 48388
rect 43192 48444 43256 48448
rect 43192 48388 43196 48444
rect 43196 48388 43252 48444
rect 43252 48388 43256 48444
rect 43192 48384 43256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 27952 47900 28016 47904
rect 27952 47844 27956 47900
rect 27956 47844 28012 47900
rect 28012 47844 28016 47900
rect 27952 47840 28016 47844
rect 28032 47900 28096 47904
rect 28032 47844 28036 47900
rect 28036 47844 28092 47900
rect 28092 47844 28096 47900
rect 28032 47840 28096 47844
rect 28112 47900 28176 47904
rect 28112 47844 28116 47900
rect 28116 47844 28172 47900
rect 28172 47844 28176 47900
rect 28112 47840 28176 47844
rect 28192 47900 28256 47904
rect 28192 47844 28196 47900
rect 28196 47844 28252 47900
rect 28252 47844 28256 47900
rect 28192 47840 28256 47844
rect 37952 47900 38016 47904
rect 37952 47844 37956 47900
rect 37956 47844 38012 47900
rect 38012 47844 38016 47900
rect 37952 47840 38016 47844
rect 38032 47900 38096 47904
rect 38032 47844 38036 47900
rect 38036 47844 38092 47900
rect 38092 47844 38096 47900
rect 38032 47840 38096 47844
rect 38112 47900 38176 47904
rect 38112 47844 38116 47900
rect 38116 47844 38172 47900
rect 38172 47844 38176 47900
rect 38112 47840 38176 47844
rect 38192 47900 38256 47904
rect 38192 47844 38196 47900
rect 38196 47844 38252 47900
rect 38252 47844 38256 47900
rect 38192 47840 38256 47844
rect 47952 47900 48016 47904
rect 47952 47844 47956 47900
rect 47956 47844 48012 47900
rect 48012 47844 48016 47900
rect 47952 47840 48016 47844
rect 48032 47900 48096 47904
rect 48032 47844 48036 47900
rect 48036 47844 48092 47900
rect 48092 47844 48096 47900
rect 48032 47840 48096 47844
rect 48112 47900 48176 47904
rect 48112 47844 48116 47900
rect 48116 47844 48172 47900
rect 48172 47844 48176 47900
rect 48112 47840 48176 47844
rect 48192 47900 48256 47904
rect 48192 47844 48196 47900
rect 48196 47844 48252 47900
rect 48252 47844 48256 47900
rect 48192 47840 48256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 32952 47356 33016 47360
rect 32952 47300 32956 47356
rect 32956 47300 33012 47356
rect 33012 47300 33016 47356
rect 32952 47296 33016 47300
rect 33032 47356 33096 47360
rect 33032 47300 33036 47356
rect 33036 47300 33092 47356
rect 33092 47300 33096 47356
rect 33032 47296 33096 47300
rect 33112 47356 33176 47360
rect 33112 47300 33116 47356
rect 33116 47300 33172 47356
rect 33172 47300 33176 47356
rect 33112 47296 33176 47300
rect 33192 47356 33256 47360
rect 33192 47300 33196 47356
rect 33196 47300 33252 47356
rect 33252 47300 33256 47356
rect 33192 47296 33256 47300
rect 42952 47356 43016 47360
rect 42952 47300 42956 47356
rect 42956 47300 43012 47356
rect 43012 47300 43016 47356
rect 42952 47296 43016 47300
rect 43032 47356 43096 47360
rect 43032 47300 43036 47356
rect 43036 47300 43092 47356
rect 43092 47300 43096 47356
rect 43032 47296 43096 47300
rect 43112 47356 43176 47360
rect 43112 47300 43116 47356
rect 43116 47300 43172 47356
rect 43172 47300 43176 47356
rect 43112 47296 43176 47300
rect 43192 47356 43256 47360
rect 43192 47300 43196 47356
rect 43196 47300 43252 47356
rect 43252 47300 43256 47356
rect 43192 47296 43256 47300
rect 24900 46956 24964 47020
rect 28764 47016 28828 47020
rect 28764 46960 28814 47016
rect 28814 46960 28828 47016
rect 28764 46956 28828 46960
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 27952 46812 28016 46816
rect 27952 46756 27956 46812
rect 27956 46756 28012 46812
rect 28012 46756 28016 46812
rect 27952 46752 28016 46756
rect 28032 46812 28096 46816
rect 28032 46756 28036 46812
rect 28036 46756 28092 46812
rect 28092 46756 28096 46812
rect 28032 46752 28096 46756
rect 28112 46812 28176 46816
rect 28112 46756 28116 46812
rect 28116 46756 28172 46812
rect 28172 46756 28176 46812
rect 28112 46752 28176 46756
rect 28192 46812 28256 46816
rect 28192 46756 28196 46812
rect 28196 46756 28252 46812
rect 28252 46756 28256 46812
rect 28192 46752 28256 46756
rect 37952 46812 38016 46816
rect 37952 46756 37956 46812
rect 37956 46756 38012 46812
rect 38012 46756 38016 46812
rect 37952 46752 38016 46756
rect 38032 46812 38096 46816
rect 38032 46756 38036 46812
rect 38036 46756 38092 46812
rect 38092 46756 38096 46812
rect 38032 46752 38096 46756
rect 38112 46812 38176 46816
rect 38112 46756 38116 46812
rect 38116 46756 38172 46812
rect 38172 46756 38176 46812
rect 38112 46752 38176 46756
rect 38192 46812 38256 46816
rect 38192 46756 38196 46812
rect 38196 46756 38252 46812
rect 38252 46756 38256 46812
rect 38192 46752 38256 46756
rect 47952 46812 48016 46816
rect 47952 46756 47956 46812
rect 47956 46756 48012 46812
rect 48012 46756 48016 46812
rect 47952 46752 48016 46756
rect 48032 46812 48096 46816
rect 48032 46756 48036 46812
rect 48036 46756 48092 46812
rect 48092 46756 48096 46812
rect 48032 46752 48096 46756
rect 48112 46812 48176 46816
rect 48112 46756 48116 46812
rect 48116 46756 48172 46812
rect 48172 46756 48176 46812
rect 48112 46752 48176 46756
rect 48192 46812 48256 46816
rect 48192 46756 48196 46812
rect 48196 46756 48252 46812
rect 48252 46756 48256 46812
rect 48192 46752 48256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 32952 46268 33016 46272
rect 32952 46212 32956 46268
rect 32956 46212 33012 46268
rect 33012 46212 33016 46268
rect 32952 46208 33016 46212
rect 33032 46268 33096 46272
rect 33032 46212 33036 46268
rect 33036 46212 33092 46268
rect 33092 46212 33096 46268
rect 33032 46208 33096 46212
rect 33112 46268 33176 46272
rect 33112 46212 33116 46268
rect 33116 46212 33172 46268
rect 33172 46212 33176 46268
rect 33112 46208 33176 46212
rect 33192 46268 33256 46272
rect 33192 46212 33196 46268
rect 33196 46212 33252 46268
rect 33252 46212 33256 46268
rect 33192 46208 33256 46212
rect 42952 46268 43016 46272
rect 42952 46212 42956 46268
rect 42956 46212 43012 46268
rect 43012 46212 43016 46268
rect 42952 46208 43016 46212
rect 43032 46268 43096 46272
rect 43032 46212 43036 46268
rect 43036 46212 43092 46268
rect 43092 46212 43096 46268
rect 43032 46208 43096 46212
rect 43112 46268 43176 46272
rect 43112 46212 43116 46268
rect 43116 46212 43172 46268
rect 43172 46212 43176 46268
rect 43112 46208 43176 46212
rect 43192 46268 43256 46272
rect 43192 46212 43196 46268
rect 43196 46212 43252 46268
rect 43252 46212 43256 46268
rect 43192 46208 43256 46212
rect 25268 45868 25332 45932
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 27952 45724 28016 45728
rect 27952 45668 27956 45724
rect 27956 45668 28012 45724
rect 28012 45668 28016 45724
rect 27952 45664 28016 45668
rect 28032 45724 28096 45728
rect 28032 45668 28036 45724
rect 28036 45668 28092 45724
rect 28092 45668 28096 45724
rect 28032 45664 28096 45668
rect 28112 45724 28176 45728
rect 28112 45668 28116 45724
rect 28116 45668 28172 45724
rect 28172 45668 28176 45724
rect 28112 45664 28176 45668
rect 28192 45724 28256 45728
rect 28192 45668 28196 45724
rect 28196 45668 28252 45724
rect 28252 45668 28256 45724
rect 28192 45664 28256 45668
rect 37952 45724 38016 45728
rect 37952 45668 37956 45724
rect 37956 45668 38012 45724
rect 38012 45668 38016 45724
rect 37952 45664 38016 45668
rect 38032 45724 38096 45728
rect 38032 45668 38036 45724
rect 38036 45668 38092 45724
rect 38092 45668 38096 45724
rect 38032 45664 38096 45668
rect 38112 45724 38176 45728
rect 38112 45668 38116 45724
rect 38116 45668 38172 45724
rect 38172 45668 38176 45724
rect 38112 45664 38176 45668
rect 38192 45724 38256 45728
rect 38192 45668 38196 45724
rect 38196 45668 38252 45724
rect 38252 45668 38256 45724
rect 38192 45664 38256 45668
rect 47952 45724 48016 45728
rect 47952 45668 47956 45724
rect 47956 45668 48012 45724
rect 48012 45668 48016 45724
rect 47952 45664 48016 45668
rect 48032 45724 48096 45728
rect 48032 45668 48036 45724
rect 48036 45668 48092 45724
rect 48092 45668 48096 45724
rect 48032 45664 48096 45668
rect 48112 45724 48176 45728
rect 48112 45668 48116 45724
rect 48116 45668 48172 45724
rect 48172 45668 48176 45724
rect 48112 45664 48176 45668
rect 48192 45724 48256 45728
rect 48192 45668 48196 45724
rect 48196 45668 48252 45724
rect 48252 45668 48256 45724
rect 48192 45664 48256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 32952 45180 33016 45184
rect 32952 45124 32956 45180
rect 32956 45124 33012 45180
rect 33012 45124 33016 45180
rect 32952 45120 33016 45124
rect 33032 45180 33096 45184
rect 33032 45124 33036 45180
rect 33036 45124 33092 45180
rect 33092 45124 33096 45180
rect 33032 45120 33096 45124
rect 33112 45180 33176 45184
rect 33112 45124 33116 45180
rect 33116 45124 33172 45180
rect 33172 45124 33176 45180
rect 33112 45120 33176 45124
rect 33192 45180 33256 45184
rect 33192 45124 33196 45180
rect 33196 45124 33252 45180
rect 33252 45124 33256 45180
rect 33192 45120 33256 45124
rect 42952 45180 43016 45184
rect 42952 45124 42956 45180
rect 42956 45124 43012 45180
rect 43012 45124 43016 45180
rect 42952 45120 43016 45124
rect 43032 45180 43096 45184
rect 43032 45124 43036 45180
rect 43036 45124 43092 45180
rect 43092 45124 43096 45180
rect 43032 45120 43096 45124
rect 43112 45180 43176 45184
rect 43112 45124 43116 45180
rect 43116 45124 43172 45180
rect 43172 45124 43176 45180
rect 43112 45120 43176 45124
rect 43192 45180 43256 45184
rect 43192 45124 43196 45180
rect 43196 45124 43252 45180
rect 43252 45124 43256 45180
rect 43192 45120 43256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 27952 44636 28016 44640
rect 27952 44580 27956 44636
rect 27956 44580 28012 44636
rect 28012 44580 28016 44636
rect 27952 44576 28016 44580
rect 28032 44636 28096 44640
rect 28032 44580 28036 44636
rect 28036 44580 28092 44636
rect 28092 44580 28096 44636
rect 28032 44576 28096 44580
rect 28112 44636 28176 44640
rect 28112 44580 28116 44636
rect 28116 44580 28172 44636
rect 28172 44580 28176 44636
rect 28112 44576 28176 44580
rect 28192 44636 28256 44640
rect 28192 44580 28196 44636
rect 28196 44580 28252 44636
rect 28252 44580 28256 44636
rect 28192 44576 28256 44580
rect 37952 44636 38016 44640
rect 37952 44580 37956 44636
rect 37956 44580 38012 44636
rect 38012 44580 38016 44636
rect 37952 44576 38016 44580
rect 38032 44636 38096 44640
rect 38032 44580 38036 44636
rect 38036 44580 38092 44636
rect 38092 44580 38096 44636
rect 38032 44576 38096 44580
rect 38112 44636 38176 44640
rect 38112 44580 38116 44636
rect 38116 44580 38172 44636
rect 38172 44580 38176 44636
rect 38112 44576 38176 44580
rect 38192 44636 38256 44640
rect 38192 44580 38196 44636
rect 38196 44580 38252 44636
rect 38252 44580 38256 44636
rect 38192 44576 38256 44580
rect 47952 44636 48016 44640
rect 47952 44580 47956 44636
rect 47956 44580 48012 44636
rect 48012 44580 48016 44636
rect 47952 44576 48016 44580
rect 48032 44636 48096 44640
rect 48032 44580 48036 44636
rect 48036 44580 48092 44636
rect 48092 44580 48096 44636
rect 48032 44576 48096 44580
rect 48112 44636 48176 44640
rect 48112 44580 48116 44636
rect 48116 44580 48172 44636
rect 48172 44580 48176 44636
rect 48112 44576 48176 44580
rect 48192 44636 48256 44640
rect 48192 44580 48196 44636
rect 48196 44580 48252 44636
rect 48252 44580 48256 44636
rect 48192 44576 48256 44580
rect 28396 44236 28460 44300
rect 30236 44236 30300 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 32952 44092 33016 44096
rect 32952 44036 32956 44092
rect 32956 44036 33012 44092
rect 33012 44036 33016 44092
rect 32952 44032 33016 44036
rect 33032 44092 33096 44096
rect 33032 44036 33036 44092
rect 33036 44036 33092 44092
rect 33092 44036 33096 44092
rect 33032 44032 33096 44036
rect 33112 44092 33176 44096
rect 33112 44036 33116 44092
rect 33116 44036 33172 44092
rect 33172 44036 33176 44092
rect 33112 44032 33176 44036
rect 33192 44092 33256 44096
rect 33192 44036 33196 44092
rect 33196 44036 33252 44092
rect 33252 44036 33256 44092
rect 33192 44032 33256 44036
rect 42952 44092 43016 44096
rect 42952 44036 42956 44092
rect 42956 44036 43012 44092
rect 43012 44036 43016 44092
rect 42952 44032 43016 44036
rect 43032 44092 43096 44096
rect 43032 44036 43036 44092
rect 43036 44036 43092 44092
rect 43092 44036 43096 44092
rect 43032 44032 43096 44036
rect 43112 44092 43176 44096
rect 43112 44036 43116 44092
rect 43116 44036 43172 44092
rect 43172 44036 43176 44092
rect 43112 44032 43176 44036
rect 43192 44092 43256 44096
rect 43192 44036 43196 44092
rect 43196 44036 43252 44092
rect 43252 44036 43256 44092
rect 43192 44032 43256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 27952 43548 28016 43552
rect 27952 43492 27956 43548
rect 27956 43492 28012 43548
rect 28012 43492 28016 43548
rect 27952 43488 28016 43492
rect 28032 43548 28096 43552
rect 28032 43492 28036 43548
rect 28036 43492 28092 43548
rect 28092 43492 28096 43548
rect 28032 43488 28096 43492
rect 28112 43548 28176 43552
rect 28112 43492 28116 43548
rect 28116 43492 28172 43548
rect 28172 43492 28176 43548
rect 28112 43488 28176 43492
rect 28192 43548 28256 43552
rect 28192 43492 28196 43548
rect 28196 43492 28252 43548
rect 28252 43492 28256 43548
rect 28192 43488 28256 43492
rect 37952 43548 38016 43552
rect 37952 43492 37956 43548
rect 37956 43492 38012 43548
rect 38012 43492 38016 43548
rect 37952 43488 38016 43492
rect 38032 43548 38096 43552
rect 38032 43492 38036 43548
rect 38036 43492 38092 43548
rect 38092 43492 38096 43548
rect 38032 43488 38096 43492
rect 38112 43548 38176 43552
rect 38112 43492 38116 43548
rect 38116 43492 38172 43548
rect 38172 43492 38176 43548
rect 38112 43488 38176 43492
rect 38192 43548 38256 43552
rect 38192 43492 38196 43548
rect 38196 43492 38252 43548
rect 38252 43492 38256 43548
rect 38192 43488 38256 43492
rect 47952 43548 48016 43552
rect 47952 43492 47956 43548
rect 47956 43492 48012 43548
rect 48012 43492 48016 43548
rect 47952 43488 48016 43492
rect 48032 43548 48096 43552
rect 48032 43492 48036 43548
rect 48036 43492 48092 43548
rect 48092 43492 48096 43548
rect 48032 43488 48096 43492
rect 48112 43548 48176 43552
rect 48112 43492 48116 43548
rect 48116 43492 48172 43548
rect 48172 43492 48176 43548
rect 48112 43488 48176 43492
rect 48192 43548 48256 43552
rect 48192 43492 48196 43548
rect 48196 43492 48252 43548
rect 48252 43492 48256 43548
rect 48192 43488 48256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 32952 43004 33016 43008
rect 32952 42948 32956 43004
rect 32956 42948 33012 43004
rect 33012 42948 33016 43004
rect 32952 42944 33016 42948
rect 33032 43004 33096 43008
rect 33032 42948 33036 43004
rect 33036 42948 33092 43004
rect 33092 42948 33096 43004
rect 33032 42944 33096 42948
rect 33112 43004 33176 43008
rect 33112 42948 33116 43004
rect 33116 42948 33172 43004
rect 33172 42948 33176 43004
rect 33112 42944 33176 42948
rect 33192 43004 33256 43008
rect 33192 42948 33196 43004
rect 33196 42948 33252 43004
rect 33252 42948 33256 43004
rect 33192 42944 33256 42948
rect 42952 43004 43016 43008
rect 42952 42948 42956 43004
rect 42956 42948 43012 43004
rect 43012 42948 43016 43004
rect 42952 42944 43016 42948
rect 43032 43004 43096 43008
rect 43032 42948 43036 43004
rect 43036 42948 43092 43004
rect 43092 42948 43096 43004
rect 43032 42944 43096 42948
rect 43112 43004 43176 43008
rect 43112 42948 43116 43004
rect 43116 42948 43172 43004
rect 43172 42948 43176 43004
rect 43112 42944 43176 42948
rect 43192 43004 43256 43008
rect 43192 42948 43196 43004
rect 43196 42948 43252 43004
rect 43252 42948 43256 43004
rect 43192 42944 43256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 27952 42460 28016 42464
rect 27952 42404 27956 42460
rect 27956 42404 28012 42460
rect 28012 42404 28016 42460
rect 27952 42400 28016 42404
rect 28032 42460 28096 42464
rect 28032 42404 28036 42460
rect 28036 42404 28092 42460
rect 28092 42404 28096 42460
rect 28032 42400 28096 42404
rect 28112 42460 28176 42464
rect 28112 42404 28116 42460
rect 28116 42404 28172 42460
rect 28172 42404 28176 42460
rect 28112 42400 28176 42404
rect 28192 42460 28256 42464
rect 28192 42404 28196 42460
rect 28196 42404 28252 42460
rect 28252 42404 28256 42460
rect 28192 42400 28256 42404
rect 37952 42460 38016 42464
rect 37952 42404 37956 42460
rect 37956 42404 38012 42460
rect 38012 42404 38016 42460
rect 37952 42400 38016 42404
rect 38032 42460 38096 42464
rect 38032 42404 38036 42460
rect 38036 42404 38092 42460
rect 38092 42404 38096 42460
rect 38032 42400 38096 42404
rect 38112 42460 38176 42464
rect 38112 42404 38116 42460
rect 38116 42404 38172 42460
rect 38172 42404 38176 42460
rect 38112 42400 38176 42404
rect 38192 42460 38256 42464
rect 38192 42404 38196 42460
rect 38196 42404 38252 42460
rect 38252 42404 38256 42460
rect 38192 42400 38256 42404
rect 47952 42460 48016 42464
rect 47952 42404 47956 42460
rect 47956 42404 48012 42460
rect 48012 42404 48016 42460
rect 47952 42400 48016 42404
rect 48032 42460 48096 42464
rect 48032 42404 48036 42460
rect 48036 42404 48092 42460
rect 48092 42404 48096 42460
rect 48032 42400 48096 42404
rect 48112 42460 48176 42464
rect 48112 42404 48116 42460
rect 48116 42404 48172 42460
rect 48172 42404 48176 42460
rect 48112 42400 48176 42404
rect 48192 42460 48256 42464
rect 48192 42404 48196 42460
rect 48196 42404 48252 42460
rect 48252 42404 48256 42460
rect 48192 42400 48256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 32952 41916 33016 41920
rect 32952 41860 32956 41916
rect 32956 41860 33012 41916
rect 33012 41860 33016 41916
rect 32952 41856 33016 41860
rect 33032 41916 33096 41920
rect 33032 41860 33036 41916
rect 33036 41860 33092 41916
rect 33092 41860 33096 41916
rect 33032 41856 33096 41860
rect 33112 41916 33176 41920
rect 33112 41860 33116 41916
rect 33116 41860 33172 41916
rect 33172 41860 33176 41916
rect 33112 41856 33176 41860
rect 33192 41916 33256 41920
rect 33192 41860 33196 41916
rect 33196 41860 33252 41916
rect 33252 41860 33256 41916
rect 33192 41856 33256 41860
rect 42952 41916 43016 41920
rect 42952 41860 42956 41916
rect 42956 41860 43012 41916
rect 43012 41860 43016 41916
rect 42952 41856 43016 41860
rect 43032 41916 43096 41920
rect 43032 41860 43036 41916
rect 43036 41860 43092 41916
rect 43092 41860 43096 41916
rect 43032 41856 43096 41860
rect 43112 41916 43176 41920
rect 43112 41860 43116 41916
rect 43116 41860 43172 41916
rect 43172 41860 43176 41916
rect 43112 41856 43176 41860
rect 43192 41916 43256 41920
rect 43192 41860 43196 41916
rect 43196 41860 43252 41916
rect 43252 41860 43256 41916
rect 43192 41856 43256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 27952 41372 28016 41376
rect 27952 41316 27956 41372
rect 27956 41316 28012 41372
rect 28012 41316 28016 41372
rect 27952 41312 28016 41316
rect 28032 41372 28096 41376
rect 28032 41316 28036 41372
rect 28036 41316 28092 41372
rect 28092 41316 28096 41372
rect 28032 41312 28096 41316
rect 28112 41372 28176 41376
rect 28112 41316 28116 41372
rect 28116 41316 28172 41372
rect 28172 41316 28176 41372
rect 28112 41312 28176 41316
rect 28192 41372 28256 41376
rect 28192 41316 28196 41372
rect 28196 41316 28252 41372
rect 28252 41316 28256 41372
rect 28192 41312 28256 41316
rect 37952 41372 38016 41376
rect 37952 41316 37956 41372
rect 37956 41316 38012 41372
rect 38012 41316 38016 41372
rect 37952 41312 38016 41316
rect 38032 41372 38096 41376
rect 38032 41316 38036 41372
rect 38036 41316 38092 41372
rect 38092 41316 38096 41372
rect 38032 41312 38096 41316
rect 38112 41372 38176 41376
rect 38112 41316 38116 41372
rect 38116 41316 38172 41372
rect 38172 41316 38176 41372
rect 38112 41312 38176 41316
rect 38192 41372 38256 41376
rect 38192 41316 38196 41372
rect 38196 41316 38252 41372
rect 38252 41316 38256 41372
rect 38192 41312 38256 41316
rect 47952 41372 48016 41376
rect 47952 41316 47956 41372
rect 47956 41316 48012 41372
rect 48012 41316 48016 41372
rect 47952 41312 48016 41316
rect 48032 41372 48096 41376
rect 48032 41316 48036 41372
rect 48036 41316 48092 41372
rect 48092 41316 48096 41372
rect 48032 41312 48096 41316
rect 48112 41372 48176 41376
rect 48112 41316 48116 41372
rect 48116 41316 48172 41372
rect 48172 41316 48176 41372
rect 48112 41312 48176 41316
rect 48192 41372 48256 41376
rect 48192 41316 48196 41372
rect 48196 41316 48252 41372
rect 48252 41316 48256 41372
rect 48192 41312 48256 41316
rect 25268 41304 25332 41308
rect 25268 41248 25282 41304
rect 25282 41248 25332 41304
rect 25268 41244 25332 41248
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 32952 40828 33016 40832
rect 32952 40772 32956 40828
rect 32956 40772 33012 40828
rect 33012 40772 33016 40828
rect 32952 40768 33016 40772
rect 33032 40828 33096 40832
rect 33032 40772 33036 40828
rect 33036 40772 33092 40828
rect 33092 40772 33096 40828
rect 33032 40768 33096 40772
rect 33112 40828 33176 40832
rect 33112 40772 33116 40828
rect 33116 40772 33172 40828
rect 33172 40772 33176 40828
rect 33112 40768 33176 40772
rect 33192 40828 33256 40832
rect 33192 40772 33196 40828
rect 33196 40772 33252 40828
rect 33252 40772 33256 40828
rect 33192 40768 33256 40772
rect 42952 40828 43016 40832
rect 42952 40772 42956 40828
rect 42956 40772 43012 40828
rect 43012 40772 43016 40828
rect 42952 40768 43016 40772
rect 43032 40828 43096 40832
rect 43032 40772 43036 40828
rect 43036 40772 43092 40828
rect 43092 40772 43096 40828
rect 43032 40768 43096 40772
rect 43112 40828 43176 40832
rect 43112 40772 43116 40828
rect 43116 40772 43172 40828
rect 43172 40772 43176 40828
rect 43112 40768 43176 40772
rect 43192 40828 43256 40832
rect 43192 40772 43196 40828
rect 43196 40772 43252 40828
rect 43252 40772 43256 40828
rect 43192 40768 43256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 27952 40284 28016 40288
rect 27952 40228 27956 40284
rect 27956 40228 28012 40284
rect 28012 40228 28016 40284
rect 27952 40224 28016 40228
rect 28032 40284 28096 40288
rect 28032 40228 28036 40284
rect 28036 40228 28092 40284
rect 28092 40228 28096 40284
rect 28032 40224 28096 40228
rect 28112 40284 28176 40288
rect 28112 40228 28116 40284
rect 28116 40228 28172 40284
rect 28172 40228 28176 40284
rect 28112 40224 28176 40228
rect 28192 40284 28256 40288
rect 28192 40228 28196 40284
rect 28196 40228 28252 40284
rect 28252 40228 28256 40284
rect 28192 40224 28256 40228
rect 37952 40284 38016 40288
rect 37952 40228 37956 40284
rect 37956 40228 38012 40284
rect 38012 40228 38016 40284
rect 37952 40224 38016 40228
rect 38032 40284 38096 40288
rect 38032 40228 38036 40284
rect 38036 40228 38092 40284
rect 38092 40228 38096 40284
rect 38032 40224 38096 40228
rect 38112 40284 38176 40288
rect 38112 40228 38116 40284
rect 38116 40228 38172 40284
rect 38172 40228 38176 40284
rect 38112 40224 38176 40228
rect 38192 40284 38256 40288
rect 38192 40228 38196 40284
rect 38196 40228 38252 40284
rect 38252 40228 38256 40284
rect 38192 40224 38256 40228
rect 47952 40284 48016 40288
rect 47952 40228 47956 40284
rect 47956 40228 48012 40284
rect 48012 40228 48016 40284
rect 47952 40224 48016 40228
rect 48032 40284 48096 40288
rect 48032 40228 48036 40284
rect 48036 40228 48092 40284
rect 48092 40228 48096 40284
rect 48032 40224 48096 40228
rect 48112 40284 48176 40288
rect 48112 40228 48116 40284
rect 48116 40228 48172 40284
rect 48172 40228 48176 40284
rect 48112 40224 48176 40228
rect 48192 40284 48256 40288
rect 48192 40228 48196 40284
rect 48196 40228 48252 40284
rect 48252 40228 48256 40284
rect 48192 40224 48256 40228
rect 21220 40156 21284 40220
rect 24900 39884 24964 39948
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 32952 39740 33016 39744
rect 32952 39684 32956 39740
rect 32956 39684 33012 39740
rect 33012 39684 33016 39740
rect 32952 39680 33016 39684
rect 33032 39740 33096 39744
rect 33032 39684 33036 39740
rect 33036 39684 33092 39740
rect 33092 39684 33096 39740
rect 33032 39680 33096 39684
rect 33112 39740 33176 39744
rect 33112 39684 33116 39740
rect 33116 39684 33172 39740
rect 33172 39684 33176 39740
rect 33112 39680 33176 39684
rect 33192 39740 33256 39744
rect 33192 39684 33196 39740
rect 33196 39684 33252 39740
rect 33252 39684 33256 39740
rect 33192 39680 33256 39684
rect 42952 39740 43016 39744
rect 42952 39684 42956 39740
rect 42956 39684 43012 39740
rect 43012 39684 43016 39740
rect 42952 39680 43016 39684
rect 43032 39740 43096 39744
rect 43032 39684 43036 39740
rect 43036 39684 43092 39740
rect 43092 39684 43096 39740
rect 43032 39680 43096 39684
rect 43112 39740 43176 39744
rect 43112 39684 43116 39740
rect 43116 39684 43172 39740
rect 43172 39684 43176 39740
rect 43112 39680 43176 39684
rect 43192 39740 43256 39744
rect 43192 39684 43196 39740
rect 43196 39684 43252 39740
rect 43252 39684 43256 39740
rect 43192 39680 43256 39684
rect 28764 39476 28828 39540
rect 24900 39340 24964 39404
rect 34100 39204 34164 39268
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 27952 39196 28016 39200
rect 27952 39140 27956 39196
rect 27956 39140 28012 39196
rect 28012 39140 28016 39196
rect 27952 39136 28016 39140
rect 28032 39196 28096 39200
rect 28032 39140 28036 39196
rect 28036 39140 28092 39196
rect 28092 39140 28096 39196
rect 28032 39136 28096 39140
rect 28112 39196 28176 39200
rect 28112 39140 28116 39196
rect 28116 39140 28172 39196
rect 28172 39140 28176 39196
rect 28112 39136 28176 39140
rect 28192 39196 28256 39200
rect 28192 39140 28196 39196
rect 28196 39140 28252 39196
rect 28252 39140 28256 39196
rect 28192 39136 28256 39140
rect 37952 39196 38016 39200
rect 37952 39140 37956 39196
rect 37956 39140 38012 39196
rect 38012 39140 38016 39196
rect 37952 39136 38016 39140
rect 38032 39196 38096 39200
rect 38032 39140 38036 39196
rect 38036 39140 38092 39196
rect 38092 39140 38096 39196
rect 38032 39136 38096 39140
rect 38112 39196 38176 39200
rect 38112 39140 38116 39196
rect 38116 39140 38172 39196
rect 38172 39140 38176 39196
rect 38112 39136 38176 39140
rect 38192 39196 38256 39200
rect 38192 39140 38196 39196
rect 38196 39140 38252 39196
rect 38252 39140 38256 39196
rect 38192 39136 38256 39140
rect 47952 39196 48016 39200
rect 47952 39140 47956 39196
rect 47956 39140 48012 39196
rect 48012 39140 48016 39196
rect 47952 39136 48016 39140
rect 48032 39196 48096 39200
rect 48032 39140 48036 39196
rect 48036 39140 48092 39196
rect 48092 39140 48096 39196
rect 48032 39136 48096 39140
rect 48112 39196 48176 39200
rect 48112 39140 48116 39196
rect 48116 39140 48172 39196
rect 48172 39140 48176 39196
rect 48112 39136 48176 39140
rect 48192 39196 48256 39200
rect 48192 39140 48196 39196
rect 48196 39140 48252 39196
rect 48252 39140 48256 39196
rect 48192 39136 48256 39140
rect 26188 38932 26252 38996
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 24716 38796 24780 38860
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 32952 38652 33016 38656
rect 32952 38596 32956 38652
rect 32956 38596 33012 38652
rect 33012 38596 33016 38652
rect 32952 38592 33016 38596
rect 33032 38652 33096 38656
rect 33032 38596 33036 38652
rect 33036 38596 33092 38652
rect 33092 38596 33096 38652
rect 33032 38592 33096 38596
rect 33112 38652 33176 38656
rect 33112 38596 33116 38652
rect 33116 38596 33172 38652
rect 33172 38596 33176 38652
rect 33112 38592 33176 38596
rect 33192 38652 33256 38656
rect 33192 38596 33196 38652
rect 33196 38596 33252 38652
rect 33252 38596 33256 38652
rect 33192 38592 33256 38596
rect 42952 38652 43016 38656
rect 42952 38596 42956 38652
rect 42956 38596 43012 38652
rect 43012 38596 43016 38652
rect 42952 38592 43016 38596
rect 43032 38652 43096 38656
rect 43032 38596 43036 38652
rect 43036 38596 43092 38652
rect 43092 38596 43096 38652
rect 43032 38592 43096 38596
rect 43112 38652 43176 38656
rect 43112 38596 43116 38652
rect 43116 38596 43172 38652
rect 43172 38596 43176 38652
rect 43112 38592 43176 38596
rect 43192 38652 43256 38656
rect 43192 38596 43196 38652
rect 43196 38596 43252 38652
rect 43252 38596 43256 38652
rect 43192 38592 43256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 27952 38108 28016 38112
rect 27952 38052 27956 38108
rect 27956 38052 28012 38108
rect 28012 38052 28016 38108
rect 27952 38048 28016 38052
rect 28032 38108 28096 38112
rect 28032 38052 28036 38108
rect 28036 38052 28092 38108
rect 28092 38052 28096 38108
rect 28032 38048 28096 38052
rect 28112 38108 28176 38112
rect 28112 38052 28116 38108
rect 28116 38052 28172 38108
rect 28172 38052 28176 38108
rect 28112 38048 28176 38052
rect 28192 38108 28256 38112
rect 28192 38052 28196 38108
rect 28196 38052 28252 38108
rect 28252 38052 28256 38108
rect 28192 38048 28256 38052
rect 37952 38108 38016 38112
rect 37952 38052 37956 38108
rect 37956 38052 38012 38108
rect 38012 38052 38016 38108
rect 37952 38048 38016 38052
rect 38032 38108 38096 38112
rect 38032 38052 38036 38108
rect 38036 38052 38092 38108
rect 38092 38052 38096 38108
rect 38032 38048 38096 38052
rect 38112 38108 38176 38112
rect 38112 38052 38116 38108
rect 38116 38052 38172 38108
rect 38172 38052 38176 38108
rect 38112 38048 38176 38052
rect 38192 38108 38256 38112
rect 38192 38052 38196 38108
rect 38196 38052 38252 38108
rect 38252 38052 38256 38108
rect 38192 38048 38256 38052
rect 47952 38108 48016 38112
rect 47952 38052 47956 38108
rect 47956 38052 48012 38108
rect 48012 38052 48016 38108
rect 47952 38048 48016 38052
rect 48032 38108 48096 38112
rect 48032 38052 48036 38108
rect 48036 38052 48092 38108
rect 48092 38052 48096 38108
rect 48032 38048 48096 38052
rect 48112 38108 48176 38112
rect 48112 38052 48116 38108
rect 48116 38052 48172 38108
rect 48172 38052 48176 38108
rect 48112 38048 48176 38052
rect 48192 38108 48256 38112
rect 48192 38052 48196 38108
rect 48196 38052 48252 38108
rect 48252 38052 48256 38108
rect 48192 38048 48256 38052
rect 28396 37708 28460 37772
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 32952 37564 33016 37568
rect 32952 37508 32956 37564
rect 32956 37508 33012 37564
rect 33012 37508 33016 37564
rect 32952 37504 33016 37508
rect 33032 37564 33096 37568
rect 33032 37508 33036 37564
rect 33036 37508 33092 37564
rect 33092 37508 33096 37564
rect 33032 37504 33096 37508
rect 33112 37564 33176 37568
rect 33112 37508 33116 37564
rect 33116 37508 33172 37564
rect 33172 37508 33176 37564
rect 33112 37504 33176 37508
rect 33192 37564 33256 37568
rect 33192 37508 33196 37564
rect 33196 37508 33252 37564
rect 33252 37508 33256 37564
rect 33192 37504 33256 37508
rect 42952 37564 43016 37568
rect 42952 37508 42956 37564
rect 42956 37508 43012 37564
rect 43012 37508 43016 37564
rect 42952 37504 43016 37508
rect 43032 37564 43096 37568
rect 43032 37508 43036 37564
rect 43036 37508 43092 37564
rect 43092 37508 43096 37564
rect 43032 37504 43096 37508
rect 43112 37564 43176 37568
rect 43112 37508 43116 37564
rect 43116 37508 43172 37564
rect 43172 37508 43176 37564
rect 43112 37504 43176 37508
rect 43192 37564 43256 37568
rect 43192 37508 43196 37564
rect 43196 37508 43252 37564
rect 43252 37508 43256 37564
rect 43192 37504 43256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 27952 37020 28016 37024
rect 27952 36964 27956 37020
rect 27956 36964 28012 37020
rect 28012 36964 28016 37020
rect 27952 36960 28016 36964
rect 28032 37020 28096 37024
rect 28032 36964 28036 37020
rect 28036 36964 28092 37020
rect 28092 36964 28096 37020
rect 28032 36960 28096 36964
rect 28112 37020 28176 37024
rect 28112 36964 28116 37020
rect 28116 36964 28172 37020
rect 28172 36964 28176 37020
rect 28112 36960 28176 36964
rect 28192 37020 28256 37024
rect 28192 36964 28196 37020
rect 28196 36964 28252 37020
rect 28252 36964 28256 37020
rect 28192 36960 28256 36964
rect 37952 37020 38016 37024
rect 37952 36964 37956 37020
rect 37956 36964 38012 37020
rect 38012 36964 38016 37020
rect 37952 36960 38016 36964
rect 38032 37020 38096 37024
rect 38032 36964 38036 37020
rect 38036 36964 38092 37020
rect 38092 36964 38096 37020
rect 38032 36960 38096 36964
rect 38112 37020 38176 37024
rect 38112 36964 38116 37020
rect 38116 36964 38172 37020
rect 38172 36964 38176 37020
rect 38112 36960 38176 36964
rect 38192 37020 38256 37024
rect 38192 36964 38196 37020
rect 38196 36964 38252 37020
rect 38252 36964 38256 37020
rect 38192 36960 38256 36964
rect 47952 37020 48016 37024
rect 47952 36964 47956 37020
rect 47956 36964 48012 37020
rect 48012 36964 48016 37020
rect 47952 36960 48016 36964
rect 48032 37020 48096 37024
rect 48032 36964 48036 37020
rect 48036 36964 48092 37020
rect 48092 36964 48096 37020
rect 48032 36960 48096 36964
rect 48112 37020 48176 37024
rect 48112 36964 48116 37020
rect 48116 36964 48172 37020
rect 48172 36964 48176 37020
rect 48112 36960 48176 36964
rect 48192 37020 48256 37024
rect 48192 36964 48196 37020
rect 48196 36964 48252 37020
rect 48252 36964 48256 37020
rect 48192 36960 48256 36964
rect 26188 36620 26252 36684
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 32952 36476 33016 36480
rect 32952 36420 32956 36476
rect 32956 36420 33012 36476
rect 33012 36420 33016 36476
rect 32952 36416 33016 36420
rect 33032 36476 33096 36480
rect 33032 36420 33036 36476
rect 33036 36420 33092 36476
rect 33092 36420 33096 36476
rect 33032 36416 33096 36420
rect 33112 36476 33176 36480
rect 33112 36420 33116 36476
rect 33116 36420 33172 36476
rect 33172 36420 33176 36476
rect 33112 36416 33176 36420
rect 33192 36476 33256 36480
rect 33192 36420 33196 36476
rect 33196 36420 33252 36476
rect 33252 36420 33256 36476
rect 33192 36416 33256 36420
rect 42952 36476 43016 36480
rect 42952 36420 42956 36476
rect 42956 36420 43012 36476
rect 43012 36420 43016 36476
rect 42952 36416 43016 36420
rect 43032 36476 43096 36480
rect 43032 36420 43036 36476
rect 43036 36420 43092 36476
rect 43092 36420 43096 36476
rect 43032 36416 43096 36420
rect 43112 36476 43176 36480
rect 43112 36420 43116 36476
rect 43116 36420 43172 36476
rect 43172 36420 43176 36476
rect 43112 36416 43176 36420
rect 43192 36476 43256 36480
rect 43192 36420 43196 36476
rect 43196 36420 43252 36476
rect 43252 36420 43256 36476
rect 43192 36416 43256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 27952 35932 28016 35936
rect 27952 35876 27956 35932
rect 27956 35876 28012 35932
rect 28012 35876 28016 35932
rect 27952 35872 28016 35876
rect 28032 35932 28096 35936
rect 28032 35876 28036 35932
rect 28036 35876 28092 35932
rect 28092 35876 28096 35932
rect 28032 35872 28096 35876
rect 28112 35932 28176 35936
rect 28112 35876 28116 35932
rect 28116 35876 28172 35932
rect 28172 35876 28176 35932
rect 28112 35872 28176 35876
rect 28192 35932 28256 35936
rect 28192 35876 28196 35932
rect 28196 35876 28252 35932
rect 28252 35876 28256 35932
rect 28192 35872 28256 35876
rect 37952 35932 38016 35936
rect 37952 35876 37956 35932
rect 37956 35876 38012 35932
rect 38012 35876 38016 35932
rect 37952 35872 38016 35876
rect 38032 35932 38096 35936
rect 38032 35876 38036 35932
rect 38036 35876 38092 35932
rect 38092 35876 38096 35932
rect 38032 35872 38096 35876
rect 38112 35932 38176 35936
rect 38112 35876 38116 35932
rect 38116 35876 38172 35932
rect 38172 35876 38176 35932
rect 38112 35872 38176 35876
rect 38192 35932 38256 35936
rect 38192 35876 38196 35932
rect 38196 35876 38252 35932
rect 38252 35876 38256 35932
rect 38192 35872 38256 35876
rect 47952 35932 48016 35936
rect 47952 35876 47956 35932
rect 47956 35876 48012 35932
rect 48012 35876 48016 35932
rect 47952 35872 48016 35876
rect 48032 35932 48096 35936
rect 48032 35876 48036 35932
rect 48036 35876 48092 35932
rect 48092 35876 48096 35932
rect 48032 35872 48096 35876
rect 48112 35932 48176 35936
rect 48112 35876 48116 35932
rect 48116 35876 48172 35932
rect 48172 35876 48176 35932
rect 48112 35872 48176 35876
rect 48192 35932 48256 35936
rect 48192 35876 48196 35932
rect 48196 35876 48252 35932
rect 48252 35876 48256 35932
rect 48192 35872 48256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 32952 35388 33016 35392
rect 32952 35332 32956 35388
rect 32956 35332 33012 35388
rect 33012 35332 33016 35388
rect 32952 35328 33016 35332
rect 33032 35388 33096 35392
rect 33032 35332 33036 35388
rect 33036 35332 33092 35388
rect 33092 35332 33096 35388
rect 33032 35328 33096 35332
rect 33112 35388 33176 35392
rect 33112 35332 33116 35388
rect 33116 35332 33172 35388
rect 33172 35332 33176 35388
rect 33112 35328 33176 35332
rect 33192 35388 33256 35392
rect 33192 35332 33196 35388
rect 33196 35332 33252 35388
rect 33252 35332 33256 35388
rect 33192 35328 33256 35332
rect 42952 35388 43016 35392
rect 42952 35332 42956 35388
rect 42956 35332 43012 35388
rect 43012 35332 43016 35388
rect 42952 35328 43016 35332
rect 43032 35388 43096 35392
rect 43032 35332 43036 35388
rect 43036 35332 43092 35388
rect 43092 35332 43096 35388
rect 43032 35328 43096 35332
rect 43112 35388 43176 35392
rect 43112 35332 43116 35388
rect 43116 35332 43172 35388
rect 43172 35332 43176 35388
rect 43112 35328 43176 35332
rect 43192 35388 43256 35392
rect 43192 35332 43196 35388
rect 43196 35332 43252 35388
rect 43252 35332 43256 35388
rect 43192 35328 43256 35332
rect 30236 35260 30300 35324
rect 18460 34988 18524 35052
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 27952 34844 28016 34848
rect 27952 34788 27956 34844
rect 27956 34788 28012 34844
rect 28012 34788 28016 34844
rect 27952 34784 28016 34788
rect 28032 34844 28096 34848
rect 28032 34788 28036 34844
rect 28036 34788 28092 34844
rect 28092 34788 28096 34844
rect 28032 34784 28096 34788
rect 28112 34844 28176 34848
rect 28112 34788 28116 34844
rect 28116 34788 28172 34844
rect 28172 34788 28176 34844
rect 28112 34784 28176 34788
rect 28192 34844 28256 34848
rect 28192 34788 28196 34844
rect 28196 34788 28252 34844
rect 28252 34788 28256 34844
rect 28192 34784 28256 34788
rect 37952 34844 38016 34848
rect 37952 34788 37956 34844
rect 37956 34788 38012 34844
rect 38012 34788 38016 34844
rect 37952 34784 38016 34788
rect 38032 34844 38096 34848
rect 38032 34788 38036 34844
rect 38036 34788 38092 34844
rect 38092 34788 38096 34844
rect 38032 34784 38096 34788
rect 38112 34844 38176 34848
rect 38112 34788 38116 34844
rect 38116 34788 38172 34844
rect 38172 34788 38176 34844
rect 38112 34784 38176 34788
rect 38192 34844 38256 34848
rect 38192 34788 38196 34844
rect 38196 34788 38252 34844
rect 38252 34788 38256 34844
rect 38192 34784 38256 34788
rect 47952 34844 48016 34848
rect 47952 34788 47956 34844
rect 47956 34788 48012 34844
rect 48012 34788 48016 34844
rect 47952 34784 48016 34788
rect 48032 34844 48096 34848
rect 48032 34788 48036 34844
rect 48036 34788 48092 34844
rect 48092 34788 48096 34844
rect 48032 34784 48096 34788
rect 48112 34844 48176 34848
rect 48112 34788 48116 34844
rect 48116 34788 48172 34844
rect 48172 34788 48176 34844
rect 48112 34784 48176 34788
rect 48192 34844 48256 34848
rect 48192 34788 48196 34844
rect 48196 34788 48252 34844
rect 48252 34788 48256 34844
rect 48192 34784 48256 34788
rect 22692 34716 22756 34780
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 32952 34300 33016 34304
rect 32952 34244 32956 34300
rect 32956 34244 33012 34300
rect 33012 34244 33016 34300
rect 32952 34240 33016 34244
rect 33032 34300 33096 34304
rect 33032 34244 33036 34300
rect 33036 34244 33092 34300
rect 33092 34244 33096 34300
rect 33032 34240 33096 34244
rect 33112 34300 33176 34304
rect 33112 34244 33116 34300
rect 33116 34244 33172 34300
rect 33172 34244 33176 34300
rect 33112 34240 33176 34244
rect 33192 34300 33256 34304
rect 33192 34244 33196 34300
rect 33196 34244 33252 34300
rect 33252 34244 33256 34300
rect 33192 34240 33256 34244
rect 42952 34300 43016 34304
rect 42952 34244 42956 34300
rect 42956 34244 43012 34300
rect 43012 34244 43016 34300
rect 42952 34240 43016 34244
rect 43032 34300 43096 34304
rect 43032 34244 43036 34300
rect 43036 34244 43092 34300
rect 43092 34244 43096 34300
rect 43032 34240 43096 34244
rect 43112 34300 43176 34304
rect 43112 34244 43116 34300
rect 43116 34244 43172 34300
rect 43172 34244 43176 34300
rect 43112 34240 43176 34244
rect 43192 34300 43256 34304
rect 43192 34244 43196 34300
rect 43196 34244 43252 34300
rect 43252 34244 43256 34300
rect 43192 34240 43256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 27952 33756 28016 33760
rect 27952 33700 27956 33756
rect 27956 33700 28012 33756
rect 28012 33700 28016 33756
rect 27952 33696 28016 33700
rect 28032 33756 28096 33760
rect 28032 33700 28036 33756
rect 28036 33700 28092 33756
rect 28092 33700 28096 33756
rect 28032 33696 28096 33700
rect 28112 33756 28176 33760
rect 28112 33700 28116 33756
rect 28116 33700 28172 33756
rect 28172 33700 28176 33756
rect 28112 33696 28176 33700
rect 28192 33756 28256 33760
rect 28192 33700 28196 33756
rect 28196 33700 28252 33756
rect 28252 33700 28256 33756
rect 28192 33696 28256 33700
rect 37952 33756 38016 33760
rect 37952 33700 37956 33756
rect 37956 33700 38012 33756
rect 38012 33700 38016 33756
rect 37952 33696 38016 33700
rect 38032 33756 38096 33760
rect 38032 33700 38036 33756
rect 38036 33700 38092 33756
rect 38092 33700 38096 33756
rect 38032 33696 38096 33700
rect 38112 33756 38176 33760
rect 38112 33700 38116 33756
rect 38116 33700 38172 33756
rect 38172 33700 38176 33756
rect 38112 33696 38176 33700
rect 38192 33756 38256 33760
rect 38192 33700 38196 33756
rect 38196 33700 38252 33756
rect 38252 33700 38256 33756
rect 38192 33696 38256 33700
rect 47952 33756 48016 33760
rect 47952 33700 47956 33756
rect 47956 33700 48012 33756
rect 48012 33700 48016 33756
rect 47952 33696 48016 33700
rect 48032 33756 48096 33760
rect 48032 33700 48036 33756
rect 48036 33700 48092 33756
rect 48092 33700 48096 33756
rect 48032 33696 48096 33700
rect 48112 33756 48176 33760
rect 48112 33700 48116 33756
rect 48116 33700 48172 33756
rect 48172 33700 48176 33756
rect 48112 33696 48176 33700
rect 48192 33756 48256 33760
rect 48192 33700 48196 33756
rect 48196 33700 48252 33756
rect 48252 33700 48256 33756
rect 48192 33696 48256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 32952 33212 33016 33216
rect 32952 33156 32956 33212
rect 32956 33156 33012 33212
rect 33012 33156 33016 33212
rect 32952 33152 33016 33156
rect 33032 33212 33096 33216
rect 33032 33156 33036 33212
rect 33036 33156 33092 33212
rect 33092 33156 33096 33212
rect 33032 33152 33096 33156
rect 33112 33212 33176 33216
rect 33112 33156 33116 33212
rect 33116 33156 33172 33212
rect 33172 33156 33176 33212
rect 33112 33152 33176 33156
rect 33192 33212 33256 33216
rect 33192 33156 33196 33212
rect 33196 33156 33252 33212
rect 33252 33156 33256 33212
rect 33192 33152 33256 33156
rect 42952 33212 43016 33216
rect 42952 33156 42956 33212
rect 42956 33156 43012 33212
rect 43012 33156 43016 33212
rect 42952 33152 43016 33156
rect 43032 33212 43096 33216
rect 43032 33156 43036 33212
rect 43036 33156 43092 33212
rect 43092 33156 43096 33212
rect 43032 33152 43096 33156
rect 43112 33212 43176 33216
rect 43112 33156 43116 33212
rect 43116 33156 43172 33212
rect 43172 33156 43176 33212
rect 43112 33152 43176 33156
rect 43192 33212 43256 33216
rect 43192 33156 43196 33212
rect 43196 33156 43252 33212
rect 43252 33156 43256 33212
rect 43192 33152 43256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 27952 32668 28016 32672
rect 27952 32612 27956 32668
rect 27956 32612 28012 32668
rect 28012 32612 28016 32668
rect 27952 32608 28016 32612
rect 28032 32668 28096 32672
rect 28032 32612 28036 32668
rect 28036 32612 28092 32668
rect 28092 32612 28096 32668
rect 28032 32608 28096 32612
rect 28112 32668 28176 32672
rect 28112 32612 28116 32668
rect 28116 32612 28172 32668
rect 28172 32612 28176 32668
rect 28112 32608 28176 32612
rect 28192 32668 28256 32672
rect 28192 32612 28196 32668
rect 28196 32612 28252 32668
rect 28252 32612 28256 32668
rect 28192 32608 28256 32612
rect 37952 32668 38016 32672
rect 37952 32612 37956 32668
rect 37956 32612 38012 32668
rect 38012 32612 38016 32668
rect 37952 32608 38016 32612
rect 38032 32668 38096 32672
rect 38032 32612 38036 32668
rect 38036 32612 38092 32668
rect 38092 32612 38096 32668
rect 38032 32608 38096 32612
rect 38112 32668 38176 32672
rect 38112 32612 38116 32668
rect 38116 32612 38172 32668
rect 38172 32612 38176 32668
rect 38112 32608 38176 32612
rect 38192 32668 38256 32672
rect 38192 32612 38196 32668
rect 38196 32612 38252 32668
rect 38252 32612 38256 32668
rect 38192 32608 38256 32612
rect 47952 32668 48016 32672
rect 47952 32612 47956 32668
rect 47956 32612 48012 32668
rect 48012 32612 48016 32668
rect 47952 32608 48016 32612
rect 48032 32668 48096 32672
rect 48032 32612 48036 32668
rect 48036 32612 48092 32668
rect 48092 32612 48096 32668
rect 48032 32608 48096 32612
rect 48112 32668 48176 32672
rect 48112 32612 48116 32668
rect 48116 32612 48172 32668
rect 48172 32612 48176 32668
rect 48112 32608 48176 32612
rect 48192 32668 48256 32672
rect 48192 32612 48196 32668
rect 48196 32612 48252 32668
rect 48252 32612 48256 32668
rect 48192 32608 48256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 32952 32124 33016 32128
rect 32952 32068 32956 32124
rect 32956 32068 33012 32124
rect 33012 32068 33016 32124
rect 32952 32064 33016 32068
rect 33032 32124 33096 32128
rect 33032 32068 33036 32124
rect 33036 32068 33092 32124
rect 33092 32068 33096 32124
rect 33032 32064 33096 32068
rect 33112 32124 33176 32128
rect 33112 32068 33116 32124
rect 33116 32068 33172 32124
rect 33172 32068 33176 32124
rect 33112 32064 33176 32068
rect 33192 32124 33256 32128
rect 33192 32068 33196 32124
rect 33196 32068 33252 32124
rect 33252 32068 33256 32124
rect 33192 32064 33256 32068
rect 42952 32124 43016 32128
rect 42952 32068 42956 32124
rect 42956 32068 43012 32124
rect 43012 32068 43016 32124
rect 42952 32064 43016 32068
rect 43032 32124 43096 32128
rect 43032 32068 43036 32124
rect 43036 32068 43092 32124
rect 43092 32068 43096 32124
rect 43032 32064 43096 32068
rect 43112 32124 43176 32128
rect 43112 32068 43116 32124
rect 43116 32068 43172 32124
rect 43172 32068 43176 32124
rect 43112 32064 43176 32068
rect 43192 32124 43256 32128
rect 43192 32068 43196 32124
rect 43196 32068 43252 32124
rect 43252 32068 43256 32124
rect 43192 32064 43256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 27952 31580 28016 31584
rect 27952 31524 27956 31580
rect 27956 31524 28012 31580
rect 28012 31524 28016 31580
rect 27952 31520 28016 31524
rect 28032 31580 28096 31584
rect 28032 31524 28036 31580
rect 28036 31524 28092 31580
rect 28092 31524 28096 31580
rect 28032 31520 28096 31524
rect 28112 31580 28176 31584
rect 28112 31524 28116 31580
rect 28116 31524 28172 31580
rect 28172 31524 28176 31580
rect 28112 31520 28176 31524
rect 28192 31580 28256 31584
rect 28192 31524 28196 31580
rect 28196 31524 28252 31580
rect 28252 31524 28256 31580
rect 28192 31520 28256 31524
rect 37952 31580 38016 31584
rect 37952 31524 37956 31580
rect 37956 31524 38012 31580
rect 38012 31524 38016 31580
rect 37952 31520 38016 31524
rect 38032 31580 38096 31584
rect 38032 31524 38036 31580
rect 38036 31524 38092 31580
rect 38092 31524 38096 31580
rect 38032 31520 38096 31524
rect 38112 31580 38176 31584
rect 38112 31524 38116 31580
rect 38116 31524 38172 31580
rect 38172 31524 38176 31580
rect 38112 31520 38176 31524
rect 38192 31580 38256 31584
rect 38192 31524 38196 31580
rect 38196 31524 38252 31580
rect 38252 31524 38256 31580
rect 38192 31520 38256 31524
rect 47952 31580 48016 31584
rect 47952 31524 47956 31580
rect 47956 31524 48012 31580
rect 48012 31524 48016 31580
rect 47952 31520 48016 31524
rect 48032 31580 48096 31584
rect 48032 31524 48036 31580
rect 48036 31524 48092 31580
rect 48092 31524 48096 31580
rect 48032 31520 48096 31524
rect 48112 31580 48176 31584
rect 48112 31524 48116 31580
rect 48116 31524 48172 31580
rect 48172 31524 48176 31580
rect 48112 31520 48176 31524
rect 48192 31580 48256 31584
rect 48192 31524 48196 31580
rect 48196 31524 48252 31580
rect 48252 31524 48256 31580
rect 48192 31520 48256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 32952 31036 33016 31040
rect 32952 30980 32956 31036
rect 32956 30980 33012 31036
rect 33012 30980 33016 31036
rect 32952 30976 33016 30980
rect 33032 31036 33096 31040
rect 33032 30980 33036 31036
rect 33036 30980 33092 31036
rect 33092 30980 33096 31036
rect 33032 30976 33096 30980
rect 33112 31036 33176 31040
rect 33112 30980 33116 31036
rect 33116 30980 33172 31036
rect 33172 30980 33176 31036
rect 33112 30976 33176 30980
rect 33192 31036 33256 31040
rect 33192 30980 33196 31036
rect 33196 30980 33252 31036
rect 33252 30980 33256 31036
rect 33192 30976 33256 30980
rect 42952 31036 43016 31040
rect 42952 30980 42956 31036
rect 42956 30980 43012 31036
rect 43012 30980 43016 31036
rect 42952 30976 43016 30980
rect 43032 31036 43096 31040
rect 43032 30980 43036 31036
rect 43036 30980 43092 31036
rect 43092 30980 43096 31036
rect 43032 30976 43096 30980
rect 43112 31036 43176 31040
rect 43112 30980 43116 31036
rect 43116 30980 43172 31036
rect 43172 30980 43176 31036
rect 43112 30976 43176 30980
rect 43192 31036 43256 31040
rect 43192 30980 43196 31036
rect 43196 30980 43252 31036
rect 43252 30980 43256 31036
rect 43192 30976 43256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 27952 30492 28016 30496
rect 27952 30436 27956 30492
rect 27956 30436 28012 30492
rect 28012 30436 28016 30492
rect 27952 30432 28016 30436
rect 28032 30492 28096 30496
rect 28032 30436 28036 30492
rect 28036 30436 28092 30492
rect 28092 30436 28096 30492
rect 28032 30432 28096 30436
rect 28112 30492 28176 30496
rect 28112 30436 28116 30492
rect 28116 30436 28172 30492
rect 28172 30436 28176 30492
rect 28112 30432 28176 30436
rect 28192 30492 28256 30496
rect 28192 30436 28196 30492
rect 28196 30436 28252 30492
rect 28252 30436 28256 30492
rect 28192 30432 28256 30436
rect 37952 30492 38016 30496
rect 37952 30436 37956 30492
rect 37956 30436 38012 30492
rect 38012 30436 38016 30492
rect 37952 30432 38016 30436
rect 38032 30492 38096 30496
rect 38032 30436 38036 30492
rect 38036 30436 38092 30492
rect 38092 30436 38096 30492
rect 38032 30432 38096 30436
rect 38112 30492 38176 30496
rect 38112 30436 38116 30492
rect 38116 30436 38172 30492
rect 38172 30436 38176 30492
rect 38112 30432 38176 30436
rect 38192 30492 38256 30496
rect 38192 30436 38196 30492
rect 38196 30436 38252 30492
rect 38252 30436 38256 30492
rect 38192 30432 38256 30436
rect 47952 30492 48016 30496
rect 47952 30436 47956 30492
rect 47956 30436 48012 30492
rect 48012 30436 48016 30492
rect 47952 30432 48016 30436
rect 48032 30492 48096 30496
rect 48032 30436 48036 30492
rect 48036 30436 48092 30492
rect 48092 30436 48096 30492
rect 48032 30432 48096 30436
rect 48112 30492 48176 30496
rect 48112 30436 48116 30492
rect 48116 30436 48172 30492
rect 48172 30436 48176 30492
rect 48112 30432 48176 30436
rect 48192 30492 48256 30496
rect 48192 30436 48196 30492
rect 48196 30436 48252 30492
rect 48252 30436 48256 30492
rect 48192 30432 48256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 32952 29948 33016 29952
rect 32952 29892 32956 29948
rect 32956 29892 33012 29948
rect 33012 29892 33016 29948
rect 32952 29888 33016 29892
rect 33032 29948 33096 29952
rect 33032 29892 33036 29948
rect 33036 29892 33092 29948
rect 33092 29892 33096 29948
rect 33032 29888 33096 29892
rect 33112 29948 33176 29952
rect 33112 29892 33116 29948
rect 33116 29892 33172 29948
rect 33172 29892 33176 29948
rect 33112 29888 33176 29892
rect 33192 29948 33256 29952
rect 33192 29892 33196 29948
rect 33196 29892 33252 29948
rect 33252 29892 33256 29948
rect 33192 29888 33256 29892
rect 42952 29948 43016 29952
rect 42952 29892 42956 29948
rect 42956 29892 43012 29948
rect 43012 29892 43016 29948
rect 42952 29888 43016 29892
rect 43032 29948 43096 29952
rect 43032 29892 43036 29948
rect 43036 29892 43092 29948
rect 43092 29892 43096 29948
rect 43032 29888 43096 29892
rect 43112 29948 43176 29952
rect 43112 29892 43116 29948
rect 43116 29892 43172 29948
rect 43172 29892 43176 29948
rect 43112 29888 43176 29892
rect 43192 29948 43256 29952
rect 43192 29892 43196 29948
rect 43196 29892 43252 29948
rect 43252 29892 43256 29948
rect 43192 29888 43256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 27952 29404 28016 29408
rect 27952 29348 27956 29404
rect 27956 29348 28012 29404
rect 28012 29348 28016 29404
rect 27952 29344 28016 29348
rect 28032 29404 28096 29408
rect 28032 29348 28036 29404
rect 28036 29348 28092 29404
rect 28092 29348 28096 29404
rect 28032 29344 28096 29348
rect 28112 29404 28176 29408
rect 28112 29348 28116 29404
rect 28116 29348 28172 29404
rect 28172 29348 28176 29404
rect 28112 29344 28176 29348
rect 28192 29404 28256 29408
rect 28192 29348 28196 29404
rect 28196 29348 28252 29404
rect 28252 29348 28256 29404
rect 28192 29344 28256 29348
rect 37952 29404 38016 29408
rect 37952 29348 37956 29404
rect 37956 29348 38012 29404
rect 38012 29348 38016 29404
rect 37952 29344 38016 29348
rect 38032 29404 38096 29408
rect 38032 29348 38036 29404
rect 38036 29348 38092 29404
rect 38092 29348 38096 29404
rect 38032 29344 38096 29348
rect 38112 29404 38176 29408
rect 38112 29348 38116 29404
rect 38116 29348 38172 29404
rect 38172 29348 38176 29404
rect 38112 29344 38176 29348
rect 38192 29404 38256 29408
rect 38192 29348 38196 29404
rect 38196 29348 38252 29404
rect 38252 29348 38256 29404
rect 38192 29344 38256 29348
rect 47952 29404 48016 29408
rect 47952 29348 47956 29404
rect 47956 29348 48012 29404
rect 48012 29348 48016 29404
rect 47952 29344 48016 29348
rect 48032 29404 48096 29408
rect 48032 29348 48036 29404
rect 48036 29348 48092 29404
rect 48092 29348 48096 29404
rect 48032 29344 48096 29348
rect 48112 29404 48176 29408
rect 48112 29348 48116 29404
rect 48116 29348 48172 29404
rect 48172 29348 48176 29404
rect 48112 29344 48176 29348
rect 48192 29404 48256 29408
rect 48192 29348 48196 29404
rect 48196 29348 48252 29404
rect 48252 29348 48256 29404
rect 48192 29344 48256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 32952 28860 33016 28864
rect 32952 28804 32956 28860
rect 32956 28804 33012 28860
rect 33012 28804 33016 28860
rect 32952 28800 33016 28804
rect 33032 28860 33096 28864
rect 33032 28804 33036 28860
rect 33036 28804 33092 28860
rect 33092 28804 33096 28860
rect 33032 28800 33096 28804
rect 33112 28860 33176 28864
rect 33112 28804 33116 28860
rect 33116 28804 33172 28860
rect 33172 28804 33176 28860
rect 33112 28800 33176 28804
rect 33192 28860 33256 28864
rect 33192 28804 33196 28860
rect 33196 28804 33252 28860
rect 33252 28804 33256 28860
rect 33192 28800 33256 28804
rect 42952 28860 43016 28864
rect 42952 28804 42956 28860
rect 42956 28804 43012 28860
rect 43012 28804 43016 28860
rect 42952 28800 43016 28804
rect 43032 28860 43096 28864
rect 43032 28804 43036 28860
rect 43036 28804 43092 28860
rect 43092 28804 43096 28860
rect 43032 28800 43096 28804
rect 43112 28860 43176 28864
rect 43112 28804 43116 28860
rect 43116 28804 43172 28860
rect 43172 28804 43176 28860
rect 43112 28800 43176 28804
rect 43192 28860 43256 28864
rect 43192 28804 43196 28860
rect 43196 28804 43252 28860
rect 43252 28804 43256 28860
rect 43192 28800 43256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 27952 28316 28016 28320
rect 27952 28260 27956 28316
rect 27956 28260 28012 28316
rect 28012 28260 28016 28316
rect 27952 28256 28016 28260
rect 28032 28316 28096 28320
rect 28032 28260 28036 28316
rect 28036 28260 28092 28316
rect 28092 28260 28096 28316
rect 28032 28256 28096 28260
rect 28112 28316 28176 28320
rect 28112 28260 28116 28316
rect 28116 28260 28172 28316
rect 28172 28260 28176 28316
rect 28112 28256 28176 28260
rect 28192 28316 28256 28320
rect 28192 28260 28196 28316
rect 28196 28260 28252 28316
rect 28252 28260 28256 28316
rect 28192 28256 28256 28260
rect 37952 28316 38016 28320
rect 37952 28260 37956 28316
rect 37956 28260 38012 28316
rect 38012 28260 38016 28316
rect 37952 28256 38016 28260
rect 38032 28316 38096 28320
rect 38032 28260 38036 28316
rect 38036 28260 38092 28316
rect 38092 28260 38096 28316
rect 38032 28256 38096 28260
rect 38112 28316 38176 28320
rect 38112 28260 38116 28316
rect 38116 28260 38172 28316
rect 38172 28260 38176 28316
rect 38112 28256 38176 28260
rect 38192 28316 38256 28320
rect 38192 28260 38196 28316
rect 38196 28260 38252 28316
rect 38252 28260 38256 28316
rect 38192 28256 38256 28260
rect 47952 28316 48016 28320
rect 47952 28260 47956 28316
rect 47956 28260 48012 28316
rect 48012 28260 48016 28316
rect 47952 28256 48016 28260
rect 48032 28316 48096 28320
rect 48032 28260 48036 28316
rect 48036 28260 48092 28316
rect 48092 28260 48096 28316
rect 48032 28256 48096 28260
rect 48112 28316 48176 28320
rect 48112 28260 48116 28316
rect 48116 28260 48172 28316
rect 48172 28260 48176 28316
rect 48112 28256 48176 28260
rect 48192 28316 48256 28320
rect 48192 28260 48196 28316
rect 48196 28260 48252 28316
rect 48252 28260 48256 28316
rect 48192 28256 48256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 32952 27772 33016 27776
rect 32952 27716 32956 27772
rect 32956 27716 33012 27772
rect 33012 27716 33016 27772
rect 32952 27712 33016 27716
rect 33032 27772 33096 27776
rect 33032 27716 33036 27772
rect 33036 27716 33092 27772
rect 33092 27716 33096 27772
rect 33032 27712 33096 27716
rect 33112 27772 33176 27776
rect 33112 27716 33116 27772
rect 33116 27716 33172 27772
rect 33172 27716 33176 27772
rect 33112 27712 33176 27716
rect 33192 27772 33256 27776
rect 33192 27716 33196 27772
rect 33196 27716 33252 27772
rect 33252 27716 33256 27772
rect 33192 27712 33256 27716
rect 42952 27772 43016 27776
rect 42952 27716 42956 27772
rect 42956 27716 43012 27772
rect 43012 27716 43016 27772
rect 42952 27712 43016 27716
rect 43032 27772 43096 27776
rect 43032 27716 43036 27772
rect 43036 27716 43092 27772
rect 43092 27716 43096 27772
rect 43032 27712 43096 27716
rect 43112 27772 43176 27776
rect 43112 27716 43116 27772
rect 43116 27716 43172 27772
rect 43172 27716 43176 27772
rect 43112 27712 43176 27716
rect 43192 27772 43256 27776
rect 43192 27716 43196 27772
rect 43196 27716 43252 27772
rect 43252 27716 43256 27772
rect 43192 27712 43256 27716
rect 18460 27508 18524 27572
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 27952 27228 28016 27232
rect 27952 27172 27956 27228
rect 27956 27172 28012 27228
rect 28012 27172 28016 27228
rect 27952 27168 28016 27172
rect 28032 27228 28096 27232
rect 28032 27172 28036 27228
rect 28036 27172 28092 27228
rect 28092 27172 28096 27228
rect 28032 27168 28096 27172
rect 28112 27228 28176 27232
rect 28112 27172 28116 27228
rect 28116 27172 28172 27228
rect 28172 27172 28176 27228
rect 28112 27168 28176 27172
rect 28192 27228 28256 27232
rect 28192 27172 28196 27228
rect 28196 27172 28252 27228
rect 28252 27172 28256 27228
rect 28192 27168 28256 27172
rect 37952 27228 38016 27232
rect 37952 27172 37956 27228
rect 37956 27172 38012 27228
rect 38012 27172 38016 27228
rect 37952 27168 38016 27172
rect 38032 27228 38096 27232
rect 38032 27172 38036 27228
rect 38036 27172 38092 27228
rect 38092 27172 38096 27228
rect 38032 27168 38096 27172
rect 38112 27228 38176 27232
rect 38112 27172 38116 27228
rect 38116 27172 38172 27228
rect 38172 27172 38176 27228
rect 38112 27168 38176 27172
rect 38192 27228 38256 27232
rect 38192 27172 38196 27228
rect 38196 27172 38252 27228
rect 38252 27172 38256 27228
rect 38192 27168 38256 27172
rect 47952 27228 48016 27232
rect 47952 27172 47956 27228
rect 47956 27172 48012 27228
rect 48012 27172 48016 27228
rect 47952 27168 48016 27172
rect 48032 27228 48096 27232
rect 48032 27172 48036 27228
rect 48036 27172 48092 27228
rect 48092 27172 48096 27228
rect 48032 27168 48096 27172
rect 48112 27228 48176 27232
rect 48112 27172 48116 27228
rect 48116 27172 48172 27228
rect 48172 27172 48176 27228
rect 48112 27168 48176 27172
rect 48192 27228 48256 27232
rect 48192 27172 48196 27228
rect 48196 27172 48252 27228
rect 48252 27172 48256 27228
rect 48192 27168 48256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 32952 26684 33016 26688
rect 32952 26628 32956 26684
rect 32956 26628 33012 26684
rect 33012 26628 33016 26684
rect 32952 26624 33016 26628
rect 33032 26684 33096 26688
rect 33032 26628 33036 26684
rect 33036 26628 33092 26684
rect 33092 26628 33096 26684
rect 33032 26624 33096 26628
rect 33112 26684 33176 26688
rect 33112 26628 33116 26684
rect 33116 26628 33172 26684
rect 33172 26628 33176 26684
rect 33112 26624 33176 26628
rect 33192 26684 33256 26688
rect 33192 26628 33196 26684
rect 33196 26628 33252 26684
rect 33252 26628 33256 26684
rect 33192 26624 33256 26628
rect 42952 26684 43016 26688
rect 42952 26628 42956 26684
rect 42956 26628 43012 26684
rect 43012 26628 43016 26684
rect 42952 26624 43016 26628
rect 43032 26684 43096 26688
rect 43032 26628 43036 26684
rect 43036 26628 43092 26684
rect 43092 26628 43096 26684
rect 43032 26624 43096 26628
rect 43112 26684 43176 26688
rect 43112 26628 43116 26684
rect 43116 26628 43172 26684
rect 43172 26628 43176 26684
rect 43112 26624 43176 26628
rect 43192 26684 43256 26688
rect 43192 26628 43196 26684
rect 43196 26628 43252 26684
rect 43252 26628 43256 26684
rect 43192 26624 43256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 27952 26140 28016 26144
rect 27952 26084 27956 26140
rect 27956 26084 28012 26140
rect 28012 26084 28016 26140
rect 27952 26080 28016 26084
rect 28032 26140 28096 26144
rect 28032 26084 28036 26140
rect 28036 26084 28092 26140
rect 28092 26084 28096 26140
rect 28032 26080 28096 26084
rect 28112 26140 28176 26144
rect 28112 26084 28116 26140
rect 28116 26084 28172 26140
rect 28172 26084 28176 26140
rect 28112 26080 28176 26084
rect 28192 26140 28256 26144
rect 28192 26084 28196 26140
rect 28196 26084 28252 26140
rect 28252 26084 28256 26140
rect 28192 26080 28256 26084
rect 37952 26140 38016 26144
rect 37952 26084 37956 26140
rect 37956 26084 38012 26140
rect 38012 26084 38016 26140
rect 37952 26080 38016 26084
rect 38032 26140 38096 26144
rect 38032 26084 38036 26140
rect 38036 26084 38092 26140
rect 38092 26084 38096 26140
rect 38032 26080 38096 26084
rect 38112 26140 38176 26144
rect 38112 26084 38116 26140
rect 38116 26084 38172 26140
rect 38172 26084 38176 26140
rect 38112 26080 38176 26084
rect 38192 26140 38256 26144
rect 38192 26084 38196 26140
rect 38196 26084 38252 26140
rect 38252 26084 38256 26140
rect 38192 26080 38256 26084
rect 47952 26140 48016 26144
rect 47952 26084 47956 26140
rect 47956 26084 48012 26140
rect 48012 26084 48016 26140
rect 47952 26080 48016 26084
rect 48032 26140 48096 26144
rect 48032 26084 48036 26140
rect 48036 26084 48092 26140
rect 48092 26084 48096 26140
rect 48032 26080 48096 26084
rect 48112 26140 48176 26144
rect 48112 26084 48116 26140
rect 48116 26084 48172 26140
rect 48172 26084 48176 26140
rect 48112 26080 48176 26084
rect 48192 26140 48256 26144
rect 48192 26084 48196 26140
rect 48196 26084 48252 26140
rect 48252 26084 48256 26140
rect 48192 26080 48256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 32952 25596 33016 25600
rect 32952 25540 32956 25596
rect 32956 25540 33012 25596
rect 33012 25540 33016 25596
rect 32952 25536 33016 25540
rect 33032 25596 33096 25600
rect 33032 25540 33036 25596
rect 33036 25540 33092 25596
rect 33092 25540 33096 25596
rect 33032 25536 33096 25540
rect 33112 25596 33176 25600
rect 33112 25540 33116 25596
rect 33116 25540 33172 25596
rect 33172 25540 33176 25596
rect 33112 25536 33176 25540
rect 33192 25596 33256 25600
rect 33192 25540 33196 25596
rect 33196 25540 33252 25596
rect 33252 25540 33256 25596
rect 33192 25536 33256 25540
rect 42952 25596 43016 25600
rect 42952 25540 42956 25596
rect 42956 25540 43012 25596
rect 43012 25540 43016 25596
rect 42952 25536 43016 25540
rect 43032 25596 43096 25600
rect 43032 25540 43036 25596
rect 43036 25540 43092 25596
rect 43092 25540 43096 25596
rect 43032 25536 43096 25540
rect 43112 25596 43176 25600
rect 43112 25540 43116 25596
rect 43116 25540 43172 25596
rect 43172 25540 43176 25596
rect 43112 25536 43176 25540
rect 43192 25596 43256 25600
rect 43192 25540 43196 25596
rect 43196 25540 43252 25596
rect 43252 25540 43256 25596
rect 43192 25536 43256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 27952 25052 28016 25056
rect 27952 24996 27956 25052
rect 27956 24996 28012 25052
rect 28012 24996 28016 25052
rect 27952 24992 28016 24996
rect 28032 25052 28096 25056
rect 28032 24996 28036 25052
rect 28036 24996 28092 25052
rect 28092 24996 28096 25052
rect 28032 24992 28096 24996
rect 28112 25052 28176 25056
rect 28112 24996 28116 25052
rect 28116 24996 28172 25052
rect 28172 24996 28176 25052
rect 28112 24992 28176 24996
rect 28192 25052 28256 25056
rect 28192 24996 28196 25052
rect 28196 24996 28252 25052
rect 28252 24996 28256 25052
rect 28192 24992 28256 24996
rect 37952 25052 38016 25056
rect 37952 24996 37956 25052
rect 37956 24996 38012 25052
rect 38012 24996 38016 25052
rect 37952 24992 38016 24996
rect 38032 25052 38096 25056
rect 38032 24996 38036 25052
rect 38036 24996 38092 25052
rect 38092 24996 38096 25052
rect 38032 24992 38096 24996
rect 38112 25052 38176 25056
rect 38112 24996 38116 25052
rect 38116 24996 38172 25052
rect 38172 24996 38176 25052
rect 38112 24992 38176 24996
rect 38192 25052 38256 25056
rect 38192 24996 38196 25052
rect 38196 24996 38252 25052
rect 38252 24996 38256 25052
rect 38192 24992 38256 24996
rect 47952 25052 48016 25056
rect 47952 24996 47956 25052
rect 47956 24996 48012 25052
rect 48012 24996 48016 25052
rect 47952 24992 48016 24996
rect 48032 25052 48096 25056
rect 48032 24996 48036 25052
rect 48036 24996 48092 25052
rect 48092 24996 48096 25052
rect 48032 24992 48096 24996
rect 48112 25052 48176 25056
rect 48112 24996 48116 25052
rect 48116 24996 48172 25052
rect 48172 24996 48176 25052
rect 48112 24992 48176 24996
rect 48192 25052 48256 25056
rect 48192 24996 48196 25052
rect 48196 24996 48252 25052
rect 48252 24996 48256 25052
rect 48192 24992 48256 24996
rect 34100 24788 34164 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 22692 17036 22756 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 24716 14316 24780 14380
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 21219 52052 21285 52053
rect 21219 51988 21220 52052
rect 21284 51988 21285 52052
rect 21219 51987 21285 51988
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 21222 40221 21282 51987
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 27944 54432 28264 54448
rect 27944 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28264 54432
rect 27944 53344 28264 54368
rect 27944 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28264 53344
rect 27944 52256 28264 53280
rect 27944 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28264 52256
rect 27944 51168 28264 52192
rect 27944 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28264 51168
rect 27944 50080 28264 51104
rect 27944 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28264 50080
rect 27944 48992 28264 50016
rect 27944 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28264 48992
rect 27944 47904 28264 48928
rect 27944 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28264 47904
rect 24899 47020 24965 47021
rect 24899 46956 24900 47020
rect 24964 46956 24965 47020
rect 24899 46955 24965 46956
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 21219 40220 21285 40221
rect 21219 40156 21220 40220
rect 21284 40156 21285 40220
rect 21219 40155 21285 40156
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 22944 39744 23264 40768
rect 24902 39949 24962 46955
rect 27944 46816 28264 47840
rect 32944 53888 33264 54448
rect 32944 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33264 53888
rect 32944 52800 33264 53824
rect 32944 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33264 52800
rect 32944 51712 33264 52736
rect 32944 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33264 51712
rect 32944 50624 33264 51648
rect 32944 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33264 50624
rect 32944 49536 33264 50560
rect 32944 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33264 49536
rect 32944 48448 33264 49472
rect 32944 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33264 48448
rect 32944 47360 33264 48384
rect 32944 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33264 47360
rect 28763 47020 28829 47021
rect 28763 46956 28764 47020
rect 28828 46956 28829 47020
rect 28763 46955 28829 46956
rect 27944 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28264 46816
rect 25267 45932 25333 45933
rect 25267 45868 25268 45932
rect 25332 45868 25333 45932
rect 25267 45867 25333 45868
rect 25270 41309 25330 45867
rect 27944 45728 28264 46752
rect 27944 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28264 45728
rect 27944 44640 28264 45664
rect 27944 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28264 44640
rect 27944 43552 28264 44576
rect 28395 44300 28461 44301
rect 28395 44236 28396 44300
rect 28460 44236 28461 44300
rect 28395 44235 28461 44236
rect 27944 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28264 43552
rect 27944 42464 28264 43488
rect 27944 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28264 42464
rect 27944 41376 28264 42400
rect 27944 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28264 41376
rect 25267 41308 25333 41309
rect 25267 41244 25268 41308
rect 25332 41244 25333 41308
rect 25267 41243 25333 41244
rect 27944 40288 28264 41312
rect 27944 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28264 40288
rect 24899 39948 24965 39949
rect 24899 39884 24900 39948
rect 24964 39884 24965 39948
rect 24899 39883 24965 39884
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 24902 39405 24962 39883
rect 24899 39404 24965 39405
rect 24899 39340 24900 39404
rect 24964 39340 24965 39404
rect 24899 39339 24965 39340
rect 27944 39200 28264 40224
rect 27944 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28264 39200
rect 26187 38996 26253 38997
rect 26187 38932 26188 38996
rect 26252 38932 26253 38996
rect 26187 38931 26253 38932
rect 24715 38860 24781 38861
rect 24715 38796 24716 38860
rect 24780 38796 24781 38860
rect 24715 38795 24781 38796
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 18459 35052 18525 35053
rect 18459 34988 18460 35052
rect 18524 34988 18525 35052
rect 18459 34987 18525 34988
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 18462 27573 18522 34987
rect 22691 34780 22757 34781
rect 22691 34716 22692 34780
rect 22756 34716 22757 34780
rect 22691 34715 22757 34716
rect 18459 27572 18525 27573
rect 18459 27508 18460 27572
rect 18524 27508 18525 27572
rect 18459 27507 18525 27508
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 22694 17101 22754 34715
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22691 17100 22757 17101
rect 22691 17036 22692 17100
rect 22756 17036 22757 17100
rect 22691 17035 22757 17036
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 24718 14381 24778 38795
rect 26190 36685 26250 38931
rect 27944 38112 28264 39136
rect 27944 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28264 38112
rect 27944 37024 28264 38048
rect 28398 37773 28458 44235
rect 28766 39541 28826 46955
rect 32944 46272 33264 47296
rect 32944 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33264 46272
rect 32944 45184 33264 46208
rect 32944 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33264 45184
rect 30235 44300 30301 44301
rect 30235 44236 30236 44300
rect 30300 44236 30301 44300
rect 30235 44235 30301 44236
rect 28763 39540 28829 39541
rect 28763 39476 28764 39540
rect 28828 39476 28829 39540
rect 28763 39475 28829 39476
rect 28395 37772 28461 37773
rect 28395 37708 28396 37772
rect 28460 37708 28461 37772
rect 28395 37707 28461 37708
rect 27944 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28264 37024
rect 26187 36684 26253 36685
rect 26187 36620 26188 36684
rect 26252 36620 26253 36684
rect 26187 36619 26253 36620
rect 27944 35936 28264 36960
rect 27944 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28264 35936
rect 27944 34848 28264 35872
rect 30238 35325 30298 44235
rect 32944 44096 33264 45120
rect 32944 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33264 44096
rect 32944 43008 33264 44032
rect 32944 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33264 43008
rect 32944 41920 33264 42944
rect 32944 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33264 41920
rect 32944 40832 33264 41856
rect 32944 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33264 40832
rect 32944 39744 33264 40768
rect 32944 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33264 39744
rect 32944 38656 33264 39680
rect 37944 54432 38264 54448
rect 37944 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38264 54432
rect 37944 53344 38264 54368
rect 37944 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38264 53344
rect 37944 52256 38264 53280
rect 37944 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38264 52256
rect 37944 51168 38264 52192
rect 37944 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38264 51168
rect 37944 50080 38264 51104
rect 37944 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38264 50080
rect 37944 48992 38264 50016
rect 37944 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38264 48992
rect 37944 47904 38264 48928
rect 37944 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38264 47904
rect 37944 46816 38264 47840
rect 37944 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38264 46816
rect 37944 45728 38264 46752
rect 37944 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38264 45728
rect 37944 44640 38264 45664
rect 37944 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38264 44640
rect 37944 43552 38264 44576
rect 37944 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38264 43552
rect 37944 42464 38264 43488
rect 37944 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38264 42464
rect 37944 41376 38264 42400
rect 37944 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38264 41376
rect 37944 40288 38264 41312
rect 37944 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38264 40288
rect 34099 39268 34165 39269
rect 34099 39204 34100 39268
rect 34164 39204 34165 39268
rect 34099 39203 34165 39204
rect 32944 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33264 38656
rect 32944 37568 33264 38592
rect 32944 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33264 37568
rect 32944 36480 33264 37504
rect 32944 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33264 36480
rect 32944 35392 33264 36416
rect 32944 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33264 35392
rect 30235 35324 30301 35325
rect 30235 35260 30236 35324
rect 30300 35260 30301 35324
rect 30235 35259 30301 35260
rect 27944 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28264 34848
rect 27944 33760 28264 34784
rect 27944 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28264 33760
rect 27944 32672 28264 33696
rect 27944 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28264 32672
rect 27944 31584 28264 32608
rect 27944 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28264 31584
rect 27944 30496 28264 31520
rect 27944 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28264 30496
rect 27944 29408 28264 30432
rect 27944 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28264 29408
rect 27944 28320 28264 29344
rect 27944 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28264 28320
rect 27944 27232 28264 28256
rect 27944 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28264 27232
rect 27944 26144 28264 27168
rect 27944 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28264 26144
rect 27944 25056 28264 26080
rect 27944 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28264 25056
rect 27944 23968 28264 24992
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 24715 14380 24781 14381
rect 24715 14316 24716 14380
rect 24780 14316 24781 14380
rect 24715 14315 24781 14316
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 34304 33264 35328
rect 32944 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33264 34304
rect 32944 33216 33264 34240
rect 32944 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33264 33216
rect 32944 32128 33264 33152
rect 32944 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33264 32128
rect 32944 31040 33264 32064
rect 32944 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33264 31040
rect 32944 29952 33264 30976
rect 32944 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33264 29952
rect 32944 28864 33264 29888
rect 32944 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33264 28864
rect 32944 27776 33264 28800
rect 32944 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33264 27776
rect 32944 26688 33264 27712
rect 32944 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33264 26688
rect 32944 25600 33264 26624
rect 32944 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33264 25600
rect 32944 24512 33264 25536
rect 34102 24853 34162 39203
rect 37944 39200 38264 40224
rect 37944 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38264 39200
rect 37944 38112 38264 39136
rect 37944 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38264 38112
rect 37944 37024 38264 38048
rect 37944 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38264 37024
rect 37944 35936 38264 36960
rect 37944 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38264 35936
rect 37944 34848 38264 35872
rect 37944 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38264 34848
rect 37944 33760 38264 34784
rect 37944 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38264 33760
rect 37944 32672 38264 33696
rect 37944 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38264 32672
rect 37944 31584 38264 32608
rect 37944 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38264 31584
rect 37944 30496 38264 31520
rect 37944 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38264 30496
rect 37944 29408 38264 30432
rect 37944 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38264 29408
rect 37944 28320 38264 29344
rect 37944 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38264 28320
rect 37944 27232 38264 28256
rect 37944 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38264 27232
rect 37944 26144 38264 27168
rect 37944 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38264 26144
rect 37944 25056 38264 26080
rect 37944 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38264 25056
rect 34099 24852 34165 24853
rect 34099 24788 34100 24852
rect 34164 24788 34165 24852
rect 34099 24787 34165 24788
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24992
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 53888 43264 54448
rect 42944 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43264 53888
rect 42944 52800 43264 53824
rect 42944 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43264 52800
rect 42944 51712 43264 52736
rect 42944 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43264 51712
rect 42944 50624 43264 51648
rect 42944 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43264 50624
rect 42944 49536 43264 50560
rect 42944 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43264 49536
rect 42944 48448 43264 49472
rect 42944 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43264 48448
rect 42944 47360 43264 48384
rect 42944 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43264 47360
rect 42944 46272 43264 47296
rect 42944 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43264 46272
rect 42944 45184 43264 46208
rect 42944 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43264 45184
rect 42944 44096 43264 45120
rect 42944 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43264 44096
rect 42944 43008 43264 44032
rect 42944 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43264 43008
rect 42944 41920 43264 42944
rect 42944 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43264 41920
rect 42944 40832 43264 41856
rect 42944 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43264 40832
rect 42944 39744 43264 40768
rect 42944 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43264 39744
rect 42944 38656 43264 39680
rect 42944 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43264 38656
rect 42944 37568 43264 38592
rect 42944 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43264 37568
rect 42944 36480 43264 37504
rect 42944 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43264 36480
rect 42944 35392 43264 36416
rect 42944 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43264 35392
rect 42944 34304 43264 35328
rect 42944 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43264 34304
rect 42944 33216 43264 34240
rect 42944 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43264 33216
rect 42944 32128 43264 33152
rect 42944 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43264 32128
rect 42944 31040 43264 32064
rect 42944 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43264 31040
rect 42944 29952 43264 30976
rect 42944 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43264 29952
rect 42944 28864 43264 29888
rect 42944 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43264 28864
rect 42944 27776 43264 28800
rect 42944 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43264 27776
rect 42944 26688 43264 27712
rect 42944 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43264 26688
rect 42944 25600 43264 26624
rect 42944 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43264 25600
rect 42944 24512 43264 25536
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 54432 48264 54448
rect 47944 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48264 54432
rect 47944 53344 48264 54368
rect 47944 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48264 53344
rect 47944 52256 48264 53280
rect 47944 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48264 52256
rect 47944 51168 48264 52192
rect 47944 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48264 51168
rect 47944 50080 48264 51104
rect 47944 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48264 50080
rect 47944 48992 48264 50016
rect 47944 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48264 48992
rect 47944 47904 48264 48928
rect 47944 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48264 47904
rect 47944 46816 48264 47840
rect 47944 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48264 46816
rect 47944 45728 48264 46752
rect 47944 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48264 45728
rect 47944 44640 48264 45664
rect 47944 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48264 44640
rect 47944 43552 48264 44576
rect 47944 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48264 43552
rect 47944 42464 48264 43488
rect 47944 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48264 42464
rect 47944 41376 48264 42400
rect 47944 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48264 41376
rect 47944 40288 48264 41312
rect 47944 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48264 40288
rect 47944 39200 48264 40224
rect 47944 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48264 39200
rect 47944 38112 48264 39136
rect 47944 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48264 38112
rect 47944 37024 48264 38048
rect 47944 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48264 37024
rect 47944 35936 48264 36960
rect 47944 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48264 35936
rect 47944 34848 48264 35872
rect 47944 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48264 34848
rect 47944 33760 48264 34784
rect 47944 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48264 33760
rect 47944 32672 48264 33696
rect 47944 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48264 32672
rect 47944 31584 48264 32608
rect 47944 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48264 31584
rect 47944 30496 48264 31520
rect 47944 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48264 30496
rect 47944 29408 48264 30432
rect 47944 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48264 29408
rect 47944 28320 48264 29344
rect 47944 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48264 28320
rect 47944 27232 48264 28256
rect 47944 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48264 27232
rect 47944 26144 48264 27168
rect 47944 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48264 26144
rect 47944 25056 48264 26080
rect 47944 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48264 25056
rect 47944 23968 48264 24992
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13432 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 10580 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 7728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 10856 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 12512 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 16836 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 8372 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 10764 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 11500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 11868 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 8280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 16652 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 16008 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 13156 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 12052 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 13064 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 14996 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 6716 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 11684 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 12696 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 11960 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 8464 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 5428 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 10856 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 7636 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 5428 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform 1 0 7360 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 36156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 37260 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 43608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 37536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 44068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 38088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 37812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 37996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 44344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 37904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 40020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 38548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 43792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 39008 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 43976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 39836 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 39468 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 38732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 44436 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 45080 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 38824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 46460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 45724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 45172 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 44344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _165_
timestamp 1676037725
transform 1 0 3680 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 5244 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1676037725
transform 1 0 4416 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1676037725
transform 1 0 8280 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 9108 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 8096 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 9108 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1676037725
transform 1 0 9936 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1676037725
transform 1 0 9844 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 19964 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1676037725
transform 1 0 13248 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1676037725
transform 1 0 13248 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 13248 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1676037725
transform 1 0 13892 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1676037725
transform 1 0 16008 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform 1 0 16836 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 16652 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 19780 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 21160 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 21988 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1676037725
transform 1 0 22448 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 21988 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 23184 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1676037725
transform 1 0 23092 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1676037725
transform 1 0 23828 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1676037725
transform 1 0 23552 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform 1 0 13432 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _195_
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _196_
timestamp 1676037725
transform 1 0 17296 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _197_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _199_
timestamp 1676037725
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _200_
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1676037725
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 20148 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 22448 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 20608 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 17572 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 14720 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 12328 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 28612 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 24380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 17572 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 38180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 36708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 38824 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 15456 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 38088 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 12512 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 37628 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 26312 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 26220 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 27048 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 32200 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 35604 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 14168 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 17296 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 36064 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 14076 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 30176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 39284 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 38088 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 33488 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 37444 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 31464 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 34684 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19688 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 19688 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19872 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17296 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 17112 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14076 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 14628 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15824 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15916 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 10672 0 1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19044 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18032 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 22816 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 17020 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 19688 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23184 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19780 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 20884 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12328 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19412 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 17848 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 20424 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17388 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 16560 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 20424 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 8924 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 15548 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 18492 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 16928 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256
timestamp 1676037725
transform 1 0 14628 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 13156 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14444 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 15364 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 15364 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14444 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14536 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 16376 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 14352 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16652 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 15548 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 17848 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257
timestamp 1676037725
transform 1 0 19412 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 14352 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 13064 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15640 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29808 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22908 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11224 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 27968 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 21896 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24748 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 23368 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 30728 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32660 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25852 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 19504 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 18584 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 22172 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 20700 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 19780 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 22448 0 1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 27416 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 28244 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 27140 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 29716 0 1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 32292 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 33396 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 32384 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 34868 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1676037725
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1676037725
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_342
timestamp 1676037725
transform 1 0 32568 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1676037725
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1676037725
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1676037725
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_485
timestamp 1676037725
transform 1 0 45724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_497
timestamp 1676037725
transform 1 0 46828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1676037725
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1676037725
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_21
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_33
timestamp 1676037725
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1676037725
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1676037725
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_157
timestamp 1676037725
transform 1 0 15548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_169
timestamp 1676037725
transform 1 0 16652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_175
timestamp 1676037725
transform 1 0 17204 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_180
timestamp 1676037725
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1676037725
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_203
timestamp 1676037725
transform 1 0 19780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_227
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_239
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1676037725
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_133
timestamp 1676037725
transform 1 0 13340 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_138
timestamp 1676037725
transform 1 0 13800 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_150
timestamp 1676037725
transform 1 0 14904 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1676037725
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp 1676037725
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_217
timestamp 1676037725
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_223
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_235
timestamp 1676037725
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_271
timestamp 1676037725
transform 1 0 26036 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_275
timestamp 1676037725
transform 1 0 26404 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_280
timestamp 1676037725
transform 1 0 26864 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_292
timestamp 1676037725
transform 1 0 27968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1676037725
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1676037725
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_203
timestamp 1676037725
transform 1 0 19780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_215
timestamp 1676037725
transform 1 0 20884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_227
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_239
timestamp 1676037725
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_11
timestamp 1676037725
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1676037725
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1676037725
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_313
timestamp 1676037725
transform 1 0 29900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_318
timestamp 1676037725
transform 1 0 30360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_9
timestamp 1676037725
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1676037725
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1676037725
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1676037725
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1676037725
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_267
timestamp 1676037725
transform 1 0 25668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_290
timestamp 1676037725
transform 1 0 27784 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_302
timestamp 1676037725
transform 1 0 28888 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_314
timestamp 1676037725
transform 1 0 29992 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_326
timestamp 1676037725
transform 1 0 31096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1676037725
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_364
timestamp 1676037725
transform 1 0 34592 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_376
timestamp 1676037725
transform 1 0 35696 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1676037725
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_247
timestamp 1676037725
transform 1 0 23828 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_259
timestamp 1676037725
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1676037725
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_9
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_291
timestamp 1676037725
transform 1 0 27876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1676037725
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1676037725
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_399
timestamp 1676037725
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1676037725
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_225
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_234
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1676037725
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_263
timestamp 1676037725
transform 1 0 25300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_275
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_287
timestamp 1676037725
transform 1 0 27508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_299
timestamp 1676037725
transform 1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1676037725
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1676037725
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1676037725
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1676037725
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_385
timestamp 1676037725
transform 1 0 36524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_397
timestamp 1676037725
transform 1 0 37628 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_409
timestamp 1676037725
transform 1 0 38732 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_417
timestamp 1676037725
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1676037725
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1676037725
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1676037725
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_262
timestamp 1676037725
transform 1 0 25208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_266
timestamp 1676037725
transform 1 0 25576 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_274
timestamp 1676037725
transform 1 0 26312 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1676037725
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_292
timestamp 1676037725
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1676037725
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1676037725
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1676037725
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1676037725
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_245
timestamp 1676037725
transform 1 0 23644 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_257
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1676037725
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_401
timestamp 1676037725
transform 1 0 37996 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_407
timestamp 1676037725
transform 1 0 38548 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_419
timestamp 1676037725
transform 1 0 39652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_431
timestamp 1676037725
transform 1 0 40756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_443
timestamp 1676037725
transform 1 0 41860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_185
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1676037725
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1676037725
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1676037725
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_389
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_395
timestamp 1676037725
transform 1 0 37444 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_400
timestamp 1676037725
transform 1 0 37904 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_412
timestamp 1676037725
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_9
timestamp 1676037725
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_399
timestamp 1676037725
transform 1 0 37812 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_411
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_423
timestamp 1676037725
transform 1 0 40020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_435
timestamp 1676037725
transform 1 0 41124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1676037725
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1676037725
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1676037725
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1676037725
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1676037725
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_23
timestamp 1676037725
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1676037725
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1676037725
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1676037725
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_313
timestamp 1676037725
transform 1 0 29900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_325
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1676037725
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1676037725
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1676037725
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1676037725
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1676037725
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_466
timestamp 1676037725
transform 1 0 43976 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_478
timestamp 1676037725
transform 1 0 45080 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_490
timestamp 1676037725
transform 1 0 46184 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1676037725
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_11
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1676037725
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_294
timestamp 1676037725
transform 1 0 28152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_249
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1676037725
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_401
timestamp 1676037725
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_406
timestamp 1676037725
transform 1 0 38456 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_412
timestamp 1676037725
transform 1 0 39008 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_424
timestamp 1676037725
transform 1 0 40112 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_436
timestamp 1676037725
transform 1 0 41216 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1676037725
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1676037725
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1676037725
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_397
timestamp 1676037725
transform 1 0 37628 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_403
timestamp 1676037725
transform 1 0 38180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_415
timestamp 1676037725
transform 1 0 39284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_465
timestamp 1676037725
transform 1 0 43884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_471
timestamp 1676037725
transform 1 0 44436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_11
timestamp 1676037725
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_23
timestamp 1676037725
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_35
timestamp 1676037725
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1676037725
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1676037725
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1676037725
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1676037725
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1676037725
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1676037725
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1676037725
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1676037725
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1676037725
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1676037725
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1676037725
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1676037725
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1676037725
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1676037725
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1676037725
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_397
timestamp 1676037725
transform 1 0 37628 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_404
timestamp 1676037725
transform 1 0 38272 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1676037725
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1676037725
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1676037725
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1676037725
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1676037725
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1676037725
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1676037725
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1676037725
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1676037725
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_9
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_220
timestamp 1676037725
transform 1 0 21344 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_232
timestamp 1676037725
transform 1 0 22448 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1676037725
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1676037725
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1676037725
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1676037725
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1676037725
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1676037725
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1676037725
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1676037725
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1676037725
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1676037725
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_427
timestamp 1676037725
transform 1 0 40388 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_439
timestamp 1676037725
transform 1 0 41492 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_451
timestamp 1676037725
transform 1 0 42596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_463
timestamp 1676037725
transform 1 0 43700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_184
timestamp 1676037725
transform 1 0 18032 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_196
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_208
timestamp 1676037725
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1676037725
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_231
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_255
timestamp 1676037725
transform 1 0 24564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_267
timestamp 1676037725
transform 1 0 25668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1676037725
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1676037725
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1676037725
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1676037725
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_411
timestamp 1676037725
transform 1 0 38916 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_423
timestamp 1676037725
transform 1 0 40020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_435
timestamp 1676037725
transform 1 0 41124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_469
timestamp 1676037725
transform 1 0 44252 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_474
timestamp 1676037725
transform 1 0 44712 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_486
timestamp 1676037725
transform 1 0 45816 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_498
timestamp 1676037725
transform 1 0 46920 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1676037725
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1676037725
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1676037725
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1676037725
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_23
timestamp 1676037725
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1676037725
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1676037725
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1676037725
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1676037725
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1676037725
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1676037725
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1676037725
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1676037725
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1676037725
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1676037725
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1676037725
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1676037725
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1676037725
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_427
timestamp 1676037725
transform 1 0 40388 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_439
timestamp 1676037725
transform 1 0 41492 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_451
timestamp 1676037725
transform 1 0 42596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_463
timestamp 1676037725
transform 1 0 43700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_11
timestamp 1676037725
transform 1 0 2116 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_23
timestamp 1676037725
transform 1 0 3220 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_35
timestamp 1676037725
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 1676037725
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1676037725
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1676037725
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1676037725
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1676037725
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1676037725
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_399
timestamp 1676037725
transform 1 0 37812 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_411
timestamp 1676037725
transform 1 0 38916 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_423
timestamp 1676037725
transform 1 0 40020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_435
timestamp 1676037725
transform 1 0 41124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_11
timestamp 1676037725
transform 1 0 2116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1676037725
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1676037725
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1676037725
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1676037725
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1676037725
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1676037725
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_463
timestamp 1676037725
transform 1 0 43700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_468
timestamp 1676037725
transform 1 0 44160 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1676037725
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1676037725
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1676037725
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1676037725
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1676037725
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1676037725
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1676037725
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1676037725
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1676037725
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1676037725
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1676037725
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1676037725
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1676037725
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1676037725
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1676037725
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_21
timestamp 1676037725
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_33
timestamp 1676037725
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_45
timestamp 1676037725
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1676037725
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1676037725
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1676037725
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_385
timestamp 1676037725
transform 1 0 36524 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1676037725
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_411
timestamp 1676037725
transform 1 0 38916 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_416
timestamp 1676037725
transform 1 0 39376 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_428
timestamp 1676037725
transform 1 0 40480 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_157
timestamp 1676037725
transform 1 0 15548 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_161
timestamp 1676037725
transform 1 0 15916 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_173
timestamp 1676037725
transform 1 0 17020 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_185
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1676037725
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1676037725
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1676037725
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_398
timestamp 1676037725
transform 1 0 37720 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_410
timestamp 1676037725
transform 1 0 38824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1676037725
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1676037725
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_457
timestamp 1676037725
transform 1 0 43148 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_465
timestamp 1676037725
transform 1 0 43884 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_470
timestamp 1676037725
transform 1 0 44344 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1676037725
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_11
timestamp 1676037725
transform 1 0 2116 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_23
timestamp 1676037725
transform 1 0 3220 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_35
timestamp 1676037725
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1676037725
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1676037725
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1676037725
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1676037725
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1676037725
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1676037725
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1676037725
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_405
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_413
timestamp 1676037725
transform 1 0 39100 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_425
timestamp 1676037725
transform 1 0 40204 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_437
timestamp 1676037725
transform 1 0 41308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1676037725
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_525
timestamp 1676037725
transform 1 0 49404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1676037725
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1676037725
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1676037725
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1676037725
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1676037725
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1676037725
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1676037725
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1676037725
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1676037725
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1676037725
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1676037725
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1676037725
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1676037725
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_501
timestamp 1676037725
transform 1 0 47196 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_525
timestamp 1676037725
transform 1 0 49404 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1676037725
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1676037725
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1676037725
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1676037725
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_404
timestamp 1676037725
transform 1 0 38272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_408
timestamp 1676037725
transform 1 0 38640 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_413
timestamp 1676037725
transform 1 0 39100 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_425
timestamp 1676037725
transform 1 0 40204 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_437
timestamp 1676037725
transform 1 0 41308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_445
timestamp 1676037725
transform 1 0 42044 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1676037725
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1676037725
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1676037725
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1676037725
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_525
timestamp 1676037725
transform 1 0 49404 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_9
timestamp 1676037725
transform 1 0 1932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1676037725
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1676037725
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1676037725
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1676037725
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1676037725
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1676037725
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1676037725
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1676037725
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1676037725
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1676037725
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1676037725
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1676037725
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1676037725
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1676037725
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1676037725
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1676037725
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1676037725
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1676037725
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1676037725
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1676037725
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1676037725
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1676037725
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1676037725
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1676037725
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1676037725
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1676037725
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1676037725
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1676037725
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1676037725
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1676037725
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1676037725
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1676037725
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1676037725
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1676037725
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_469
timestamp 1676037725
transform 1 0 44252 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_475
timestamp 1676037725
transform 1 0 44804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_487
timestamp 1676037725
transform 1 0 45908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_499
timestamp 1676037725
transform 1 0 47012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1676037725
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_525
timestamp 1676037725
transform 1 0 49404 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_164
timestamp 1676037725
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1676037725
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1676037725
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1676037725
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1676037725
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1676037725
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_409
timestamp 1676037725
transform 1 0 38732 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_414
timestamp 1676037725
transform 1 0 39192 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1676037725
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1676037725
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_21
timestamp 1676037725
transform 1 0 3036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_33
timestamp 1676037725
transform 1 0 4140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp 1676037725
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1676037725
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_141
timestamp 1676037725
transform 1 0 14076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_144
timestamp 1676037725
transform 1 0 14352 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_150
timestamp 1676037725
transform 1 0 14904 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1676037725
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_198
timestamp 1676037725
transform 1 0 19320 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_211
timestamp 1676037725
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1676037725
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1676037725
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1676037725
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1676037725
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1676037725
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1676037725
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_477
timestamp 1676037725
transform 1 0 44988 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_482
timestamp 1676037725
transform 1 0 45448 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_494
timestamp 1676037725
transform 1 0 46552 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_502
timestamp 1676037725
transform 1 0 47288 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_521
timestamp 1676037725
transform 1 0 49036 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_525
timestamp 1676037725
transform 1 0 49404 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1676037725
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_164
timestamp 1676037725
transform 1 0 16192 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_172
timestamp 1676037725
transform 1 0 16928 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_211
timestamp 1676037725
transform 1 0 20516 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_224
timestamp 1676037725
transform 1 0 21712 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_236
timestamp 1676037725
transform 1 0 22816 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1676037725
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1676037725
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1676037725
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1676037725
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_394
timestamp 1676037725
transform 1 0 37352 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_406
timestamp 1676037725
transform 1 0 38456 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_418
timestamp 1676037725
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1676037725
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1676037725
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1676037725
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1676037725
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1676037725
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_175
timestamp 1676037725
transform 1 0 17204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_196
timestamp 1676037725
transform 1 0 19136 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1676037725
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_236
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_252
timestamp 1676037725
transform 1 0 24288 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_255
timestamp 1676037725
transform 1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_268
timestamp 1676037725
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_299
timestamp 1676037725
transform 1 0 28612 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_309
timestamp 1676037725
transform 1 0 29532 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_321
timestamp 1676037725
transform 1 0 30636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_333
timestamp 1676037725
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1676037725
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1676037725
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_525
timestamp 1676037725
transform 1 0 49404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1676037725
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_167
timestamp 1676037725
transform 1 0 16468 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1676037725
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_203
timestamp 1676037725
transform 1 0 19780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_227
timestamp 1676037725
transform 1 0 21988 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_234
timestamp 1676037725
transform 1 0 22632 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1676037725
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1676037725
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_314
timestamp 1676037725
transform 1 0 29992 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_326
timestamp 1676037725
transform 1 0 31096 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_338
timestamp 1676037725
transform 1 0 32200 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_350
timestamp 1676037725
transform 1 0 33304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1676037725
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1676037725
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1676037725
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1676037725
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1676037725
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1676037725
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_497
timestamp 1676037725
transform 1 0 46828 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_509
timestamp 1676037725
transform 1 0 47932 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_21
timestamp 1676037725
transform 1 0 3036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_33
timestamp 1676037725
transform 1 0 4140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_45
timestamp 1676037725
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1676037725
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_188
timestamp 1676037725
transform 1 0 18400 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_200
timestamp 1676037725
transform 1 0 19504 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_230
timestamp 1676037725
transform 1 0 22264 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_245
timestamp 1676037725
transform 1 0 23644 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_257
timestamp 1676037725
transform 1 0 24748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_269
timestamp 1676037725
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1676037725
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_301
timestamp 1676037725
transform 1 0 28796 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_307
timestamp 1676037725
transform 1 0 29348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_319
timestamp 1676037725
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1676037725
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_398
timestamp 1676037725
transform 1 0 37720 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_410
timestamp 1676037725
transform 1 0 38824 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_422
timestamp 1676037725
transform 1 0 39928 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_434
timestamp 1676037725
transform 1 0 41032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1676037725
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_525
timestamp 1676037725
transform 1 0 49404 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_125
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_130
timestamp 1676037725
transform 1 0 13064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_154
timestamp 1676037725
transform 1 0 15272 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_183
timestamp 1676037725
transform 1 0 17940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_219
timestamp 1676037725
transform 1 0 21252 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_231
timestamp 1676037725
transform 1 0 22356 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_239
timestamp 1676037725
transform 1 0 23092 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_264
timestamp 1676037725
transform 1 0 25392 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_281
timestamp 1676037725
transform 1 0 26956 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_293
timestamp 1676037725
transform 1 0 28060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1676037725
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1676037725
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1676037725
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1676037725
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1676037725
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1676037725
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1676037725
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_483
timestamp 1676037725
transform 1 0 45540 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_495
timestamp 1676037725
transform 1 0 46644 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_507
timestamp 1676037725
transform 1 0 47748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_519
timestamp 1676037725
transform 1 0 48852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1676037725
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_101
timestamp 1676037725
transform 1 0 10396 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1676037725
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_140
timestamp 1676037725
transform 1 0 13984 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_153
timestamp 1676037725
transform 1 0 15180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_182
timestamp 1676037725
transform 1 0 17848 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_206
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_243
timestamp 1676037725
transform 1 0 23460 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_254
timestamp 1676037725
transform 1 0 24472 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_266
timestamp 1676037725
transform 1 0 25576 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1676037725
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_301
timestamp 1676037725
transform 1 0 28796 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_314
timestamp 1676037725
transform 1 0 29992 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_326
timestamp 1676037725
transform 1 0 31096 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1676037725
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_342
timestamp 1676037725
transform 1 0 32568 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_354
timestamp 1676037725
transform 1 0 33672 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_366
timestamp 1676037725
transform 1 0 34776 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_378
timestamp 1676037725
transform 1 0 35880 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1676037725
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_401
timestamp 1676037725
transform 1 0 37996 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_406
timestamp 1676037725
transform 1 0 38456 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_418
timestamp 1676037725
transform 1 0 39560 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_430
timestamp 1676037725
transform 1 0 40664 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_442
timestamp 1676037725
transform 1 0 41768 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_469
timestamp 1676037725
transform 1 0 44252 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_474
timestamp 1676037725
transform 1 0 44712 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_486
timestamp 1676037725
transform 1 0 45816 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_498
timestamp 1676037725
transform 1 0 46920 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_517
timestamp 1676037725
transform 1 0 48668 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_521
timestamp 1676037725
transform 1 0 49036 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_525
timestamp 1676037725
transform 1 0 49404 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1676037725
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_71
timestamp 1676037725
transform 1 0 7636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_76
timestamp 1676037725
transform 1 0 8096 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_105
timestamp 1676037725
transform 1 0 10764 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_110
timestamp 1676037725
transform 1 0 11224 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_122
timestamp 1676037725
transform 1 0 12328 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 1676037725
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_169
timestamp 1676037725
transform 1 0 16652 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_212
timestamp 1676037725
transform 1 0 20608 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_216
timestamp 1676037725
transform 1 0 20976 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_226
timestamp 1676037725
transform 1 0 21896 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_278
timestamp 1676037725
transform 1 0 26680 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_286
timestamp 1676037725
transform 1 0 27416 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_291
timestamp 1676037725
transform 1 0 27876 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1676037725
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_331
timestamp 1676037725
transform 1 0 31556 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_344
timestamp 1676037725
transform 1 0 32752 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1676037725
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1676037725
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1676037725
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1676037725
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1676037725
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1676037725
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_121
timestamp 1676037725
transform 1 0 12236 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1676037725
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_182
timestamp 1676037725
transform 1 0 17848 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_194
timestamp 1676037725
transform 1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_218
timestamp 1676037725
transform 1 0 21160 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_236
timestamp 1676037725
transform 1 0 22816 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_244
timestamp 1676037725
transform 1 0 23552 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_265
timestamp 1676037725
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1676037725
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_315
timestamp 1676037725
transform 1 0 30084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_328
timestamp 1676037725
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_348
timestamp 1676037725
transform 1 0 33120 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1676037725
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1676037725
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1676037725
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1676037725
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_525
timestamp 1676037725
transform 1 0 49404 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1676037725
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_150
timestamp 1676037725
transform 1 0 14904 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_158
timestamp 1676037725
transform 1 0 15640 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_182
timestamp 1676037725
transform 1 0 17848 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1676037725
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_202
timestamp 1676037725
transform 1 0 19688 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_206
timestamp 1676037725
transform 1 0 20056 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_216
timestamp 1676037725
transform 1 0 20976 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_240
timestamp 1676037725
transform 1 0 23184 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_246
timestamp 1676037725
transform 1 0 23736 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_276
timestamp 1676037725
transform 1 0 26496 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_297
timestamp 1676037725
transform 1 0 28428 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1676037725
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_331
timestamp 1676037725
transform 1 0 31556 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_338
timestamp 1676037725
transform 1 0 32200 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1676037725
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1676037725
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1676037725
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1676037725
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_143
timestamp 1676037725
transform 1 0 14260 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_153
timestamp 1676037725
transform 1 0 15180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1676037725
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_186
timestamp 1676037725
transform 1 0 18216 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_201
timestamp 1676037725
transform 1 0 19596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1676037725
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_251
timestamp 1676037725
transform 1 0 24196 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_272
timestamp 1676037725
transform 1 0 26128 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_303
timestamp 1676037725
transform 1 0 28980 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_310
timestamp 1676037725
transform 1 0 29624 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1676037725
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_342
timestamp 1676037725
transform 1 0 32568 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_346
timestamp 1676037725
transform 1 0 32936 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_367
timestamp 1676037725
transform 1 0 34868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_379
timestamp 1676037725
transform 1 0 35972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_420
timestamp 1676037725
transform 1 0 39744 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_435
timestamp 1676037725
transform 1 0 41124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_525
timestamp 1676037725
transform 1 0 49404 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_152
timestamp 1676037725
transform 1 0 15088 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_176
timestamp 1676037725
transform 1 0 17296 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_184
timestamp 1676037725
transform 1 0 18032 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_225
timestamp 1676037725
transform 1 0 21804 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_240
timestamp 1676037725
transform 1 0 23184 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1676037725
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_271
timestamp 1676037725
transform 1 0 26036 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_283
timestamp 1676037725
transform 1 0 27140 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_289
timestamp 1676037725
transform 1 0 27692 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_302
timestamp 1676037725
transform 1 0 28888 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_320
timestamp 1676037725
transform 1 0 30544 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_341
timestamp 1676037725
transform 1 0 32476 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1676037725
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_370
timestamp 1676037725
transform 1 0 35144 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1676037725
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1676037725
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1676037725
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1676037725
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1676037725
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1676037725
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1676037725
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1676037725
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1676037725
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_129
timestamp 1676037725
transform 1 0 12972 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_139
timestamp 1676037725
transform 1 0 13892 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_152
timestamp 1676037725
transform 1 0 15088 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_156
timestamp 1676037725
transform 1 0 15456 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1676037725
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_175
timestamp 1676037725
transform 1 0 17204 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_191
timestamp 1676037725
transform 1 0 18676 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_215
timestamp 1676037725
transform 1 0 20884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_247
timestamp 1676037725
transform 1 0 23828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1676037725
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_303
timestamp 1676037725
transform 1 0 28980 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_311
timestamp 1676037725
transform 1 0 29716 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1676037725
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_348
timestamp 1676037725
transform 1 0 33120 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_355
timestamp 1676037725
transform 1 0 33764 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_383
timestamp 1676037725
transform 1 0 36340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_408
timestamp 1676037725
transform 1 0 38640 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_420
timestamp 1676037725
transform 1 0 39744 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_432
timestamp 1676037725
transform 1 0 40848 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_438
timestamp 1676037725
transform 1 0 41400 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1676037725
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1676037725
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1676037725
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1676037725
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1676037725
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1676037725
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_521
timestamp 1676037725
transform 1 0 49036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_525
timestamp 1676037725
transform 1 0 49404 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1676037725
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_117
timestamp 1676037725
transform 1 0 11868 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_163
timestamp 1676037725
transform 1 0 16100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_178
timestamp 1676037725
transform 1 0 17480 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1676037725
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_208
timestamp 1676037725
transform 1 0 20240 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_232
timestamp 1676037725
transform 1 0 22448 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_240
timestamp 1676037725
transform 1 0 23184 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1676037725
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_276
timestamp 1676037725
transform 1 0 26496 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_284
timestamp 1676037725
transform 1 0 27232 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_296
timestamp 1676037725
transform 1 0 28336 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_300
timestamp 1676037725
transform 1 0 28704 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1676037725
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_320
timestamp 1676037725
transform 1 0 30544 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_333
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_346
timestamp 1676037725
transform 1 0 32936 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_350
timestamp 1676037725
transform 1 0 33304 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1676037725
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_387
timestamp 1676037725
transform 1 0 36708 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_399
timestamp 1676037725
transform 1 0 37812 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_411
timestamp 1676037725
transform 1 0 38916 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_426
timestamp 1676037725
transform 1 0 40296 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_438
timestamp 1676037725
transform 1 0 41400 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_450
timestamp 1676037725
transform 1 0 42504 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_462
timestamp 1676037725
transform 1 0 43608 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_474
timestamp 1676037725
transform 1 0 44712 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_94
timestamp 1676037725
transform 1 0 9752 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_106
timestamp 1676037725
transform 1 0 10856 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_129
timestamp 1676037725
transform 1 0 12972 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_150
timestamp 1676037725
transform 1 0 14904 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1676037725
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_175
timestamp 1676037725
transform 1 0 17204 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_178
timestamp 1676037725
transform 1 0 17480 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_191
timestamp 1676037725
transform 1 0 18676 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1676037725
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1676037725
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_230
timestamp 1676037725
transform 1 0 22264 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_245
timestamp 1676037725
transform 1 0 23644 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_249
timestamp 1676037725
transform 1 0 24012 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_270
timestamp 1676037725
transform 1 0 25944 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1676037725
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_293
timestamp 1676037725
transform 1 0 28060 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_315
timestamp 1676037725
transform 1 0 30084 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 1676037725
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_350
timestamp 1676037725
transform 1 0 33304 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_358
timestamp 1676037725
transform 1 0 34040 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_379
timestamp 1676037725
transform 1 0 35972 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1676037725
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_404
timestamp 1676037725
transform 1 0 38272 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_416
timestamp 1676037725
transform 1 0 39376 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_428
timestamp 1676037725
transform 1 0 40480 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_440
timestamp 1676037725
transform 1 0 41584 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_525
timestamp 1676037725
transform 1 0 49404 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1676037725
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1676037725
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_96
timestamp 1676037725
transform 1 0 9936 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_108
timestamp 1676037725
transform 1 0 11040 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_116
timestamp 1676037725
transform 1 0 11776 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1676037725
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1676037725
transform 1 0 14444 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_155
timestamp 1676037725
transform 1 0 15364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_175
timestamp 1676037725
transform 1 0 17204 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_181
timestamp 1676037725
transform 1 0 17756 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_219
timestamp 1676037725
transform 1 0 21252 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_227
timestamp 1676037725
transform 1 0 21988 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_275
timestamp 1676037725
transform 1 0 26404 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_283
timestamp 1676037725
transform 1 0 27140 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1676037725
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_313
timestamp 1676037725
transform 1 0 29900 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_334
timestamp 1676037725
transform 1 0 31832 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_347
timestamp 1676037725
transform 1 0 33028 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1676037725
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_388
timestamp 1676037725
transform 1 0 36800 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_412
timestamp 1676037725
transform 1 0 39008 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1676037725
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1676037725
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1676037725
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1676037725
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_121
timestamp 1676037725
transform 1 0 12236 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1676037725
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_155
timestamp 1676037725
transform 1 0 15364 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1676037725
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_191
timestamp 1676037725
transform 1 0 18676 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_204
timestamp 1676037725
transform 1 0 19872 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_212
timestamp 1676037725
transform 1 0 20608 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1676037725
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_236
timestamp 1676037725
transform 1 0 22816 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1676037725
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_306
timestamp 1676037725
transform 1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_331
timestamp 1676037725
transform 1 0 31556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_360
timestamp 1676037725
transform 1 0 34224 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1676037725
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_401
timestamp 1676037725
transform 1 0 37996 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_413
timestamp 1676037725
transform 1 0 39100 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_425
timestamp 1676037725
transform 1 0 40204 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_437
timestamp 1676037725
transform 1 0 41308 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_445
timestamp 1676037725
transform 1 0 42044 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_525
timestamp 1676037725
transform 1 0 49404 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1676037725
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_154
timestamp 1676037725
transform 1 0 15272 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_180
timestamp 1676037725
transform 1 0 17664 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1676037725
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_201
timestamp 1676037725
transform 1 0 19596 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_211
timestamp 1676037725
transform 1 0 20516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_218
timestamp 1676037725
transform 1 0 21160 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1676037725
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_246
timestamp 1676037725
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_282
timestamp 1676037725
transform 1 0 27048 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_297
timestamp 1676037725
transform 1 0 28428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1676037725
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_341
timestamp 1676037725
transform 1 0 32476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_354
timestamp 1676037725
transform 1 0 33672 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1676037725
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_371
timestamp 1676037725
transform 1 0 35236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_392
timestamp 1676037725
transform 1 0 37168 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_405
timestamp 1676037725
transform 1 0 38364 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1676037725
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_21
timestamp 1676037725
transform 1 0 3036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_33
timestamp 1676037725
transform 1 0 4140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_45
timestamp 1676037725
transform 1 0 5244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_53
timestamp 1676037725
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_77
timestamp 1676037725
transform 1 0 8188 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_83
timestamp 1676037725
transform 1 0 8740 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_95
timestamp 1676037725
transform 1 0 9844 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_107
timestamp 1676037725
transform 1 0 10948 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_130
timestamp 1676037725
transform 1 0 13064 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_142
timestamp 1676037725
transform 1 0 14168 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_175
timestamp 1676037725
transform 1 0 17204 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_179
timestamp 1676037725
transform 1 0 17572 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_192
timestamp 1676037725
transform 1 0 18768 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_203
timestamp 1676037725
transform 1 0 19780 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_209
timestamp 1676037725
transform 1 0 20332 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1676037725
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_250
timestamp 1676037725
transform 1 0 24104 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_263
timestamp 1676037725
transform 1 0 25300 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1676037725
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_303
timestamp 1676037725
transform 1 0 28980 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1676037725
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_367
timestamp 1676037725
transform 1 0 34868 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_380
timestamp 1676037725
transform 1 0 36064 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_404
timestamp 1676037725
transform 1 0 38272 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_521
timestamp 1676037725
transform 1 0 49036 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_525
timestamp 1676037725
transform 1 0 49404 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp 1676037725
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_81
timestamp 1676037725
transform 1 0 8556 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_132
timestamp 1676037725
transform 1 0 13248 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_173
timestamp 1676037725
transform 1 0 17020 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_179
timestamp 1676037725
transform 1 0 17572 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1676037725
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_224
timestamp 1676037725
transform 1 0 21712 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_237
timestamp 1676037725
transform 1 0 22908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1676037725
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_270
timestamp 1676037725
transform 1 0 25944 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_276
timestamp 1676037725
transform 1 0 26496 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_291
timestamp 1676037725
transform 1 0 27876 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1676037725
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_331
timestamp 1676037725
transform 1 0 31556 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_335
timestamp 1676037725
transform 1 0 31924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_339
timestamp 1676037725
transform 1 0 32292 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_356
timestamp 1676037725
transform 1 0 33856 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_378
timestamp 1676037725
transform 1 0 35880 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_391
timestamp 1676037725
transform 1 0 37076 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_152
timestamp 1676037725
transform 1 0 15088 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_165
timestamp 1676037725
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_192
timestamp 1676037725
transform 1 0 18768 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_200
timestamp 1676037725
transform 1 0 19504 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1676037725
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_247
timestamp 1676037725
transform 1 0 23828 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_260
timestamp 1676037725
transform 1 0 25024 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_267
timestamp 1676037725
transform 1 0 25668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1676037725
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_292
timestamp 1676037725
transform 1 0 27968 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_296
timestamp 1676037725
transform 1 0 28336 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_334
timestamp 1676037725
transform 1 0 31832 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_343
timestamp 1676037725
transform 1 0 32660 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_353
timestamp 1676037725
transform 1 0 33580 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_366
timestamp 1676037725
transform 1 0 34776 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1676037725
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_401
timestamp 1676037725
transform 1 0 37996 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_404
timestamp 1676037725
transform 1 0 38272 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_525
timestamp 1676037725
transform 1 0 49404 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1676037725
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_103
timestamp 1676037725
transform 1 0 10580 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_127
timestamp 1676037725
transform 1 0 12788 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_135
timestamp 1676037725
transform 1 0 13524 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_147
timestamp 1676037725
transform 1 0 14628 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_151
timestamp 1676037725
transform 1 0 14996 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_157
timestamp 1676037725
transform 1 0 15548 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_178
timestamp 1676037725
transform 1 0 17480 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_184
timestamp 1676037725
transform 1 0 18032 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1676037725
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_201
timestamp 1676037725
transform 1 0 19596 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_211
timestamp 1676037725
transform 1 0 20516 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_224
timestamp 1676037725
transform 1 0 21712 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_237
timestamp 1676037725
transform 1 0 22908 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1676037725
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_281
timestamp 1676037725
transform 1 0 26956 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1676037725
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_320
timestamp 1676037725
transform 1 0 30544 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_349
timestamp 1676037725
transform 1 0 33212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_362
timestamp 1676037725
transform 1 0 34408 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_391
timestamp 1676037725
transform 1 0 37076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_397
timestamp 1676037725
transform 1 0 37628 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1676037725
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1676037725
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1676037725
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1676037725
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_21
timestamp 1676037725
transform 1 0 3036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_33
timestamp 1676037725
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_45
timestamp 1676037725
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_53
timestamp 1676037725
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_152
timestamp 1676037725
transform 1 0 15088 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_158
timestamp 1676037725
transform 1 0 15640 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_166
timestamp 1676037725
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_177
timestamp 1676037725
transform 1 0 17388 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_194
timestamp 1676037725
transform 1 0 18952 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_200
timestamp 1676037725
transform 1 0 19504 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1676037725
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_229
timestamp 1676037725
transform 1 0 22172 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_239
timestamp 1676037725
transform 1 0 23092 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_252
timestamp 1676037725
transform 1 0 24288 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_275
timestamp 1676037725
transform 1 0 26404 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_292
timestamp 1676037725
transform 1 0 27968 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_318
timestamp 1676037725
transform 1 0 30360 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_324
timestamp 1676037725
transform 1 0 30912 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 1676037725
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_359
timestamp 1676037725
transform 1 0 34132 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_383
timestamp 1676037725
transform 1 0 36340 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_401
timestamp 1676037725
transform 1 0 37996 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_404
timestamp 1676037725
transform 1 0 38272 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1676037725
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1676037725
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1676037725
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1676037725
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_517
timestamp 1676037725
transform 1 0 48668 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_525
timestamp 1676037725
transform 1 0 49404 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_117
timestamp 1676037725
transform 1 0 11868 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_123
timestamp 1676037725
transform 1 0 12420 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_129
timestamp 1676037725
transform 1 0 12972 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_159
timestamp 1676037725
transform 1 0 15732 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_183
timestamp 1676037725
transform 1 0 17940 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_191
timestamp 1676037725
transform 1 0 18676 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_208
timestamp 1676037725
transform 1 0 20240 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_235
timestamp 1676037725
transform 1 0 22724 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1676037725
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_261
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_265
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_275
timestamp 1676037725
transform 1 0 26404 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_288
timestamp 1676037725
transform 1 0 27600 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_292
timestamp 1676037725
transform 1 0 27968 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_302
timestamp 1676037725
transform 1 0 28888 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_320
timestamp 1676037725
transform 1 0 30544 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_333
timestamp 1676037725
transform 1 0 31740 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_339
timestamp 1676037725
transform 1 0 32292 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_351
timestamp 1676037725
transform 1 0 33396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1676037725
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_369
timestamp 1676037725
transform 1 0 35052 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_393
timestamp 1676037725
transform 1 0 37260 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_399
timestamp 1676037725
transform 1 0 37812 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_412
timestamp 1676037725
transform 1 0 39008 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1676037725
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1676037725
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1676037725
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_121
timestamp 1676037725
transform 1 0 12236 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_126
timestamp 1676037725
transform 1 0 12696 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_134
timestamp 1676037725
transform 1 0 13432 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_146
timestamp 1676037725
transform 1 0 14536 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_157
timestamp 1676037725
transform 1 0 15548 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_165
timestamp 1676037725
transform 1 0 16284 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_189
timestamp 1676037725
transform 1 0 18492 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_213
timestamp 1676037725
transform 1 0 20700 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1676037725
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_240
timestamp 1676037725
transform 1 0 23184 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_253
timestamp 1676037725
transform 1 0 24380 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_266
timestamp 1676037725
transform 1 0 25576 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1676037725
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_298
timestamp 1676037725
transform 1 0 28520 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_304
timestamp 1676037725
transform 1 0 29072 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_314
timestamp 1676037725
transform 1 0 29992 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_326
timestamp 1676037725
transform 1 0 31096 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_332
timestamp 1676037725
transform 1 0 31648 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_348
timestamp 1676037725
transform 1 0 33120 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_377
timestamp 1676037725
transform 1 0 35788 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_389
timestamp 1676037725
transform 1 0 36892 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_415
timestamp 1676037725
transform 1 0 39284 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_427
timestamp 1676037725
transform 1 0 40388 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_439
timestamp 1676037725
transform 1 0 41492 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_517
timestamp 1676037725
transform 1 0 48668 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_521
timestamp 1676037725
transform 1 0 49036 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_525
timestamp 1676037725
transform 1 0 49404 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1676037725
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_117
timestamp 1676037725
transform 1 0 11868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_129
timestamp 1676037725
transform 1 0 12972 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_149
timestamp 1676037725
transform 1 0 14812 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_160
timestamp 1676037725
transform 1 0 15824 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_167
timestamp 1676037725
transform 1 0 16468 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_176
timestamp 1676037725
transform 1 0 17296 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_188
timestamp 1676037725
transform 1 0 18400 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1676037725
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_208
timestamp 1676037725
transform 1 0 20240 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_223
timestamp 1676037725
transform 1 0 21620 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_278
timestamp 1676037725
transform 1 0 26680 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_284
timestamp 1676037725
transform 1 0 27232 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_297
timestamp 1676037725
transform 1 0 28428 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1676037725
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_331
timestamp 1676037725
transform 1 0 31556 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_355
timestamp 1676037725
transform 1 0 33764 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_387
timestamp 1676037725
transform 1 0 36708 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_399
timestamp 1676037725
transform 1 0 37812 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_411
timestamp 1676037725
transform 1 0 38916 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_119
timestamp 1676037725
transform 1 0 12052 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_131
timestamp 1676037725
transform 1 0 13156 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_143
timestamp 1676037725
transform 1 0 14260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_155
timestamp 1676037725
transform 1 0 15364 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_166
timestamp 1676037725
transform 1 0 16376 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_191
timestamp 1676037725
transform 1 0 18676 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_214
timestamp 1676037725
transform 1 0 20792 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_221
timestamp 1676037725
transform 1 0 21436 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_247
timestamp 1676037725
transform 1 0 23828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1676037725
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_294
timestamp 1676037725
transform 1 0 28152 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_309
timestamp 1676037725
transform 1 0 29532 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1676037725
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_370
timestamp 1676037725
transform 1 0 35144 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_378
timestamp 1676037725
transform 1 0 35880 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 1676037725
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_404
timestamp 1676037725
transform 1 0 38272 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_416
timestamp 1676037725
transform 1 0 39376 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_428
timestamp 1676037725
transform 1 0 40480 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_440
timestamp 1676037725
transform 1 0 41584 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_517
timestamp 1676037725
transform 1 0 48668 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_525
timestamp 1676037725
transform 1 0 49404 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_21
timestamp 1676037725
transform 1 0 3036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_149
timestamp 1676037725
transform 1 0 14812 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_155
timestamp 1676037725
transform 1 0 15364 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_167
timestamp 1676037725
transform 1 0 16468 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_174
timestamp 1676037725
transform 1 0 17112 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_181
timestamp 1676037725
transform 1 0 17756 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_194
timestamp 1676037725
transform 1 0 18952 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_202
timestamp 1676037725
transform 1 0 19688 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_228
timestamp 1676037725
transform 1 0 22080 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_243
timestamp 1676037725
transform 1 0 23460 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_264
timestamp 1676037725
transform 1 0 25392 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_271
timestamp 1676037725
transform 1 0 26036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_277
timestamp 1676037725
transform 1 0 26588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_281
timestamp 1676037725
transform 1 0 26956 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_285
timestamp 1676037725
transform 1 0 27324 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1676037725
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_322
timestamp 1676037725
transform 1 0 30728 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_346
timestamp 1676037725
transform 1 0 32936 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1676037725
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_369
timestamp 1676037725
transform 1 0 35052 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_390
timestamp 1676037725
transform 1 0 36984 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_402
timestamp 1676037725
transform 1 0 38088 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_414
timestamp 1676037725
transform 1 0 39192 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1676037725
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1676037725
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1676037725
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1676037725
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1676037725
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1676037725
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1676037725
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_45
timestamp 1676037725
transform 1 0 5244 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_77
timestamp 1676037725
transform 1 0 8188 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_84
timestamp 1676037725
transform 1 0 8832 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_96
timestamp 1676037725
transform 1 0 9936 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_108
timestamp 1676037725
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1676037725
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_198
timestamp 1676037725
transform 1 0 19320 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_222
timestamp 1676037725
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_231
timestamp 1676037725
transform 1 0 22356 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_252
timestamp 1676037725
transform 1 0 24288 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1676037725
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_286
timestamp 1676037725
transform 1 0 27416 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_298
timestamp 1676037725
transform 1 0 28520 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_306
timestamp 1676037725
transform 1 0 29256 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_328
timestamp 1676037725
transform 1 0 31280 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_359
timestamp 1676037725
transform 1 0 34132 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_370
timestamp 1676037725
transform 1 0 35144 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_383
timestamp 1676037725
transform 1 0 36340 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1676037725
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1676037725
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1676037725
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_517
timestamp 1676037725
transform 1 0 48668 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_525
timestamp 1676037725
transform 1 0 49404 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_35
timestamp 1676037725
transform 1 0 4324 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_40
timestamp 1676037725
transform 1 0 4784 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_46
timestamp 1676037725
transform 1 0 5336 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_51
timestamp 1676037725
transform 1 0 5796 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_63
timestamp 1676037725
transform 1 0 6900 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_75
timestamp 1676037725
transform 1 0 8004 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_117
timestamp 1676037725
transform 1 0 11868 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_122
timestamp 1676037725
transform 1 0 12328 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_130
timestamp 1676037725
transform 1 0 13064 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_138
timestamp 1676037725
transform 1 0 13800 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_159
timestamp 1676037725
transform 1 0 15732 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_166
timestamp 1676037725
transform 1 0 16376 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1676037725
transform 1 0 18952 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_232
timestamp 1676037725
transform 1 0 22448 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_257
timestamp 1676037725
transform 1 0 24748 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_278
timestamp 1676037725
transform 1 0 26680 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_290
timestamp 1676037725
transform 1 0 27784 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1676037725
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1676037725
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_320
timestamp 1676037725
transform 1 0 30544 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_349
timestamp 1676037725
transform 1 0 33212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1676037725
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1676037725
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1676037725
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1676037725
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1676037725
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1676037725
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_21
timestamp 1676037725
transform 1 0 3036 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_32
timestamp 1676037725
transform 1 0 4048 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_44
timestamp 1676037725
transform 1 0 5152 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_49
timestamp 1676037725
transform 1 0 5612 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_65
timestamp 1676037725
transform 1 0 7084 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_77
timestamp 1676037725
transform 1 0 8188 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_89
timestamp 1676037725
transform 1 0 9292 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_97
timestamp 1676037725
transform 1 0 10028 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_102
timestamp 1676037725
transform 1 0 10488 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1676037725
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_155
timestamp 1676037725
transform 1 0 15364 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_159
timestamp 1676037725
transform 1 0 15732 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_166
timestamp 1676037725
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_184
timestamp 1676037725
transform 1 0 18032 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_208
timestamp 1676037725
transform 1 0 20240 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_212
timestamp 1676037725
transform 1 0 20608 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_222
timestamp 1676037725
transform 1 0 21528 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_236
timestamp 1676037725
transform 1 0 22816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_240
timestamp 1676037725
transform 1 0 23184 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_262
timestamp 1676037725
transform 1 0 25208 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_269
timestamp 1676037725
transform 1 0 25852 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_277
timestamp 1676037725
transform 1 0 26588 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_292
timestamp 1676037725
transform 1 0 27968 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_320
timestamp 1676037725
transform 1 0 30544 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_333
timestamp 1676037725
transform 1 0 31740 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_341
timestamp 1676037725
transform 1 0 32476 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_351
timestamp 1676037725
transform 1 0 33396 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_364
timestamp 1676037725
transform 1 0 34592 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_386
timestamp 1676037725
transform 1 0 36616 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_404
timestamp 1676037725
transform 1 0 38272 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_416
timestamp 1676037725
transform 1 0 39376 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_428
timestamp 1676037725
transform 1 0 40480 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_440
timestamp 1676037725
transform 1 0 41584 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_521
timestamp 1676037725
transform 1 0 49036 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_525
timestamp 1676037725
transform 1 0 49404 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_21
timestamp 1676037725
transform 1 0 3036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_69
timestamp 1676037725
transform 1 0 7452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_81
timestamp 1676037725
transform 1 0 8556 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_125
timestamp 1676037725
transform 1 0 12604 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_129
timestamp 1676037725
transform 1 0 12972 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_137
timestamp 1676037725
transform 1 0 13708 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1676037725
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_203
timestamp 1676037725
transform 1 0 19780 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_225
timestamp 1676037725
transform 1 0 21804 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_232
timestamp 1676037725
transform 1 0 22448 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_240
timestamp 1676037725
transform 1 0 23184 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1676037725
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_275
timestamp 1676037725
transform 1 0 26404 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_288
timestamp 1676037725
transform 1 0 27600 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_295
timestamp 1676037725
transform 1 0 28244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_302
timestamp 1676037725
transform 1 0 28888 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_320
timestamp 1676037725
transform 1 0 30544 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_324
timestamp 1676037725
transform 1 0 30912 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_334
timestamp 1676037725
transform 1 0 31832 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_342
timestamp 1676037725
transform 1 0 32568 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_353
timestamp 1676037725
transform 1 0 33580 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_360
timestamp 1676037725
transform 1 0 34224 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_414
timestamp 1676037725
transform 1 0 39192 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_65
timestamp 1676037725
transform 1 0 7084 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_72
timestamp 1676037725
transform 1 0 7728 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_84
timestamp 1676037725
transform 1 0 8832 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_96
timestamp 1676037725
transform 1 0 9936 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_108
timestamp 1676037725
transform 1 0 11040 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_117
timestamp 1676037725
transform 1 0 11868 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_121
timestamp 1676037725
transform 1 0 12236 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_129
timestamp 1676037725
transform 1 0 12972 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_134
timestamp 1676037725
transform 1 0 13432 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_146
timestamp 1676037725
transform 1 0 14536 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_158
timestamp 1676037725
transform 1 0 15640 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_166
timestamp 1676037725
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_187
timestamp 1676037725
transform 1 0 18308 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_194
timestamp 1676037725
transform 1 0 18952 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_222
timestamp 1676037725
transform 1 0 21528 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_229
timestamp 1676037725
transform 1 0 22172 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_239
timestamp 1676037725
transform 1 0 23092 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_252
timestamp 1676037725
transform 1 0 24288 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_265
timestamp 1676037725
transform 1 0 25484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1676037725
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_292
timestamp 1676037725
transform 1 0 27968 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_320
timestamp 1676037725
transform 1 0 30544 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_324
timestamp 1676037725
transform 1 0 30912 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1676037725
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_341
timestamp 1676037725
transform 1 0 32476 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_351
timestamp 1676037725
transform 1 0 33396 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_364
timestamp 1676037725
transform 1 0 34592 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_372
timestamp 1676037725
transform 1 0 35328 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_377
timestamp 1676037725
transform 1 0 35788 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_390
timestamp 1676037725
transform 1 0 36984 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_404
timestamp 1676037725
transform 1 0 38272 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_412
timestamp 1676037725
transform 1 0 39008 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_423
timestamp 1676037725
transform 1 0 40020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_435
timestamp 1676037725
transform 1 0 41124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1676037725
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_517
timestamp 1676037725
transform 1 0 48668 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_525
timestamp 1676037725
transform 1 0 49404 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_105
timestamp 1676037725
transform 1 0 10764 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_110
timestamp 1676037725
transform 1 0 11224 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_122
timestamp 1676037725
transform 1 0 12328 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_134
timestamp 1676037725
transform 1 0 13432 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1676037725
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_202
timestamp 1676037725
transform 1 0 19688 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_210
timestamp 1676037725
transform 1 0 20424 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_220
timestamp 1676037725
transform 1 0 21344 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_244
timestamp 1676037725
transform 1 0 23552 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_259
timestamp 1676037725
transform 1 0 24932 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_269
timestamp 1676037725
transform 1 0 25852 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_282
timestamp 1676037725
transform 1 0 27048 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1676037725
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_313
timestamp 1676037725
transform 1 0 29900 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_323
timestamp 1676037725
transform 1 0 30820 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_334
timestamp 1676037725
transform 1 0 31832 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_340
timestamp 1676037725
transform 1 0 32384 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_353
timestamp 1676037725
transform 1 0 33580 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1676037725
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_369
timestamp 1676037725
transform 1 0 35052 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_391
timestamp 1676037725
transform 1 0 37076 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_404
timestamp 1676037725
transform 1 0 38272 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_416
timestamp 1676037725
transform 1 0 39376 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_513
timestamp 1676037725
transform 1 0 48300 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_21
timestamp 1676037725
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_33
timestamp 1676037725
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_45
timestamp 1676037725
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1676037725
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_117
timestamp 1676037725
transform 1 0 11868 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_121
timestamp 1676037725
transform 1 0 12236 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_133
timestamp 1676037725
transform 1 0 13340 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_145
timestamp 1676037725
transform 1 0 14444 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_157
timestamp 1676037725
transform 1 0 15548 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_165
timestamp 1676037725
transform 1 0 16284 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_201
timestamp 1676037725
transform 1 0 19596 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1676037725
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_248
timestamp 1676037725
transform 1 0 23920 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_256
timestamp 1676037725
transform 1 0 24656 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1676037725
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_296
timestamp 1676037725
transform 1 0 28336 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_300
timestamp 1676037725
transform 1 0 28704 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_310
timestamp 1676037725
transform 1 0 29624 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_334
timestamp 1676037725
transform 1 0 31832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_348
timestamp 1676037725
transform 1 0 33120 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_360
timestamp 1676037725
transform 1 0 34224 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_383
timestamp 1676037725
transform 1 0 36340 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_525
timestamp 1676037725
transform 1 0 49404 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1676037725
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_203
timestamp 1676037725
transform 1 0 19780 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_207
timestamp 1676037725
transform 1 0 20148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_220
timestamp 1676037725
transform 1 0 21344 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_228
timestamp 1676037725
transform 1 0 22080 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1676037725
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_268
timestamp 1676037725
transform 1 0 25760 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_292
timestamp 1676037725
transform 1 0 27968 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1676037725
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_320
timestamp 1676037725
transform 1 0 30544 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_346
timestamp 1676037725
transform 1 0 32936 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_359
timestamp 1676037725
transform 1 0 34132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_376
timestamp 1676037725
transform 1 0 35696 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_405
timestamp 1676037725
transform 1 0 38364 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_415
timestamp 1676037725
transform 1 0 39284 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1676037725
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1676037725
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1676037725
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1676037725
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_124
timestamp 1676037725
transform 1 0 12512 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_136
timestamp 1676037725
transform 1 0 13616 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_148
timestamp 1676037725
transform 1 0 14720 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_160
timestamp 1676037725
transform 1 0 15824 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_201
timestamp 1676037725
transform 1 0 19596 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_222
timestamp 1676037725
transform 1 0 21528 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_236
timestamp 1676037725
transform 1 0 22816 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_260
timestamp 1676037725
transform 1 0 25024 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1676037725
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1676037725
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_292
timestamp 1676037725
transform 1 0 27968 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_304
timestamp 1676037725
transform 1 0 29072 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_328
timestamp 1676037725
transform 1 0 31280 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_345
timestamp 1676037725
transform 1 0 32844 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_366
timestamp 1676037725
transform 1 0 34776 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_379
timestamp 1676037725
transform 1 0 35972 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_401
timestamp 1676037725
transform 1 0 37996 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_413
timestamp 1676037725
transform 1 0 39100 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_425
timestamp 1676037725
transform 1 0 40204 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_437
timestamp 1676037725
transform 1 0 41308 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_445
timestamp 1676037725
transform 1 0 42044 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_521
timestamp 1676037725
transform 1 0 49036 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_525
timestamp 1676037725
transform 1 0 49404 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1676037725
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_201
timestamp 1676037725
transform 1 0 19596 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_211
timestamp 1676037725
transform 1 0 20516 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_219
timestamp 1676037725
transform 1 0 21252 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_225
timestamp 1676037725
transform 1 0 21804 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_229
timestamp 1676037725
transform 1 0 22172 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_250
timestamp 1676037725
transform 1 0 24104 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_281
timestamp 1676037725
transform 1 0 26956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_302
timestamp 1676037725
transform 1 0 28888 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_343
timestamp 1676037725
transform 1 0 32660 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_356
timestamp 1676037725
transform 1 0 33856 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_376
timestamp 1676037725
transform 1 0 35696 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_391
timestamp 1676037725
transform 1 0 37076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_403
timestamp 1676037725
transform 1 0 38180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_415
timestamp 1676037725
transform 1 0 39284 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_521
timestamp 1676037725
transform 1 0 49036 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_245
timestamp 1676037725
transform 1 0 23644 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_255
timestamp 1676037725
transform 1 0 24564 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_265
timestamp 1676037725
transform 1 0 25484 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_278
timestamp 1676037725
transform 1 0 26680 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_292
timestamp 1676037725
transform 1 0 27968 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_304
timestamp 1676037725
transform 1 0 29072 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_314
timestamp 1676037725
transform 1 0 29992 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_327
timestamp 1676037725
transform 1 0 31188 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_360
timestamp 1676037725
transform 1 0 34224 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_525
timestamp 1676037725
transform 1 0 49404 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_93
timestamp 1676037725
transform 1 0 9660 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_99
timestamp 1676037725
transform 1 0 10212 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_111
timestamp 1676037725
transform 1 0 11316 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_123
timestamp 1676037725
transform 1 0 12420 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_131
timestamp 1676037725
transform 1 0 13156 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_136
timestamp 1676037725
transform 1 0 13616 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_207
timestamp 1676037725
transform 1 0 20148 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_219
timestamp 1676037725
transform 1 0 21252 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_231
timestamp 1676037725
transform 1 0 22356 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_243
timestamp 1676037725
transform 1 0 23460 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_261
timestamp 1676037725
transform 1 0 25116 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_284
timestamp 1676037725
transform 1 0 27232 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_297
timestamp 1676037725
transform 1 0 28428 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1676037725
transform 1 0 29072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_320
timestamp 1676037725
transform 1 0 30544 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_332
timestamp 1676037725
transform 1 0 31648 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_353
timestamp 1676037725
transform 1 0 33580 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_361
timestamp 1676037725
transform 1 0 34316 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_376
timestamp 1676037725
transform 1 0 35696 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_388
timestamp 1676037725
transform 1 0 36800 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_400
timestamp 1676037725
transform 1 0 37904 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_412
timestamp 1676037725
transform 1 0 39008 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_21
timestamp 1676037725
transform 1 0 3036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_33
timestamp 1676037725
transform 1 0 4140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_45
timestamp 1676037725
transform 1 0 5244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1676037725
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_131
timestamp 1676037725
transform 1 0 13156 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_135
timestamp 1676037725
transform 1 0 13524 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_143
timestamp 1676037725
transform 1 0 14260 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_87_153
timestamp 1676037725
transform 1 0 15180 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_166
timestamp 1676037725
transform 1 0 16376 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_222
timestamp 1676037725
transform 1 0 21528 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_231
timestamp 1676037725
transform 1 0 22356 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_243
timestamp 1676037725
transform 1 0 23460 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_255
timestamp 1676037725
transform 1 0 24564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_267
timestamp 1676037725
transform 1 0 25668 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_287
timestamp 1676037725
transform 1 0 27508 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_308
timestamp 1676037725
transform 1 0 29440 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_321
timestamp 1676037725
transform 1 0 30636 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_334
timestamp 1676037725
transform 1 0 31832 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_348
timestamp 1676037725
transform 1 0 33120 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_374
timestamp 1676037725
transform 1 0 35512 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_386
timestamp 1676037725
transform 1 0 36616 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_521
timestamp 1676037725
transform 1 0 49036 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_525
timestamp 1676037725
transform 1 0 49404 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_73
timestamp 1676037725
transform 1 0 7820 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_80
timestamp 1676037725
transform 1 0 8464 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_129
timestamp 1676037725
transform 1 0 12972 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_136
timestamp 1676037725
transform 1 0 13616 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_173
timestamp 1676037725
transform 1 0 17020 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_181
timestamp 1676037725
transform 1 0 17756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_193
timestamp 1676037725
transform 1 0 18860 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_229
timestamp 1676037725
transform 1 0 22172 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_236
timestamp 1676037725
transform 1 0 22816 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_248
timestamp 1676037725
transform 1 0 23920 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_299
timestamp 1676037725
transform 1 0 28612 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_322
timestamp 1676037725
transform 1 0 30728 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_335
timestamp 1676037725
transform 1 0 31924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_347
timestamp 1676037725
transform 1 0 33028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_359
timestamp 1676037725
transform 1 0 34132 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_21
timestamp 1676037725
transform 1 0 3036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_33
timestamp 1676037725
transform 1 0 4140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_45
timestamp 1676037725
transform 1 0 5244 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_53
timestamp 1676037725
transform 1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_91
timestamp 1676037725
transform 1 0 9476 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_95
timestamp 1676037725
transform 1 0 9844 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_100
timestamp 1676037725
transform 1 0 10304 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_131
timestamp 1676037725
transform 1 0 13156 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_136
timestamp 1676037725
transform 1 0 13616 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_148
timestamp 1676037725
transform 1 0 14720 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_160
timestamp 1676037725
transform 1 0 15824 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_175
timestamp 1676037725
transform 1 0 17204 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_187
timestamp 1676037725
transform 1 0 18308 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_199
timestamp 1676037725
transform 1 0 19412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_211
timestamp 1676037725
transform 1 0 20516 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_231
timestamp 1676037725
transform 1 0 22356 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_243
timestamp 1676037725
transform 1 0 23460 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_255
timestamp 1676037725
transform 1 0 24564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_267
timestamp 1676037725
transform 1 0 25668 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_276
timestamp 1676037725
transform 1 0 26496 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_288
timestamp 1676037725
transform 1 0 27600 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_292
timestamp 1676037725
transform 1 0 27968 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_296
timestamp 1676037725
transform 1 0 28336 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_308
timestamp 1676037725
transform 1 0 29440 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_320
timestamp 1676037725
transform 1 0 30544 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_324
timestamp 1676037725
transform 1 0 30912 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_334
timestamp 1676037725
transform 1 0 31832 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_521
timestamp 1676037725
transform 1 0 49036 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_525
timestamp 1676037725
transform 1 0 49404 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1676037725
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_91
timestamp 1676037725
transform 1 0 9476 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_103
timestamp 1676037725
transform 1 0 10580 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_115
timestamp 1676037725
transform 1 0 11684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_127
timestamp 1676037725
transform 1 0 12788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1676037725
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1676037725
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1676037725
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1676037725
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_437
timestamp 1676037725
transform 1 0 41308 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_461
timestamp 1676037725
transform 1 0 43516 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_473
timestamp 1676037725
transform 1 0 44620 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1676037725
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1676037725
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1676037725
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1676037725
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_77
timestamp 1676037725
transform 1 0 8188 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_82
timestamp 1676037725
transform 1 0 8648 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_94
timestamp 1676037725
transform 1 0 9752 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_106
timestamp 1676037725
transform 1 0 10856 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1676037725
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_521
timestamp 1676037725
transform 1 0 49036 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_525
timestamp 1676037725
transform 1 0 49404 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_22
timestamp 1676037725
transform 1 0 3128 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_33
timestamp 1676037725
transform 1 0 4140 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_50
timestamp 1676037725
transform 1 0 5704 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_78
timestamp 1676037725
transform 1 0 8280 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_89
timestamp 1676037725
transform 1 0 9292 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_106
timestamp 1676037725
transform 1 0 10856 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_134
timestamp 1676037725
transform 1 0 13432 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_145
timestamp 1676037725
transform 1 0 14444 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_162
timestamp 1676037725
transform 1 0 16008 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_190
timestamp 1676037725
transform 1 0 18584 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_236
timestamp 1676037725
transform 1 0 22816 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_244
timestamp 1676037725
transform 1 0 23552 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1676037725
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1676037725
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1676037725
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1676037725
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_511
timestamp 1676037725
transform 1 0 48116 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_11
timestamp 1676037725
transform 1 0 2116 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_29
timestamp 1676037725
transform 1 0 3772 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_37
timestamp 1676037725
transform 1 0 4508 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_61
timestamp 1676037725
transform 1 0 6716 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_65
timestamp 1676037725
transform 1 0 7084 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_85
timestamp 1676037725
transform 1 0 8924 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_141
timestamp 1676037725
transform 1 0 14076 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_166
timestamp 1676037725
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_197
timestamp 1676037725
transform 1 0 19228 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_201
timestamp 1676037725
transform 1 0 19596 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_218
timestamp 1676037725
transform 1 0 21160 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_230
timestamp 1676037725
transform 1 0 22264 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_238
timestamp 1676037725
transform 1 0 23000 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_243
timestamp 1676037725
transform 1 0 23460 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_251
timestamp 1676037725
transform 1 0 24196 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_263
timestamp 1676037725
transform 1 0 25300 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_275
timestamp 1676037725
transform 1 0 26404 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1676037725
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1676037725
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_511
timestamp 1676037725
transform 1 0 48116 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_525
timestamp 1676037725
transform 1 0 49404 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1676037725
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_45
timestamp 1676037725
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1676037725
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1676037725
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_101
timestamp 1676037725
transform 1 0 10396 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_118
timestamp 1676037725
transform 1 0 11960 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_138
timestamp 1676037725
transform 1 0 13800 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_157
timestamp 1676037725
transform 1 0 15548 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_174
timestamp 1676037725
transform 1 0 17112 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1676037725
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_215
timestamp 1676037725
transform 1 0 20884 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_232
timestamp 1676037725
transform 1 0 22448 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_239
timestamp 1676037725
transform 1 0 23092 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_243
timestamp 1676037725
transform 1 0 23460 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_247
timestamp 1676037725
transform 1 0 23828 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1676037725
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1676037725
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1676037725
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_289
timestamp 1676037725
transform 1 0 27692 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_297
timestamp 1676037725
transform 1 0 28428 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_303
timestamp 1676037725
transform 1 0 28980 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_321
timestamp 1676037725
transform 1 0 30636 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_327
timestamp 1676037725
transform 1 0 31188 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_331
timestamp 1676037725
transform 1 0 31556 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_343
timestamp 1676037725
transform 1 0 32660 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_355
timestamp 1676037725
transform 1 0 33764 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_359
timestamp 1676037725
transform 1 0 34132 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1676037725
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_377
timestamp 1676037725
transform 1 0 35788 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_383
timestamp 1676037725
transform 1 0 36340 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_387
timestamp 1676037725
transform 1 0 36708 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_399
timestamp 1676037725
transform 1 0 37812 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_411
timestamp 1676037725
transform 1 0 38916 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_415
timestamp 1676037725
transform 1 0 39284 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1676037725
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1676037725
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1676037725
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_457
timestamp 1676037725
transform 1 0 43148 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_465
timestamp 1676037725
transform 1 0 43884 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_472
timestamp 1676037725
transform 1 0 44528 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_495
timestamp 1676037725
transform 1 0 46644 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_500
timestamp 1676037725
transform 1 0 47104 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_508
timestamp 1676037725
transform 1 0 47840 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_521
timestamp 1676037725
transform 1 0 49036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_121
timestamp 1676037725
transform 1 0 12236 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_177
timestamp 1676037725
transform 1 0 17388 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_194
timestamp 1676037725
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_222
timestamp 1676037725
transform 1 0 21528 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_236
timestamp 1676037725
transform 1 0 22816 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_243
timestamp 1676037725
transform 1 0 23460 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_257
timestamp 1676037725
transform 1 0 24748 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_268
timestamp 1676037725
transform 1 0 25760 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_275
timestamp 1676037725
transform 1 0 26404 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1676037725
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_286
timestamp 1676037725
transform 1 0 27416 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_293
timestamp 1676037725
transform 1 0 28060 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_300
timestamp 1676037725
transform 1 0 28704 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_309
timestamp 1676037725
transform 1 0 29532 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_314
timestamp 1676037725
transform 1 0 29992 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_321
timestamp 1676037725
transform 1 0 30636 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_328
timestamp 1676037725
transform 1 0 31280 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_342
timestamp 1676037725
transform 1 0 32568 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_356
timestamp 1676037725
transform 1 0 33856 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_365
timestamp 1676037725
transform 1 0 34684 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_369
timestamp 1676037725
transform 1 0 35052 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_380
timestamp 1676037725
transform 1 0 36064 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_387
timestamp 1676037725
transform 1 0 36708 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1676037725
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_398
timestamp 1676037725
transform 1 0 37720 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_405
timestamp 1676037725
transform 1 0 38364 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_412
timestamp 1676037725
transform 1 0 39008 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_421
timestamp 1676037725
transform 1 0 39836 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_426
timestamp 1676037725
transform 1 0 40296 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_433
timestamp 1676037725
transform 1 0 40940 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_445
timestamp 1676037725
transform 1 0 42044 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_471
timestamp 1676037725
transform 1 0 44436 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_475
timestamp 1676037725
transform 1 0 44804 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_477
timestamp 1676037725
transform 1 0 44988 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_483
timestamp 1676037725
transform 1 0 45540 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_493
timestamp 1676037725
transform 1 0 46460 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_501
timestamp 1676037725
transform 1 0 47196 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_511
timestamp 1676037725
transform 1 0 48116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_519
timestamp 1676037725
transform 1 0 48852 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 49128 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input7 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 1564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input28
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input32
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 49128 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1676037725
transform 1 0 49036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 49036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 49128 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform 1 0 49036 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform 1 0 49036 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 49036 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 49128 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 49036 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 49036 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 49036 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 1676037725
transform 1 0 49036 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 49128 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform 1 0 49036 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 49036 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform 1 0 49036 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 49128 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 49128 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform 1 0 49036 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 49128 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 49128 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 48484 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 49036 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform 1 0 49036 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 49128 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 49036 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform 1 0 49036 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform 1 0 49036 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 49128 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 49036 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 21988 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 28428 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 28704 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 29716 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1676037725
transform 1 0 30360 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 31004 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1676037725
transform 1 0 31280 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 32292 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1676037725
transform 1 0 32936 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1676037725
transform 1 0 33580 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1676037725
transform 1 0 33856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1676037725
transform 1 0 22816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1676037725
transform 1 0 34868 0 1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1676037725
transform 1 0 35144 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1676037725
transform 1 0 36432 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1676037725
transform 1 0 36432 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 37444 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 38088 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1676037725
transform 1 0 38732 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 39008 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 40020 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 40664 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1676037725
transform 1 0 22540 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1676037725
transform 1 0 23184 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 23828 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1676037725
transform 1 0 24840 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1676037725
transform 1 0 25484 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1676037725
transform 1 0 26128 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 27140 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1676037725
transform 1 0 27784 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1676037725
transform 1 0 35420 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1676037725
transform 1 0 38640 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input96
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1676037725
transform 1 0 45356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform 1 0 42596 0 -1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1676037725
transform 1 0 48484 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input100
timestamp 1676037725
transform 1 0 48484 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform 1 0 47932 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1676037725
transform 1 0 47748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input103
timestamp 1676037725
transform 1 0 45908 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1676037725
transform 1 0 46828 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1676037725
transform 1 0 46736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform 1 0 47748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 1676037725
transform 1 0 48484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1676037725
transform 1 0 48668 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1676037725
transform 1 0 44160 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input110
timestamp 1676037725
transform 1 0 45172 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1656 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 1564 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 1564 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 1564 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 1564 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 1564 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 1564 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 1564 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 1564 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 1564 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 1564 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 1564 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 1564 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 1564 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 1564 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 1564 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 1564 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 47932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 47932 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 47932 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 47932 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 47932 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 47932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 47932 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 47932 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 47932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 47932 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 47932 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 47932 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 47932 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 47932 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 2300 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 9384 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 10488 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 11960 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 12328 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 14536 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 2024 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 14904 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 15640 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 17112 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 17480 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 19688 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 20056 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 20976 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 4232 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 5336 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 22172 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 49864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 49864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 49864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 49864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 49864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 49864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 49864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 49864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 49864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 49864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 49864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 49864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 49864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 49864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 49864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 49864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 49864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 49864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 49864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 49864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 49864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 49864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 49864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 49864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 49864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 49864 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 49864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 49864 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 49864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 49864 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 49864 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 49864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 49864 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 49864 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 49864 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 49864 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 49864 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 49864 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 49864 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 49864 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 49864 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 49864 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 49864 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 49864 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 49864 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 49864 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 49864 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 49864 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 49864 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 49864 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 49864 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 49864 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 49864 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 49864 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 49864 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24380 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24656 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22448 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20240 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21804 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20608 0 1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18400 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19872 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21712 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24564 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24840 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24748 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23184 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27600 0 -1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 26128 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27048 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27416 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24564 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27416 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29900 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31096 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33304 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33672 0 -1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34500 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 35144 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34960 0 1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37444 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35144 0 1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31924 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31280 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29716 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29992 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27324 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 28244 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29624 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 27416 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28520 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29900 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29992 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29716 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28244 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 41400 0 1 51136
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29440 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30728 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32384 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32936 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29440 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31280 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34500 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35144 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37260 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 35052 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35144 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32476 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32384 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34960 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34960 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35328 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37168 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34132 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34500 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33028 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32568 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32568 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24656 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24104 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24380 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24288 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23644 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19964 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19044 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19504 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20608 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21344 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18216 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14812 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15456 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15824 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13524 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13064 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14444 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15640 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16100 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27508 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24196 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 22356 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__258
timestamp 1676037725
transform 1 0 25392 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26772 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23552 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18124 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27600 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__211
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20792 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15272 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26772 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__214
timestamp 1676037725
transform 1 0 18676 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13064 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25116 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23460 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__216
timestamp 1676037725
transform 1 0 22632 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19688 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20884 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20700 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__259
timestamp 1676037725
transform 1 0 21160 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 19412 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20516 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19504 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13064 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27600 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25024 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 22264 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23736 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__260
timestamp 1676037725
transform 1 0 22172 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18492 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17020 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27784 0 1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24932 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 23000 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__261
timestamp 1676037725
transform 1 0 21528 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13156 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29808 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28336 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24564 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 25760 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29900 0 1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28336 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__212
timestamp 1676037725
transform 1 0 18676 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20516 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18308 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__213
timestamp 1676037725
transform 1 0 28612 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28336 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26220 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__215
timestamp 1676037725
transform 1 0 25576 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25852 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30360 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36156 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 25760 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30912 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__217
timestamp 1676037725
transform 1 0 26680 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33304 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37996 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 27508 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32568 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 32016 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 31004 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40020 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 36248 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32752 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28244 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35512 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33028 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__224
timestamp 1676037725
transform 1 0 34040 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40848 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34684 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36064 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 38640 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 30912 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__227
timestamp 1676037725
transform 1 0 32292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36708 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 37444 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 38824 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41124 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34592 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 33304 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 33580 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__218
timestamp 1676037725
transform 1 0 33488 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 30912 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32752 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33948 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 38272 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32108 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 31004 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 26128 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36064 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30452 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__219
timestamp 1676037725
transform 1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33396 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38180 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 31004 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 25852 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32200 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37444 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28796 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24932 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__222
timestamp 1676037725
transform 1 0 27416 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27600 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32108 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29992 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__223
timestamp 1676037725
transform 1 0 28980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37996 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__225
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28428 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31924 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28704 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__226
timestamp 1676037725
transform 1 0 27600 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27232 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30452 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38272 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__228
timestamp 1676037725
transform 1 0 28796 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27692 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35144 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27968 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26220 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38456 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 29716 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 31004 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__234
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 31096 0 1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27324 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32568 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38364 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33764 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28060 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__244
timestamp 1676037725
transform 1 0 25208 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 25208 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 39192 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 32292 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33764 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__252
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33028 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 39652 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 31004 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37536 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34960 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__253
timestamp 1676037725
transform 1 0 34868 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35788 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38180 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36064 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28060 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 29348 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 25576 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38640 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__230
timestamp 1676037725
transform 1 0 35512 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36248 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27968 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 38640 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38272 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 32292 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32752 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27140 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37536 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37812 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 31924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33120 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26680 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 35236 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36156 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 29072 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28704 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__235
timestamp 1676037725
transform 1 0 23828 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24472 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25668 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__236
timestamp 1676037725
transform 1 0 23552 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__237
timestamp 1676037725
transform 1 0 25760 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27048 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__238
timestamp 1676037725
transform 1 0 24196 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22908 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__239
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17480 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21068 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18952 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__240
timestamp 1676037725
transform 1 0 17296 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20148 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 21528 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__242
timestamp 1676037725
transform 1 0 20884 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 26220 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__243
timestamp 1676037725
transform 1 0 22356 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15272 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__245
timestamp 1676037725
transform 1 0 13524 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11960 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__246
timestamp 1676037725
transform 1 0 15456 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12696 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__247
timestamp 1676037725
transform 1 0 14720 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11960 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12880 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12420 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__248
timestamp 1676037725
transform 1 0 12788 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10212 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__249
timestamp 1676037725
transform 1 0 16192 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11960 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__250
timestamp 1676037725
transform 1 0 15456 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12236 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23460 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__251
timestamp 1676037725
transform 1 0 19872 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13248 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 29440 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 34592 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 39744 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 44896 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 56200 49294 57000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 2320 51000 2440 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 56200 1638 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 39040 800 39160 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 39856 800 39976 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 42304 800 42424 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 43936 800 44056 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 44752 800 44872 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 46384 800 46504 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 47200 800 47320 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 48832 800 48952 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 49648 800 49768 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 51280 800 51400 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 30064 800 30184 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 31696 800 31816 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 34960 800 35080 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 27616 51000 27736 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 35776 51000 35896 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 36592 51000 36712 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 37408 51000 37528 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 38224 51000 38344 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 39040 51000 39160 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 39856 51000 39976 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 40672 51000 40792 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 41488 51000 41608 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 42304 51000 42424 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 43120 51000 43240 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 28432 51000 28552 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 43936 51000 44056 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 44752 51000 44872 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 45568 51000 45688 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 46384 51000 46504 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 47200 51000 47320 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 48016 51000 48136 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 48832 51000 48952 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 49648 51000 49768 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 50464 51000 50584 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 51280 51000 51400 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 29248 51000 29368 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 30064 51000 30184 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 30880 51000 31000 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 31696 51000 31816 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 32512 51000 32632 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 33328 51000 33448 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 34144 51000 34264 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 34960 51000 35080 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 3136 51000 3256 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 11296 51000 11416 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 12112 51000 12232 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 12928 51000 13048 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 13744 51000 13864 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 14560 51000 14680 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 15376 51000 15496 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 16192 51000 16312 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 17008 51000 17128 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 17824 51000 17944 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 18640 51000 18760 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 3952 51000 4072 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 19456 51000 19576 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 20272 51000 20392 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 21088 51000 21208 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 22720 51000 22840 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 23536 51000 23656 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 24352 51000 24472 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 25168 51000 25288 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 25984 51000 26104 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 26800 51000 26920 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 4768 51000 4888 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 5584 51000 5704 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 6400 51000 6520 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 7216 51000 7336 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 8032 51000 8152 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 8848 51000 8968 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 9664 51000 9784 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 10480 51000 10600 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 56200 21602 57000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 56200 28042 57000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 56200 28686 57000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 56200 29330 57000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 56200 29974 57000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 56200 30618 57000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 56200 31262 57000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 56200 31906 57000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 56200 32550 57000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 56200 33194 57000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 56200 33838 57000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 56200 22246 57000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 56200 34482 57000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 56200 35126 57000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 56200 35770 57000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 56200 36414 57000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 56200 37058 57000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 56200 37702 57000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 56200 38346 57000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 56200 38990 57000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 56200 39634 57000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 56200 40278 57000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 56200 22890 57000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 56200 23534 57000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 56200 24178 57000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 56200 24822 57000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 56200 25466 57000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 56200 26110 57000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 56200 26754 57000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 56200 27398 57000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 56200 2282 57000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 56200 8722 57000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 56200 10654 57000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 56200 11298 57000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 56200 11942 57000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 56200 12586 57000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 56200 13230 57000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 56200 13874 57000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 56200 14518 57000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 56200 2926 57000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 56200 15806 57000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 56200 16450 57000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 56200 17094 57000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 56200 17738 57000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 56200 18382 57000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 56200 19670 57000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 56200 20958 57000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 56200 3570 57000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 56200 4214 57000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 56200 5502 57000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 56200 6146 57000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 56200 6790 57000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 56200 7434 57000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 56200 8078 57000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 56200 42210 57000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 200 nsew signal input
flabel metal2 s 42798 56200 42854 57000 0 FreeSans 224 90 0 0 reset_top_in
port 201 nsew signal input
flabel metal3 s 50200 52096 51000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal3 s 50200 52912 51000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal3 s 50200 53728 51000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal3 s 50200 54544 51000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 56200 43498 57000 0 FreeSans 224 90 0 0 test_enable_top_in
port 206 nsew signal input
flabel metal2 s 45374 56200 45430 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 56200 46074 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 56200 46718 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 56200 47362 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 56200 48006 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 56200 48650 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 56200 44142 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 56200 44786 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal3 s 0 52096 800 52216 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal3 s 0 53728 800 53848 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 54400 25484 54400 0 VGND
rlabel metal1 25484 53856 25484 53856 0 VPWR
rlabel metal1 22172 19482 22172 19482 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 20976 18598 20976 18598 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 18906 19482 18906 19482 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 16974 13362 16974 13362 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal2 23874 39100 23874 39100 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal2 21482 29478 21482 29478 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 23414 37740 23414 37740 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 18722 34068 18722 34068 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 20838 31858 20838 31858 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 18860 28730 18860 28730 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 18262 31858 18262 31858 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 17894 33422 17894 33422 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal2 17434 29920 17434 29920 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal2 16422 28492 16422 28492 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 18860 36210 18860 36210 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 16054 31969 16054 31969 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 15916 30022 15916 30022 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 21298 33354 21298 33354 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 17434 32742 17434 32742 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 13110 35122 13110 35122 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 15134 33558 15134 33558 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 27098 21022 27098 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 21528 26758 21528 26758 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 16238 33490 16238 33490 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18124 34034 18124 34034 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18676 33966 18676 33966 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18400 32198 18400 32198 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19780 31858 19780 31858 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19412 33898 19412 33898 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 20562 28186 20562 28186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 22310 29274 22310 29274 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 19826 29342 19826 29342 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15594 35802 15594 35802 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18492 26350 18492 26350 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 19182 26486 19182 26486 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15824 35734 15824 35734 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18170 33490 18170 33490 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17848 33626 17848 33626 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17066 27540 17066 27540 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15824 35462 15824 35462 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 17434 32368 17434 32368 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 17618 27370 17618 27370 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 18768 27438 18768 27438 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 18630 26911 18630 26911 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 11362 34034 11362 34034 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15594 27438 15594 27438 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 17434 19346 17434 19346 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 11822 35156 11822 35156 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17710 36278 17710 36278 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15594 33091 15594 33091 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17986 28186 17986 28186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14720 30770 14720 30770 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 14858 30906 14858 30906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 16974 28288 16974 28288 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 15778 29954 15778 29954 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 15870 29036 15870 29036 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 14766 35904 14766 35904 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14398 34102 14398 34102 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13248 34374 13248 34374 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14628 34714 14628 34714 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16790 35122 16790 35122 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20654 33626 20654 33626 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 16054 30226 16054 30226 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13892 34714 13892 34714 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13708 35054 13708 35054 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 14766 33422 14766 33422 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 15594 33626 15594 33626 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 13294 34646 13294 34646 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 22678 8058 22678 8058 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 21482 4590 21482 4590 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 25944 11050 25944 11050 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 26979 12410 26979 12410 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 25438 9112 25438 9112 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 21528 4522 21528 4522 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 24702 6289 24702 6289 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel via1 25507 12410 25507 12410 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 27508 8262 27508 8262 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 19412 11662 19412 11662 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 21022 11526 21022 11526 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel via1 24725 12410 24725 12410 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 24183 12818 24183 12818 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 19228 13158 19228 13158 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel via1 23575 12954 23575 12954 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 2254 1588 2254 1588 0 ccff_head
rlabel metal1 49312 51986 49312 51986 0 ccff_head_1
rlabel metal3 49734 2380 49734 2380 0 ccff_tail
rlabel metal1 1886 52530 1886 52530 0 ccff_tail_0
rlabel metal3 820 3196 820 3196 0 chanx_left_in[0]
rlabel metal3 820 11356 820 11356 0 chanx_left_in[10]
rlabel metal3 820 12172 820 12172 0 chanx_left_in[11]
rlabel metal3 820 12988 820 12988 0 chanx_left_in[12]
rlabel metal3 820 13804 820 13804 0 chanx_left_in[13]
rlabel metal3 820 14620 820 14620 0 chanx_left_in[14]
rlabel metal3 820 15436 820 15436 0 chanx_left_in[15]
rlabel metal3 820 16252 820 16252 0 chanx_left_in[16]
rlabel metal3 820 17068 820 17068 0 chanx_left_in[17]
rlabel metal3 1142 17884 1142 17884 0 chanx_left_in[18]
rlabel metal3 820 18700 820 18700 0 chanx_left_in[19]
rlabel metal3 820 4012 820 4012 0 chanx_left_in[1]
rlabel metal3 820 19516 820 19516 0 chanx_left_in[20]
rlabel metal3 820 20332 820 20332 0 chanx_left_in[21]
rlabel metal3 820 21148 820 21148 0 chanx_left_in[22]
rlabel metal3 820 21964 820 21964 0 chanx_left_in[23]
rlabel metal3 820 22780 820 22780 0 chanx_left_in[24]
rlabel metal3 820 23596 820 23596 0 chanx_left_in[25]
rlabel metal3 820 24412 820 24412 0 chanx_left_in[26]
rlabel metal3 820 25228 820 25228 0 chanx_left_in[27]
rlabel metal3 1188 26044 1188 26044 0 chanx_left_in[28]
rlabel metal3 820 26860 820 26860 0 chanx_left_in[29]
rlabel metal3 820 4828 820 4828 0 chanx_left_in[2]
rlabel metal3 820 5644 820 5644 0 chanx_left_in[3]
rlabel metal3 820 6460 820 6460 0 chanx_left_in[4]
rlabel metal3 820 7276 820 7276 0 chanx_left_in[5]
rlabel metal3 1142 8092 1142 8092 0 chanx_left_in[6]
rlabel metal3 820 8908 820 8908 0 chanx_left_in[7]
rlabel metal3 820 9724 820 9724 0 chanx_left_in[8]
rlabel metal3 820 10540 820 10540 0 chanx_left_in[9]
rlabel metal3 1004 27676 1004 27676 0 chanx_left_out[0]
rlabel metal2 2806 35955 2806 35955 0 chanx_left_out[10]
rlabel metal3 1004 36652 1004 36652 0 chanx_left_out[11]
rlabel metal3 1004 37468 1004 37468 0 chanx_left_out[12]
rlabel metal3 1004 38284 1004 38284 0 chanx_left_out[13]
rlabel metal3 1004 39100 1004 39100 0 chanx_left_out[14]
rlabel metal3 1372 39916 1372 39916 0 chanx_left_out[15]
rlabel metal3 1004 40732 1004 40732 0 chanx_left_out[16]
rlabel metal3 1004 41548 1004 41548 0 chanx_left_out[17]
rlabel metal3 1004 42364 1004 42364 0 chanx_left_out[18]
rlabel metal3 1004 43180 1004 43180 0 chanx_left_out[19]
rlabel metal3 1004 28492 1004 28492 0 chanx_left_out[1]
rlabel metal3 1372 43996 1372 43996 0 chanx_left_out[20]
rlabel metal3 1004 44812 1004 44812 0 chanx_left_out[21]
rlabel metal3 1004 45628 1004 45628 0 chanx_left_out[22]
rlabel metal3 1004 46444 1004 46444 0 chanx_left_out[23]
rlabel metal3 1004 47260 1004 47260 0 chanx_left_out[24]
rlabel metal3 1004 48076 1004 48076 0 chanx_left_out[25]
rlabel metal3 1004 48892 1004 48892 0 chanx_left_out[26]
rlabel metal3 1004 49708 1004 49708 0 chanx_left_out[27]
rlabel metal3 1004 50524 1004 50524 0 chanx_left_out[28]
rlabel metal3 1004 51340 1004 51340 0 chanx_left_out[29]
rlabel metal3 1004 29308 1004 29308 0 chanx_left_out[2]
rlabel metal3 1004 30124 1004 30124 0 chanx_left_out[3]
rlabel metal3 1004 30940 1004 30940 0 chanx_left_out[4]
rlabel metal3 1004 31756 1004 31756 0 chanx_left_out[5]
rlabel metal3 1004 32572 1004 32572 0 chanx_left_out[6]
rlabel metal3 1004 33388 1004 33388 0 chanx_left_out[7]
rlabel metal3 1372 34204 1372 34204 0 chanx_left_out[8]
rlabel metal3 1004 35020 1004 35020 0 chanx_left_out[9]
rlabel metal2 49358 27863 49358 27863 0 chanx_right_in_0[0]
rlabel metal1 48714 36142 48714 36142 0 chanx_right_in_0[10]
rlabel metal2 49082 36703 49082 36703 0 chanx_right_in_0[11]
rlabel metal2 49358 37655 49358 37655 0 chanx_right_in_0[12]
rlabel via2 49174 38267 49174 38267 0 chanx_right_in_0[13]
rlabel metal2 49174 39219 49174 39219 0 chanx_right_in_0[14]
rlabel metal2 49082 39967 49082 39967 0 chanx_right_in_0[15]
rlabel metal2 49358 40919 49358 40919 0 chanx_right_in_0[16]
rlabel via2 49082 41565 49082 41565 0 chanx_right_in_0[17]
rlabel metal2 49082 42517 49082 42517 0 chanx_right_in_0[18]
rlabel metal2 49174 43231 49174 43231 0 chanx_right_in_0[19]
rlabel via2 49082 28509 49082 28509 0 chanx_right_in_0[1]
rlabel metal2 49358 44183 49358 44183 0 chanx_right_in_0[20]
rlabel via2 49082 44829 49082 44829 0 chanx_right_in_0[21]
rlabel metal2 49082 45781 49082 45781 0 chanx_right_in_0[22]
rlabel metal2 49082 46495 49082 46495 0 chanx_right_in_0[23]
rlabel metal2 49358 47447 49358 47447 0 chanx_right_in_0[24]
rlabel via2 49358 48093 49358 48093 0 chanx_right_in_0[25]
rlabel metal2 49082 49045 49082 49045 0 chanx_right_in_0[26]
rlabel metal2 49358 49759 49358 49759 0 chanx_right_in_0[27]
rlabel metal2 49358 50711 49358 50711 0 chanx_right_in_0[28]
rlabel via2 48530 51357 48530 51357 0 chanx_right_in_0[29]
rlabel metal2 49174 29427 49174 29427 0 chanx_right_in_0[2]
rlabel metal2 49082 30175 49082 30175 0 chanx_right_in_0[3]
rlabel metal2 49358 31127 49358 31127 0 chanx_right_in_0[4]
rlabel via2 49082 31773 49082 31773 0 chanx_right_in_0[5]
rlabel metal2 49082 32725 49082 32725 0 chanx_right_in_0[6]
rlabel metal2 49174 33439 49174 33439 0 chanx_right_in_0[7]
rlabel metal2 49358 34391 49358 34391 0 chanx_right_in_0[8]
rlabel via2 49082 35037 49082 35037 0 chanx_right_in_0[9]
rlabel metal3 49734 3196 49734 3196 0 chanx_right_out_0[0]
rlabel metal2 49174 11509 49174 11509 0 chanx_right_out_0[10]
rlabel metal3 49734 12172 49734 12172 0 chanx_right_out_0[11]
rlabel metal3 49734 12988 49734 12988 0 chanx_right_out_0[12]
rlabel via2 49174 13821 49174 13821 0 chanx_right_out_0[13]
rlabel metal2 49174 14773 49174 14773 0 chanx_right_out_0[14]
rlabel metal3 49734 15436 49734 15436 0 chanx_right_out_0[15]
rlabel metal2 49174 16371 49174 16371 0 chanx_right_out_0[16]
rlabel via2 49174 17085 49174 17085 0 chanx_right_out_0[17]
rlabel metal2 49174 18037 49174 18037 0 chanx_right_out_0[18]
rlabel metal3 49734 18700 49734 18700 0 chanx_right_out_0[19]
rlabel via2 49174 4029 49174 4029 0 chanx_right_out_0[1]
rlabel metal3 49734 19516 49734 19516 0 chanx_right_out_0[20]
rlabel via2 49174 20349 49174 20349 0 chanx_right_out_0[21]
rlabel metal2 49174 21301 49174 21301 0 chanx_right_out_0[22]
rlabel metal3 49734 21964 49734 21964 0 chanx_right_out_0[23]
rlabel metal3 49734 22780 49734 22780 0 chanx_right_out_0[24]
rlabel via2 49174 23613 49174 23613 0 chanx_right_out_0[25]
rlabel metal2 49174 24565 49174 24565 0 chanx_right_out_0[26]
rlabel metal3 49734 25228 49734 25228 0 chanx_right_out_0[27]
rlabel metal2 48392 26044 48392 26044 0 chanx_right_out_0[28]
rlabel via2 49174 26877 49174 26877 0 chanx_right_out_0[29]
rlabel metal2 49174 4981 49174 4981 0 chanx_right_out_0[2]
rlabel metal3 49734 5644 49734 5644 0 chanx_right_out_0[3]
rlabel metal3 49734 6460 49734 6460 0 chanx_right_out_0[4]
rlabel via2 49174 7293 49174 7293 0 chanx_right_out_0[5]
rlabel metal2 49174 8245 49174 8245 0 chanx_right_out_0[6]
rlabel metal3 49734 8908 49734 8908 0 chanx_right_out_0[7]
rlabel metal3 49734 9724 49734 9724 0 chanx_right_out_0[8]
rlabel via2 49174 10557 49174 10557 0 chanx_right_out_0[9]
rlabel metal1 21896 53074 21896 53074 0 chany_top_in[0]
rlabel metal2 28244 56236 28244 56236 0 chany_top_in[10]
rlabel metal1 28796 53550 28796 53550 0 chany_top_in[11]
rlabel metal1 29624 54162 29624 54162 0 chany_top_in[12]
rlabel metal2 30176 56236 30176 56236 0 chany_top_in[13]
rlabel metal2 30590 55711 30590 55711 0 chany_top_in[14]
rlabel metal1 31372 53550 31372 53550 0 chany_top_in[15]
rlabel metal1 32200 54162 32200 54162 0 chany_top_in[16]
rlabel metal2 32522 55711 32522 55711 0 chany_top_in[17]
rlabel metal2 33166 55711 33166 55711 0 chany_top_in[18]
rlabel metal1 33948 53550 33948 53550 0 chany_top_in[19]
rlabel metal1 22632 53550 22632 53550 0 chany_top_in[1]
rlabel metal1 34684 53618 34684 53618 0 chany_top_in[20]
rlabel metal1 35144 54162 35144 54162 0 chany_top_in[21]
rlabel metal1 36294 54162 36294 54162 0 chany_top_in[22]
rlabel metal1 36524 53550 36524 53550 0 chany_top_in[23]
rlabel metal1 37352 54162 37352 54162 0 chany_top_in[24]
rlabel metal2 37674 55711 37674 55711 0 chany_top_in[25]
rlabel metal2 38318 55711 38318 55711 0 chany_top_in[26]
rlabel metal1 39100 53550 39100 53550 0 chany_top_in[27]
rlabel metal1 39928 54162 39928 54162 0 chany_top_in[28]
rlabel metal2 40250 55711 40250 55711 0 chany_top_in[29]
rlabel metal1 22816 54162 22816 54162 0 chany_top_in[2]
rlabel metal1 23460 54162 23460 54162 0 chany_top_in[3]
rlabel metal1 24104 54162 24104 54162 0 chany_top_in[4]
rlabel metal1 24932 54162 24932 54162 0 chany_top_in[5]
rlabel metal1 25576 54162 25576 54162 0 chany_top_in[6]
rlabel metal2 26082 55209 26082 55209 0 chany_top_in[7]
rlabel metal1 27048 54162 27048 54162 0 chany_top_in[8]
rlabel metal2 27370 55711 27370 55711 0 chany_top_in[9]
rlabel metal1 2530 53142 2530 53142 0 chany_top_out[0]
rlabel metal1 8556 54230 8556 54230 0 chany_top_out[10]
rlabel metal1 9614 52530 9614 52530 0 chany_top_out[11]
rlabel metal1 10120 53006 10120 53006 0 chany_top_out[12]
rlabel metal1 10672 54230 10672 54230 0 chany_top_out[13]
rlabel metal2 11270 54920 11270 54920 0 chany_top_out[14]
rlabel metal1 12190 52530 12190 52530 0 chany_top_out[15]
rlabel metal1 12834 53006 12834 53006 0 chany_top_out[16]
rlabel metal2 13202 55711 13202 55711 0 chany_top_out[17]
rlabel metal1 13708 54230 13708 54230 0 chany_top_out[18]
rlabel metal1 14766 52530 14766 52530 0 chany_top_out[19]
rlabel metal2 2898 54920 2898 54920 0 chany_top_out[1]
rlabel metal1 15272 53006 15272 53006 0 chany_top_out[20]
rlabel metal1 15824 54230 15824 54230 0 chany_top_out[21]
rlabel metal2 16422 54920 16422 54920 0 chany_top_out[22]
rlabel metal1 17342 52530 17342 52530 0 chany_top_out[23]
rlabel metal1 17986 53006 17986 53006 0 chany_top_out[24]
rlabel metal2 18354 54920 18354 54920 0 chany_top_out[25]
rlabel metal1 18860 54230 18860 54230 0 chany_top_out[26]
rlabel metal1 19918 53006 19918 53006 0 chany_top_out[27]
rlabel metal1 20424 54094 20424 54094 0 chany_top_out[28]
rlabel metal1 21436 53482 21436 53482 0 chany_top_out[29]
rlabel metal1 3404 54230 3404 54230 0 chany_top_out[2]
rlabel metal1 4508 52530 4508 52530 0 chany_top_out[3]
rlabel metal1 4968 53006 4968 53006 0 chany_top_out[4]
rlabel metal2 5474 55158 5474 55158 0 chany_top_out[5]
rlabel metal2 6118 54920 6118 54920 0 chany_top_out[6]
rlabel metal2 6762 54376 6762 54376 0 chany_top_out[7]
rlabel metal1 7682 53006 7682 53006 0 chany_top_out[8]
rlabel metal2 8050 55711 8050 55711 0 chany_top_out[9]
rlabel metal1 19366 38250 19366 38250 0 clknet_0_prog_clk
rlabel metal1 12696 5746 12696 5746 0 clknet_4_0_0_prog_clk
rlabel metal1 27508 42126 27508 42126 0 clknet_4_10_0_prog_clk
rlabel metal1 27646 40086 27646 40086 0 clknet_4_11_0_prog_clk
rlabel metal2 32706 15273 32706 15273 0 clknet_4_12_0_prog_clk
rlabel metal1 32844 33422 32844 33422 0 clknet_4_13_0_prog_clk
rlabel metal1 33028 40562 33028 40562 0 clknet_4_14_0_prog_clk
rlabel metal1 39376 51374 39376 51374 0 clknet_4_15_0_prog_clk
rlabel metal1 21160 9554 21160 9554 0 clknet_4_1_0_prog_clk
rlabel metal1 14214 35122 14214 35122 0 clknet_4_2_0_prog_clk
rlabel metal2 21390 32368 21390 32368 0 clknet_4_3_0_prog_clk
rlabel metal2 14490 38930 14490 38930 0 clknet_4_4_0_prog_clk
rlabel metal1 19688 38930 19688 38930 0 clknet_4_5_0_prog_clk
rlabel metal1 20608 40562 20608 40562 0 clknet_4_6_0_prog_clk
rlabel metal2 23322 42976 23322 42976 0 clknet_4_7_0_prog_clk
rlabel metal2 27094 13329 27094 13329 0 clknet_4_8_0_prog_clk
rlabel metal1 29440 38318 29440 38318 0 clknet_4_9_0_prog_clk
rlabel metal2 5566 1622 5566 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 8878 1622 8878 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 12190 1622 12190 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 15502 1622 15502 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 32062 1588 32062 1588 0 gfpga_pad_io_soc_in[0]
rlabel metal2 35374 1588 35374 1588 0 gfpga_pad_io_soc_in[1]
rlabel metal2 38686 1588 38686 1588 0 gfpga_pad_io_soc_in[2]
rlabel metal2 41998 1588 41998 1588 0 gfpga_pad_io_soc_in[3]
rlabel metal2 18814 1622 18814 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 22126 1622 22126 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 25438 1622 25438 1622 0 gfpga_pad_io_soc_out[2]
rlabel metal2 28750 1860 28750 1860 0 gfpga_pad_io_soc_out[3]
rlabel metal2 45310 1554 45310 1554 0 isol_n
rlabel metal2 9706 3944 9706 3944 0 net1
rlabel metal1 10120 16626 10120 16626 0 net10
rlabel metal1 47978 53040 47978 53040 0 net100
rlabel metal1 43470 53686 43470 53686 0 net101
rlabel metal1 47104 52870 47104 52870 0 net102
rlabel metal2 45862 54434 45862 54434 0 net103
rlabel metal1 38870 53958 38870 53958 0 net104
rlabel metal1 41469 53482 41469 53482 0 net105
rlabel metal1 38893 54298 38893 54298 0 net106
rlabel metal2 48714 50796 48714 50796 0 net107
rlabel metal2 48898 50558 48898 50558 0 net108
rlabel metal1 41400 53618 41400 53618 0 net109
rlabel metal2 2070 17119 2070 17119 0 net11
rlabel metal1 23414 52428 23414 52428 0 net110
rlabel metal1 39997 2618 39997 2618 0 net111
rlabel metal2 1702 46036 1702 46036 0 net112
rlabel metal2 11178 29376 11178 29376 0 net113
rlabel metal1 1794 36176 1794 36176 0 net114
rlabel metal2 1794 36550 1794 36550 0 net115
rlabel metal2 1794 38148 1794 38148 0 net116
rlabel metal1 15318 39814 15318 39814 0 net117
rlabel metal1 1794 39440 1794 39440 0 net118
rlabel metal1 1794 40052 1794 40052 0 net119
rlabel metal1 14260 18054 14260 18054 0 net12
rlabel metal2 12282 40902 12282 40902 0 net120
rlabel metal1 12190 41242 12190 41242 0 net121
rlabel metal1 8556 42670 8556 42670 0 net122
rlabel metal1 1794 43316 1794 43316 0 net123
rlabel metal2 11086 29546 11086 29546 0 net124
rlabel metal1 1794 44302 1794 44302 0 net125
rlabel metal2 11086 44404 11086 44404 0 net126
rlabel metal2 12282 44914 12282 44914 0 net127
rlabel metal2 8694 44982 8694 44982 0 net128
rlabel metal2 4094 45526 4094 45526 0 net129
rlabel metal1 4347 18598 4347 18598 0 net13
rlabel metal2 11086 47124 11086 47124 0 net130
rlabel metal2 5842 46580 5842 46580 0 net131
rlabel metal2 5750 46852 5750 46852 0 net132
rlabel metal2 5658 47974 5658 47974 0 net133
rlabel metal1 4692 51374 4692 51374 0 net134
rlabel metal2 8694 30362 8694 30362 0 net135
rlabel metal1 4600 30226 4600 30226 0 net136
rlabel metal1 4347 31314 4347 31314 0 net137
rlabel metal2 12742 32062 12742 32062 0 net138
rlabel metal2 16698 33830 16698 33830 0 net139
rlabel metal2 25346 5405 25346 5405 0 net14
rlabel metal2 8602 35564 8602 35564 0 net140
rlabel metal2 10994 34748 10994 34748 0 net141
rlabel metal1 2277 35054 2277 35054 0 net142
rlabel metal2 36478 6460 36478 6460 0 net143
rlabel metal2 38318 16797 38318 16797 0 net144
rlabel metal1 45816 19210 45816 19210 0 net145
rlabel metal1 40802 17578 40802 17578 0 net146
rlabel metal1 44114 18666 44114 18666 0 net147
rlabel metal1 41584 19210 41584 19210 0 net148
rlabel metal1 44482 21930 44482 21930 0 net149
rlabel metal1 9430 19686 9430 19686 0 net15
rlabel metal1 44068 20842 44068 20842 0 net150
rlabel metal2 42826 19278 42826 19278 0 net151
rlabel metal2 47058 20910 47058 20910 0 net152
rlabel metal2 45126 21420 45126 21420 0 net153
rlabel metal1 37812 10506 37812 10506 0 net154
rlabel metal2 46966 22202 46966 22202 0 net155
rlabel metal2 44206 22542 44206 22542 0 net156
rlabel metal2 44298 23630 44298 23630 0 net157
rlabel metal2 44758 24412 44758 24412 0 net158
rlabel metal2 45310 25466 45310 25466 0 net159
rlabel metal1 9384 20230 9384 20230 0 net16
rlabel metal1 47426 23698 47426 23698 0 net160
rlabel metal1 47886 24786 47886 24786 0 net161
rlabel metal1 46966 25262 46966 25262 0 net162
rlabel metal2 46506 28492 46506 28492 0 net163
rlabel metal2 46782 29070 46782 29070 0 net164
rlabel metal1 37536 11050 37536 11050 0 net165
rlabel metal2 43838 10234 43838 10234 0 net166
rlabel metal2 38410 9690 38410 9690 0 net167
rlabel metal2 38594 10302 38594 10302 0 net168
rlabel metal2 37766 11152 37766 11152 0 net169
rlabel metal1 10948 21318 10948 21318 0 net17
rlabel metal1 45310 16626 45310 16626 0 net170
rlabel metal2 38502 12988 38502 12988 0 net171
rlabel metal1 38364 16626 38364 16626 0 net172
rlabel metal1 2530 53006 2530 53006 0 net173
rlabel metal1 7406 54128 7406 54128 0 net174
rlabel metal1 9706 52462 9706 52462 0 net175
rlabel metal1 11178 53074 11178 53074 0 net176
rlabel metal1 10258 54162 10258 54162 0 net177
rlabel metal1 10718 53516 10718 53516 0 net178
rlabel metal1 13018 52462 13018 52462 0 net179
rlabel metal1 10580 21862 10580 21862 0 net18
rlabel metal1 12834 53108 12834 53108 0 net180
rlabel metal1 13892 53550 13892 53550 0 net181
rlabel metal1 13156 54162 13156 54162 0 net182
rlabel metal1 15824 52462 15824 52462 0 net183
rlabel metal2 2070 49028 2070 49028 0 net184
rlabel metal1 15180 53074 15180 53074 0 net185
rlabel metal1 15134 49810 15134 49810 0 net186
rlabel metal1 15870 53618 15870 53618 0 net187
rlabel metal1 18400 52462 18400 52462 0 net188
rlabel metal1 18630 53074 18630 53074 0 net189
rlabel metal1 3358 23154 3358 23154 0 net19
rlabel metal1 17710 53482 17710 53482 0 net190
rlabel metal1 18906 54162 18906 54162 0 net191
rlabel metal1 21252 52666 21252 52666 0 net192
rlabel metal1 21114 54162 21114 54162 0 net193
rlabel metal1 21206 53584 21206 53584 0 net194
rlabel metal1 3036 54162 3036 54162 0 net195
rlabel metal1 4600 52462 4600 52462 0 net196
rlabel metal1 5290 53074 5290 53074 0 net197
rlabel metal1 4876 54162 4876 54162 0 net198
rlabel metal1 5474 53516 5474 53516 0 net199
rlabel metal2 49174 51612 49174 51612 0 net2
rlabel metal1 3404 23766 3404 23766 0 net20
rlabel metal1 7682 52462 7682 52462 0 net200
rlabel metal1 8694 53074 8694 53074 0 net201
rlabel metal1 7958 53550 7958 53550 0 net202
rlabel metal1 6831 2414 6831 2414 0 net203
rlabel metal1 10212 2414 10212 2414 0 net204
rlabel metal1 13294 2414 13294 2414 0 net205
rlabel metal2 17894 3434 17894 3434 0 net206
rlabel metal2 19642 4522 19642 4522 0 net207
rlabel metal2 22218 4012 22218 4012 0 net208
rlabel metal2 25254 4012 25254 4012 0 net209
rlabel metal1 15088 36006 15088 36006 0 net21
rlabel metal2 28842 4318 28842 4318 0 net210
rlabel metal1 21206 41106 21206 41106 0 net211
rlabel metal2 20470 44846 20470 44846 0 net212
rlabel metal2 28750 44676 28750 44676 0 net213
rlabel metal1 18722 40154 18722 40154 0 net214
rlabel metal1 26036 39406 26036 39406 0 net215
rlabel metal1 21482 39406 21482 39406 0 net216
rlabel metal1 27784 39610 27784 39610 0 net217
rlabel metal2 33718 34680 33718 34680 0 net218
rlabel metal1 34914 34102 34914 34102 0 net219
rlabel metal1 2668 25330 2668 25330 0 net22
rlabel metal2 32246 38624 32246 38624 0 net220
rlabel metal1 29578 35054 29578 35054 0 net221
rlabel metal1 27830 32878 27830 32878 0 net222
rlabel metal1 29394 31450 29394 31450 0 net223
rlabel metal1 33856 37434 33856 37434 0 net224
rlabel metal1 29394 29614 29394 29614 0 net225
rlabel metal1 27738 31450 27738 31450 0 net226
rlabel metal1 32476 33490 32476 33490 0 net227
rlabel metal1 28566 41242 28566 41242 0 net228
rlabel metal2 29578 33694 29578 33694 0 net229
rlabel metal1 13156 36890 13156 36890 0 net23
rlabel metal1 35052 34170 35052 34170 0 net230
rlabel metal1 32614 31314 32614 31314 0 net231
rlabel metal1 33120 32946 33120 32946 0 net232
rlabel metal2 29118 29648 29118 29648 0 net233
rlabel metal1 34132 44914 34132 44914 0 net234
rlabel metal1 24518 32878 24518 32878 0 net235
rlabel metal1 24380 33966 24380 33966 0 net236
rlabel metal2 25990 34544 25990 34544 0 net237
rlabel metal2 24978 30906 24978 30906 0 net238
rlabel metal2 22218 36278 22218 36278 0 net239
rlabel metal1 14812 37298 14812 37298 0 net24
rlabel metal1 17526 37876 17526 37876 0 net240
rlabel metal1 21390 37434 21390 37434 0 net241
rlabel metal1 20608 37230 20608 37230 0 net242
rlabel metal2 22402 29444 22402 29444 0 net243
rlabel metal1 26956 40494 26956 40494 0 net244
rlabel metal1 14214 33966 14214 33966 0 net245
rlabel metal1 15778 39066 15778 39066 0 net246
rlabel metal1 14812 39610 14812 39610 0 net247
rlabel metal1 12972 37842 12972 37842 0 net248
rlabel metal1 15916 41582 15916 41582 0 net249
rlabel metal1 37904 10642 37904 10642 0 net25
rlabel metal2 15962 43588 15962 43588 0 net250
rlabel metal1 19320 47022 19320 47022 0 net251
rlabel metal2 34178 45764 34178 45764 0 net252
rlabel metal1 35236 43282 35236 43282 0 net253
rlabel metal1 23322 30362 23322 30362 0 net254
rlabel metal2 22218 30430 22218 30430 0 net255
rlabel metal1 14214 32878 14214 32878 0 net256
rlabel metal2 18998 33643 18998 33643 0 net257
rlabel metal1 25070 38794 25070 38794 0 net258
rlabel metal1 20332 40426 20332 40426 0 net259
rlabel metal2 17250 6221 17250 6221 0 net26
rlabel metal1 21298 44506 21298 44506 0 net260
rlabel metal2 18538 46478 18538 46478 0 net261
rlabel metal1 25024 42670 25024 42670 0 net262
rlabel metal1 9384 6630 9384 6630 0 net27
rlabel metal1 11040 7174 11040 7174 0 net28
rlabel metal1 14007 8330 14007 8330 0 net29
rlabel metal1 8280 3366 8280 3366 0 net3
rlabel metal1 15226 8806 15226 8806 0 net30
rlabel metal1 8234 9894 8234 9894 0 net31
rlabel metal1 38548 16082 38548 16082 0 net32
rlabel metal2 36570 30158 36570 30158 0 net33
rlabel metal2 49266 36584 49266 36584 0 net34
rlabel via2 48346 36635 48346 36635 0 net35
rlabel metal1 45540 37774 45540 37774 0 net36
rlabel metal2 49266 38046 49266 38046 0 net37
rlabel metal2 49266 39100 49266 39100 0 net38
rlabel metal2 15870 39032 15870 39032 0 net39
rlabel metal1 11914 11594 11914 11594 0 net4
rlabel metal2 49174 40698 49174 40698 0 net40
rlabel metal2 49266 40426 49266 40426 0 net41
rlabel metal2 47242 41480 47242 41480 0 net42
rlabel metal2 49266 43690 49266 43690 0 net43
rlabel metal1 45540 28424 45540 28424 0 net44
rlabel metal1 45540 44438 45540 44438 0 net45
rlabel metal2 47426 42840 47426 42840 0 net46
rlabel metal1 48944 45798 48944 45798 0 net47
rlabel metal1 20102 35054 20102 35054 0 net48
rlabel metal2 42826 46444 42826 46444 0 net49
rlabel metal1 32936 17170 32936 17170 0 net5
rlabel metal2 43378 46410 43378 46410 0 net50
rlabel metal1 45540 49096 45540 49096 0 net51
rlabel metal2 43470 48382 43470 48382 0 net52
rlabel metal2 42826 49232 42826 49232 0 net53
rlabel metal1 48806 51306 48806 51306 0 net54
rlabel metal1 45540 29648 45540 29648 0 net55
rlabel metal2 49266 29920 49266 29920 0 net56
rlabel metal1 49174 31212 49174 31212 0 net57
rlabel metal1 45540 31892 45540 31892 0 net58
rlabel metal1 19734 33014 19734 33014 0 net59
rlabel metal2 1886 22780 1886 22780 0 net6
rlabel metal1 16974 34680 16974 34680 0 net60
rlabel metal1 48300 34714 48300 34714 0 net61
rlabel metal2 48346 34969 48346 34969 0 net62
rlabel metal1 23690 52870 23690 52870 0 net63
rlabel metal2 27876 53516 27876 53516 0 net64
rlabel metal1 28704 53414 28704 53414 0 net65
rlabel metal1 29440 53958 29440 53958 0 net66
rlabel metal1 30498 50694 30498 50694 0 net67
rlabel metal1 30912 53958 30912 53958 0 net68
rlabel metal1 30912 53414 30912 53414 0 net69
rlabel metal1 1794 13804 1794 13804 0 net7
rlabel metal1 32660 50490 32660 50490 0 net70
rlabel metal1 32798 53958 32798 53958 0 net71
rlabel metal2 33626 51918 33626 51918 0 net72
rlabel metal1 32844 53414 32844 53414 0 net73
rlabel metal1 23138 53414 23138 53414 0 net74
rlabel metal1 32430 53482 32430 53482 0 net75
rlabel metal1 32614 54094 32614 54094 0 net76
rlabel metal1 31970 54230 31970 54230 0 net77
rlabel metal1 32982 53686 32982 53686 0 net78
rlabel metal2 37490 54298 37490 54298 0 net79
rlabel metal1 11776 14790 11776 14790 0 net8
rlabel metal1 35052 54026 35052 54026 0 net80
rlabel metal1 36938 54162 36938 54162 0 net81
rlabel metal1 37122 49946 37122 49946 0 net82
rlabel metal1 38134 54230 38134 54230 0 net83
rlabel metal2 40710 54264 40710 54264 0 net84
rlabel metal1 24012 53958 24012 53958 0 net85
rlabel metal1 23230 54264 23230 54264 0 net86
rlabel metal1 23874 54060 23874 54060 0 net87
rlabel metal1 27508 54298 27508 54298 0 net88
rlabel metal1 25806 53958 25806 53958 0 net89
rlabel metal1 35558 19346 35558 19346 0 net9
rlabel metal1 28336 54094 28336 54094 0 net90
rlabel metal1 27324 53958 27324 53958 0 net91
rlabel metal2 28428 53958 28428 53958 0 net92
rlabel metal2 24794 9146 24794 9146 0 net93
rlabel metal1 31004 2346 31004 2346 0 net94
rlabel metal1 38962 2516 38962 2516 0 net95
rlabel metal1 38870 2448 38870 2448 0 net96
rlabel metal1 24932 8466 24932 8466 0 net97
rlabel metal1 21482 5644 21482 5644 0 net98
rlabel metal1 42596 52530 42596 52530 0 net99
rlabel metal2 48622 2098 48622 2098 0 prog_clk
rlabel metal1 42412 54230 42412 54230 0 prog_reset_top_in
rlabel metal2 48530 52309 48530 52309 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel via2 48530 52989 48530 52989 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 48208 53550 48208 53550 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 47840 53142 47840 53142 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 29670 34714 29670 34714 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal2 24978 43826 24978 43826 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal2 24794 38794 24794 38794 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 27002 41718 27002 41718 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal1 21206 39474 21206 39474 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal2 20194 43486 20194 43486 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel metal1 20884 37774 20884 37774 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 21436 43418 21436 43418 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 21574 46342 21574 46342 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal1 21712 44710 21712 44710 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 20608 46478 20608 46478 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal2 21482 47974 21482 47974 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 23138 39474 23138 39474 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal1 19780 47702 19780 47702 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal1 25530 46478 25530 46478 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal2 25162 40437 25162 40437 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal2 26634 44676 26634 44676 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal2 21942 42330 21942 42330 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal2 26450 43843 26450 43843 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 20608 42602 20608 42602 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal1 21206 47124 21206 47124 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal1 29440 47090 29440 47090 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal1 23552 47566 23552 47566 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal1 27416 48042 27416 48042 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal1 28513 49606 28513 49606 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 26634 46954 26634 46954 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal1 19734 40086 19734 40086 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel metal1 27186 41582 27186 41582 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 18814 40494 18814 40494 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal1 32338 48008 32338 48008 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel metal1 26726 39474 26726 39474 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal1 21620 40154 21620 40154 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 20378 39508 20378 39508 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal1 21252 45322 21252 45322 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal1 33902 42806 33902 42806 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel metal2 34178 45186 34178 45186 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 29210 43384 29210 43384 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal2 39238 40664 39238 40664 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal2 34086 39712 34086 39712 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal1 34086 38182 34086 38182 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 33258 39950 33258 39950 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal1 32338 36278 32338 36278 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal1 32522 39610 32522 39610 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal1 32982 38250 32982 38250 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal1 34132 41174 34132 41174 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal1 32890 46512 32890 46512 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal2 32706 40131 32706 40131 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal1 30176 35530 30176 35530 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal1 27324 39338 27324 39338 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal1 29578 39610 29578 39610 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal1 32706 35190 32706 35190 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal1 27278 37774 27278 37774 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 28888 37978 28888 37978 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal1 34086 32402 34086 32402 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal1 29532 39950 29532 39950 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal1 30028 34374 30028 34374 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal1 36110 39066 36110 39066 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel via2 28934 31875 28934 31875 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal2 35466 38624 35466 38624 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal2 32154 32334 32154 32334 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal2 30866 37162 30866 37162 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 28421 34374 28421 34374 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 37030 39304 37030 39304 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal2 37766 39712 37766 39712 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal1 30866 48178 30866 48178 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel metal1 41216 51782 41216 51782 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 34270 47532 34270 47532 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal2 36846 43248 36846 43248 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal1 32430 37128 32430 37128 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal1 38318 40562 38318 40562 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 36340 41038 36340 41038 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 36800 36890 36800 36890 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel metal1 35328 36074 35328 36074 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 34684 36822 34684 36822 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 33580 38862 33580 38862 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal1 37122 37128 37122 37128 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 34730 34986 34730 34986 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal1 33120 34034 33120 34034 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 36432 35802 36432 35802 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 37352 34374 37352 34374 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal1 30728 34034 30728 34034 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal1 34960 33830 34960 33830 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 33580 32742 33580 32742 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal2 33534 49878 33534 49878 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal1 32292 48790 32292 48790 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 32062 47260 32062 47260 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 24702 35598 24702 35598 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel metal1 28106 33286 28106 33286 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 23322 36686 23322 36686 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal2 25898 36652 25898 36652 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 25530 36346 25530 36346 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 25668 36686 25668 36686 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal2 23966 34884 23966 34884 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 25898 34714 25898 34714 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal2 21390 35122 21390 35122 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 24702 32198 24702 32198 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 19451 34374 19451 34374 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal2 21482 33728 21482 33728 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 19596 35734 19596 35734 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal1 20286 34510 20286 34510 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 22402 36278 22402 36278 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal2 21298 35292 21298 35292 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20286 31212 20286 31212 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal1 23920 34714 23920 34714 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal2 31602 44302 31602 44302 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal1 33258 44336 33258 44336 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 34362 43690 34362 43690 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 15778 33864 15778 33864 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal1 15318 31722 15318 31722 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 17296 37298 17296 37298 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 18446 35632 18446 35632 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 15088 37638 15088 37638 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal2 16146 36992 16146 36992 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 14812 38250 14812 38250 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal1 14352 35598 14352 35598 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 16560 40426 16560 40426 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal2 16238 38896 16238 38896 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 17434 43656 17434 43656 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal1 17526 40698 17526 40698 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 20010 44676 20010 44676 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel metal1 35420 45866 35420 45866 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal1 39652 45390 39652 45390 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 34638 45390 34638 45390 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 40250 44268 40250 44268 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 38456 44914 38456 44914 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 14628 40970 14628 40970 0 sb_1__0_.mux_left_track_1.out
rlabel metal2 27278 46019 27278 46019 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27370 44846 27370 44846 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24150 39066 24150 39066 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22402 41208 22402 41208 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23782 44982 23782 44982 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23644 41242 23644 41242 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 18538 41174 18538 41174 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7544 43214 7544 43214 0 sb_1__0_.mux_left_track_11.out
rlabel metal2 21022 47294 21022 47294 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 45832 21482 45832 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20378 43622 20378 43622 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19688 40698 19688 40698 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 18630 44268 18630 44268 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19044 42670 19044 42670 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13294 41548 13294 41548 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18032 37162 18032 37162 0 sb_1__0_.mux_left_track_13.out
rlabel metal1 25760 48790 25760 48790 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 25070 47430 25070 47430 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21758 44370 21758 44370 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18952 43282 18952 43282 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19596 43418 19596 43418 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17894 41582 17894 41582 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 6854 44846 6854 44846 0 sb_1__0_.mux_left_track_21.out
rlabel metal2 22494 48926 22494 48926 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23920 47226 23920 47226 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18860 44710 18860 44710 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22034 47872 22034 47872 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18998 45050 18998 45050 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14996 45458 14996 45458 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 14996 38726 14996 38726 0 sb_1__0_.mux_left_track_29.out
rlabel metal2 26358 47736 26358 47736 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27324 45322 27324 45322 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24840 39610 24840 39610 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25898 45560 25898 45560 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24196 42534 24196 42534 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19734 39916 19734 39916 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 13524 36788 13524 36788 0 sb_1__0_.mux_left_track_3.out
rlabel metal1 26220 48314 26220 48314 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26082 41786 26082 41786 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21298 42636 21298 42636 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20332 41514 20332 41514 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20792 40970 20792 40970 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17388 32402 17388 32402 0 sb_1__0_.mux_left_track_37.out
rlabel metal2 27600 50388 27600 50388 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 28382 47430 28382 47430 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21160 47022 21160 47022 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22034 45730 22034 45730 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18860 40494 18860 40494 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 15272 37978 15272 37978 0 sb_1__0_.mux_left_track_45.out
rlabel metal1 30636 49130 30636 49130 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 29026 48382 29026 48382 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28014 44506 28014 44506 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16330 41990 16330 41990 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9476 40086 9476 40086 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 23966 43758 23966 43758 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25898 40698 25898 40698 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18400 38998 18400 38998 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17342 39610 17342 39610 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 16974 39814 16974 39814 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8004 31722 8004 31722 0 sb_1__0_.mux_left_track_53.out
rlabel metal1 32338 49708 32338 49708 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24058 40494 24058 40494 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25898 39984 25898 39984 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20148 36822 20148 36822 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13501 43622 13501 43622 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 24150 40018 24150 40018 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25070 38522 25070 38522 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19872 38522 19872 38522 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22770 39576 22770 39576 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20516 39338 20516 39338 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17618 38250 17618 38250 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 39008 35462 39008 35462 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 31096 44506 31096 44506 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33994 44336 33994 44336 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27968 36550 27968 36550 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33718 42738 33718 42738 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33718 41480 33718 41480 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 33672 40052 33672 40052 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 44666 28118 44666 28118 0 sb_1__0_.mux_right_track_10.out
rlabel metal1 34316 48518 34316 48518 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33258 44778 33258 44778 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34040 39066 34040 39066 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33994 37230 33994 37230 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38456 38386 38456 38386 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38686 38216 38686 38216 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39698 35972 39698 35972 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 44574 29070 44574 29070 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 36340 42126 36340 42126 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36386 42262 36386 42262 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30590 35598 30590 35598 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34454 34918 34454 34918 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33810 35258 33810 35258 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 35328 35258 35328 35258 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43976 30702 43976 30702 0 sb_1__0_.mux_right_track_2.out
rlabel metal1 32982 45526 32982 45526 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32660 45594 32660 45594 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28428 35190 28428 35190 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37260 42262 37260 42262 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 33442 42024 33442 42024 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39882 35054 39882 35054 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39422 27098 39422 27098 0 sb_1__0_.mux_right_track_20.out
rlabel metal1 30590 43758 30590 43758 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30590 43690 30590 43690 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27278 31926 27278 31926 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32706 36482 32706 36482 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32177 36074 32177 36074 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37214 36074 37214 36074 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 43930 25194 43930 25194 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 29302 41174 29302 41174 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29670 41242 29670 41242 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26726 32810 26726 32810 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32614 36567 32614 36567 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 31786 34476 31786 34476 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33810 35190 33810 35190 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 42228 19414 42228 19414 0 sb_1__0_.mux_right_track_36.out
rlabel metal1 31050 40562 31050 40562 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 31142 40494 31142 40494 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33534 32334 33534 32334 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33902 31756 33902 31756 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35696 32266 35696 32266 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 45862 31416 45862 31416 0 sb_1__0_.mux_right_track_4.out
rlabel metal1 36156 43418 36156 43418 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35742 43418 35742 43418 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 31970 35292 31970 35292 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37490 37842 37490 37842 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37168 37910 37168 37910 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 40480 33490 40480 33490 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43838 16558 43838 16558 0 sb_1__0_.mux_right_track_44.out
rlabel metal2 31418 36380 31418 36380 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32338 30600 32338 30600 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33672 31994 33672 31994 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40250 15062 40250 15062 0 sb_1__0_.mux_right_track_52.out
rlabel metal1 30774 32538 30774 32538 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29072 31178 29072 31178 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34500 23698 34500 23698 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 44206 32096 44206 32096 0 sb_1__0_.mux_right_track_6.out
rlabel metal1 37122 44778 37122 44778 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 37122 46002 37122 46002 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38318 38318 38318 38318 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33074 33558 33074 33558 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 39330 39474 39330 39474 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38364 38522 38364 38522 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 41354 37060 41354 37060 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 25024 53550 25024 53550 0 sb_1__0_.mux_top_track_0.out
rlabel metal2 34914 47396 34914 47396 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36938 47770 36938 47770 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24794 41321 24794 41321 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28060 43690 28060 43690 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35006 47770 35006 47770 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 28796 43962 28796 43962 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 29072 48586 29072 48586 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 25070 44506 25070 44506 0 sb_1__0_.mux_top_track_10.out
rlabel metal2 36570 41321 36570 41321 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37720 40698 37720 40698 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 31786 39168 31786 39168 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28520 34170 28520 34170 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 29762 39508 29762 39508 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 27232 44982 27232 44982 0 sb_1__0_.mux_top_track_12.out
rlabel metal2 39146 38658 39146 38658 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37720 37978 37720 37978 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32384 34374 32384 34374 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34017 38454 34017 38454 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26956 43418 26956 43418 0 sb_1__0_.mux_top_track_14.out
rlabel metal2 38778 38522 38778 38522 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36708 36550 36708 36550 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32982 32538 32982 32538 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 39270 28612 39270 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21620 49810 21620 49810 0 sb_1__0_.mux_top_track_16.out
rlabel metal1 37950 34714 37950 34714 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37858 34476 37858 34476 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33304 31994 33304 31994 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32706 37094 32706 37094 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23690 41446 23690 41446 0 sb_1__0_.mux_top_track_18.out
rlabel metal1 36064 32538 36064 32538 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35420 32198 35420 32198 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29486 33966 29486 33966 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 26956 34102 26956 34102 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 25668 53074 25668 53074 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 35144 48314 35144 48314 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37858 47226 37858 47226 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30084 44506 30084 44506 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34684 49402 34684 49402 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 31096 45322 31096 45322 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29348 50490 29348 50490 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17664 44506 17664 44506 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 25622 37910 25622 37910 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24748 33082 24748 33082 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 44200 20838 44200 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18216 45322 18216 45322 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 24150 37978 24150 37978 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 34170 24104 34170 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21252 41276 21252 41276 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19366 46138 19366 46138 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 25484 38318 25484 38318 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23506 35258 23506 35258 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19688 41400 19688 41400 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19228 42534 19228 42534 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 23368 37230 23368 37230 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23966 30906 23966 30906 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19964 39270 19964 39270 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17526 42568 17526 42568 0 sb_1__0_.mux_top_track_28.out
rlabel metal2 21206 33626 21206 33626 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17618 42670 17618 42670 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16146 46954 16146 46954 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 20286 31994 20286 31994 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17756 37638 17756 37638 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15226 44506 15226 44506 0 sb_1__0_.mux_top_track_32.out
rlabel metal1 20148 33014 20148 33014 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18262 37978 18262 37978 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15502 44234 15502 44234 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 21896 32538 21896 32538 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19780 37094 19780 37094 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16652 42534 16652 42534 0 sb_1__0_.mux_top_track_36.out
rlabel metal1 24380 36890 24380 36890 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21942 29274 21942 29274 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21988 36550 21988 36550 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23782 52530 23782 52530 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 33442 44506 33442 44506 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34914 44438 34914 44438 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 30866 44472 30866 44472 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 40698 28612 40698 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 28428 45050 28428 45050 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12006 45458 12006 45458 0 sb_1__0_.mux_top_track_40.out
rlabel metal1 15088 33830 15088 33830 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13248 41650 13248 41650 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11638 47974 11638 47974 0 sb_1__0_.mux_top_track_42.out
rlabel metal1 16974 35802 16974 35802 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15272 39066 15272 39066 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10994 45322 10994 45322 0 sb_1__0_.mux_top_track_44.out
rlabel metal1 15548 36346 15548 36346 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13570 40154 13570 40154 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9936 44506 9936 44506 0 sb_1__0_.mux_top_track_46.out
rlabel metal1 12880 32538 12880 32538 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 41446 12466 41446 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10120 51306 10120 51306 0 sb_1__0_.mux_top_track_48.out
rlabel metal1 17894 39066 17894 39066 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14398 41786 14398 41786 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9568 51986 9568 51986 0 sb_1__0_.mux_top_track_50.out
rlabel metal1 17986 39610 17986 39610 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15364 43418 15364 43418 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9936 52938 9936 52938 0 sb_1__0_.mux_top_track_58.out
rlabel metal2 20746 46172 20746 46172 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16698 47226 16698 47226 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24058 53142 24058 53142 0 sb_1__0_.mux_top_track_6.out
rlabel metal2 37490 44812 37490 44812 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39238 45390 39238 45390 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32890 41242 32890 41242 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37444 45254 37444 45254 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 33626 45594 33626 45594 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33074 48212 33074 48212 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24150 52326 24150 52326 0 sb_1__0_.mux_top_track_8.out
rlabel metal1 37904 44914 37904 44914 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 39698 44642 39698 44642 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31878 40018 31878 40018 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36938 44506 36938 44506 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35604 44506 35604 44506 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 35834 44217 35834 44217 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45402 55413 45402 55413 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 46046 55711 46046 55711 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46736 53550 46736 53550 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 47564 54162 47564 54162 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal2 47978 55711 47978 55711 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48668 53550 48668 53550 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44206 53550 44206 53550 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 44988 54162 44988 54162 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal3 3787 52156 3787 52156 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 2154 52972 2154 52972 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1211 53788 1211 53788 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 2062 54604 2062 54604 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 57000
<< end >>
