magic
tech sky130A
magscale 1 2
timestamp 1681685501
<< viali >>
rect 9137 24361 9171 24395
rect 37933 24361 37967 24395
rect 42441 24361 42475 24395
rect 44741 24361 44775 24395
rect 46857 24361 46891 24395
rect 23857 24293 23891 24327
rect 36921 24293 36955 24327
rect 39405 24293 39439 24327
rect 47961 24293 47995 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 16865 24225 16899 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25053 24225 25087 24259
rect 25237 24225 25271 24259
rect 26341 24225 26375 24259
rect 27721 24225 27755 24259
rect 29745 24225 29779 24259
rect 31677 24225 31711 24259
rect 2053 24157 2087 24191
rect 3893 24157 3927 24191
rect 4169 24157 4203 24191
rect 4629 24157 4663 24191
rect 6469 24157 6503 24191
rect 6745 24157 6779 24191
rect 7297 24157 7331 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 11897 24157 11931 24191
rect 12449 24157 12483 24191
rect 14473 24157 14507 24191
rect 15117 24157 15151 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22017 24157 22051 24191
rect 24041 24157 24075 24191
rect 27629 24157 27663 24191
rect 28549 24157 28583 24191
rect 30021 24157 30055 24191
rect 31033 24157 31067 24191
rect 32321 24157 32355 24191
rect 33425 24157 33459 24191
rect 34897 24157 34931 24191
rect 36001 24157 36035 24191
rect 37657 24157 37691 24191
rect 38485 24157 38519 24191
rect 40049 24157 40083 24191
rect 41153 24157 41187 24191
rect 42073 24157 42107 24191
rect 44373 24157 44407 24191
rect 45201 24157 45235 24191
rect 45937 24157 45971 24191
rect 46673 24157 46707 24191
rect 47225 24157 47259 24191
rect 47777 24157 47811 24191
rect 48605 24157 48639 24191
rect 17141 24089 17175 24123
rect 19073 24089 19107 24123
rect 34345 24089 34379 24123
rect 38117 24089 38151 24123
rect 39589 24089 39623 24123
rect 1593 24021 1627 24055
rect 1685 24021 1719 24055
rect 3985 24021 4019 24055
rect 6561 24021 6595 24055
rect 11713 24021 11747 24055
rect 14289 24021 14323 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 25789 24021 25823 24055
rect 26157 24021 26191 24055
rect 26249 24021 26283 24055
rect 27169 24021 27203 24055
rect 27537 24021 27571 24055
rect 28273 24021 28307 24055
rect 29193 24021 29227 24055
rect 32965 24021 32999 24055
rect 34069 24021 34103 24055
rect 35541 24021 35575 24055
rect 36645 24021 36679 24055
rect 37473 24021 37507 24055
rect 39129 24021 39163 24055
rect 40693 24021 40727 24055
rect 41797 24021 41831 24055
rect 44189 24021 44223 24055
rect 45385 24021 45419 24055
rect 46121 24021 46155 24055
rect 49249 24021 49283 24055
rect 1777 23817 1811 23851
rect 6469 23817 6503 23851
rect 12357 23817 12391 23851
rect 24225 23817 24259 23851
rect 36645 23817 36679 23851
rect 39313 23817 39347 23851
rect 41061 23817 41095 23851
rect 46305 23817 46339 23851
rect 47593 23817 47627 23851
rect 48145 23817 48179 23851
rect 3985 23749 4019 23783
rect 7205 23749 7239 23783
rect 9137 23749 9171 23783
rect 10977 23749 11011 23783
rect 14289 23749 14323 23783
rect 17877 23749 17911 23783
rect 21189 23749 21223 23783
rect 30665 23749 30699 23783
rect 33517 23749 33551 23783
rect 33701 23749 33735 23783
rect 36001 23749 36035 23783
rect 36185 23749 36219 23783
rect 37933 23749 37967 23783
rect 38485 23749 38519 23783
rect 38669 23749 38703 23783
rect 39221 23749 39255 23783
rect 43269 23749 43303 23783
rect 46213 23749 46247 23783
rect 2145 23681 2179 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6561 23681 6595 23715
rect 7113 23681 7147 23715
rect 7941 23681 7975 23715
rect 9873 23681 9907 23715
rect 12265 23681 12299 23715
rect 13277 23681 13311 23715
rect 15117 23681 15151 23715
rect 17049 23681 17083 23715
rect 18705 23681 18739 23715
rect 21005 23681 21039 23715
rect 29561 23681 29595 23715
rect 31493 23681 31527 23715
rect 32321 23681 32355 23715
rect 34345 23681 34379 23715
rect 34805 23681 34839 23715
rect 36829 23681 36863 23715
rect 37657 23681 37691 23715
rect 39957 23681 39991 23715
rect 40877 23681 40911 23715
rect 41429 23681 41463 23715
rect 42625 23681 42659 23715
rect 43729 23681 43763 23715
rect 44833 23681 44867 23715
rect 45569 23681 45603 23715
rect 46765 23681 46799 23715
rect 47317 23681 47351 23715
rect 47961 23681 47995 23715
rect 48697 23681 48731 23715
rect 5457 23613 5491 23647
rect 7389 23613 7423 23647
rect 12541 23613 12575 23647
rect 16129 23613 16163 23647
rect 18981 23613 19015 23647
rect 22017 23613 22051 23647
rect 22293 23613 22327 23647
rect 24869 23613 24903 23647
rect 25145 23613 25179 23647
rect 27169 23613 27203 23647
rect 27445 23613 27479 23647
rect 42073 23613 42107 23647
rect 6745 23545 6779 23579
rect 29377 23545 29411 23579
rect 30205 23545 30239 23579
rect 37473 23545 37507 23579
rect 1593 23477 1627 23511
rect 2237 23477 2271 23511
rect 11529 23477 11563 23511
rect 11897 23477 11931 23511
rect 20453 23477 20487 23511
rect 21649 23477 21683 23511
rect 23765 23477 23799 23511
rect 26617 23477 26651 23511
rect 28917 23477 28951 23511
rect 29929 23477 29963 23511
rect 30113 23477 30147 23511
rect 30757 23477 30791 23511
rect 31309 23477 31343 23511
rect 31861 23477 31895 23511
rect 32965 23477 32999 23511
rect 34161 23477 34195 23511
rect 35449 23477 35483 23511
rect 40601 23477 40635 23511
rect 44373 23477 44407 23511
rect 45017 23477 45051 23511
rect 45753 23477 45787 23511
rect 46949 23477 46983 23511
rect 49341 23477 49375 23511
rect 3617 23273 3651 23307
rect 3801 23273 3835 23307
rect 11069 23273 11103 23307
rect 11786 23273 11820 23307
rect 13645 23273 13679 23307
rect 13921 23273 13955 23307
rect 19441 23273 19475 23307
rect 25789 23273 25823 23307
rect 29009 23273 29043 23307
rect 29377 23273 29411 23307
rect 33609 23273 33643 23307
rect 34161 23273 34195 23307
rect 39589 23273 39623 23307
rect 44005 23273 44039 23307
rect 44649 23273 44683 23307
rect 49341 23273 49375 23307
rect 14933 23205 14967 23239
rect 18889 23205 18923 23239
rect 3433 23137 3467 23171
rect 4813 23137 4847 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11529 23137 11563 23171
rect 13277 23137 13311 23171
rect 16497 23137 16531 23171
rect 20085 23137 20119 23171
rect 22569 23137 22603 23171
rect 25145 23137 25179 23171
rect 26341 23137 26375 23171
rect 27261 23137 27295 23171
rect 27537 23137 27571 23171
rect 30021 23137 30055 23171
rect 31493 23137 31527 23171
rect 40049 23137 40083 23171
rect 47501 23137 47535 23171
rect 1777 23069 1811 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9321 23069 9355 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 19625 23069 19659 23103
rect 22293 23069 22327 23103
rect 26249 23069 26283 23103
rect 29745 23069 29779 23103
rect 32137 23069 32171 23103
rect 33149 23069 33183 23103
rect 34069 23069 34103 23103
rect 34989 23069 35023 23103
rect 38945 23069 38979 23103
rect 39221 23069 39255 23103
rect 40325 23069 40359 23103
rect 42901 23069 42935 23103
rect 43361 23069 43395 23103
rect 46213 23069 46247 23103
rect 47685 23069 47719 23103
rect 47961 23069 47995 23103
rect 48697 23069 48731 23103
rect 2789 23001 2823 23035
rect 4077 23001 4111 23035
rect 4537 23001 4571 23035
rect 9597 23001 9631 23035
rect 14381 23001 14415 23035
rect 17417 23001 17451 23035
rect 20361 23001 20395 23035
rect 25053 23001 25087 23035
rect 33425 23001 33459 23035
rect 35173 23001 35207 23035
rect 35633 23001 35667 23035
rect 36553 23001 36587 23035
rect 4169 22933 4203 22967
rect 4629 22933 4663 22967
rect 9045 22933 9079 22967
rect 14473 22933 14507 22967
rect 21833 22933 21867 22967
rect 24041 22933 24075 22967
rect 24593 22933 24627 22967
rect 24961 22933 24995 22967
rect 26157 22933 26191 22967
rect 26893 22933 26927 22967
rect 31953 22933 31987 22967
rect 32413 22933 32447 22967
rect 32597 22933 32631 22967
rect 32965 22933 32999 22967
rect 36093 22933 36127 22967
rect 37841 22933 37875 22967
rect 38761 22933 38795 22967
rect 42717 22933 42751 22967
rect 46857 22933 46891 22967
rect 48145 22933 48179 22967
rect 18613 22729 18647 22763
rect 21465 22729 21499 22763
rect 25789 22729 25823 22763
rect 26433 22729 26467 22763
rect 27629 22729 27663 22763
rect 31033 22729 31067 22763
rect 33241 22729 33275 22763
rect 36829 22729 36863 22763
rect 37473 22729 37507 22763
rect 43269 22729 43303 22763
rect 47777 22729 47811 22763
rect 10701 22661 10735 22695
rect 16129 22661 16163 22695
rect 17141 22661 17175 22695
rect 22201 22661 22235 22695
rect 26525 22661 26559 22695
rect 26801 22661 26835 22695
rect 28641 22661 28675 22695
rect 33793 22661 33827 22695
rect 36553 22661 36587 22695
rect 41797 22661 41831 22695
rect 47685 22661 47719 22695
rect 1777 22593 1811 22627
rect 3801 22593 3835 22627
rect 4813 22593 4847 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 7941 22593 7975 22627
rect 9781 22593 9815 22627
rect 11805 22593 11839 22627
rect 14565 22593 14599 22627
rect 15025 22593 15059 22627
rect 19257 22593 19291 22627
rect 19717 22593 19751 22627
rect 22477 22593 22511 22627
rect 25697 22593 25731 22627
rect 27537 22593 27571 22627
rect 30941 22593 30975 22627
rect 31861 22593 31895 22627
rect 32413 22593 32447 22627
rect 33149 22593 33183 22627
rect 34253 22593 34287 22627
rect 34529 22593 34563 22627
rect 35633 22593 35667 22627
rect 36369 22593 36403 22627
rect 37381 22593 37415 22627
rect 37841 22593 37875 22627
rect 40877 22593 40911 22627
rect 41521 22593 41555 22627
rect 42625 22593 42659 22627
rect 43913 22593 43947 22627
rect 48053 22593 48087 22627
rect 48329 22593 48363 22627
rect 49065 22593 49099 22627
rect 2789 22525 2823 22559
rect 3893 22525 3927 22559
rect 4077 22525 4111 22559
rect 5089 22525 5123 22559
rect 7297 22525 7331 22559
rect 8677 22525 8711 22559
rect 12449 22525 12483 22559
rect 12725 22525 12759 22559
rect 16865 22525 16899 22559
rect 19993 22525 20027 22559
rect 21925 22525 21959 22559
rect 23121 22525 23155 22559
rect 23397 22525 23431 22559
rect 25881 22525 25915 22559
rect 27721 22525 27755 22559
rect 28365 22525 28399 22559
rect 30113 22525 30147 22559
rect 31125 22525 31159 22559
rect 33609 22525 33643 22559
rect 38117 22525 38151 22559
rect 44557 22525 44591 22559
rect 6745 22457 6779 22491
rect 27169 22457 27203 22491
rect 30573 22457 30607 22491
rect 31677 22457 31711 22491
rect 3433 22389 3467 22423
rect 6469 22389 6503 22423
rect 11897 22389 11931 22423
rect 14197 22389 14231 22423
rect 19073 22389 19107 22423
rect 24869 22389 24903 22423
rect 25329 22389 25363 22423
rect 32505 22389 32539 22423
rect 35725 22389 35759 22423
rect 39589 22389 39623 22423
rect 40693 22389 40727 22423
rect 41337 22389 41371 22423
rect 48513 22389 48547 22423
rect 49249 22389 49283 22423
rect 14473 22185 14507 22219
rect 27537 22185 27571 22219
rect 28641 22185 28675 22219
rect 29653 22185 29687 22219
rect 29837 22185 29871 22219
rect 9045 22117 9079 22151
rect 20085 22117 20119 22151
rect 22293 22117 22327 22151
rect 24593 22117 24627 22151
rect 48421 22117 48455 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 7297 22049 7331 22083
rect 9781 22049 9815 22083
rect 9965 22049 9999 22083
rect 11253 22049 11287 22083
rect 13369 22049 13403 22083
rect 15669 22049 15703 22083
rect 17141 22049 17175 22083
rect 22661 22049 22695 22083
rect 23765 22049 23799 22083
rect 23949 22049 23983 22083
rect 25237 22049 25271 22083
rect 29193 22049 29227 22083
rect 30757 22049 30791 22083
rect 31861 22049 31895 22083
rect 32045 22049 32079 22083
rect 32229 22049 32263 22083
rect 39221 22049 39255 22083
rect 1777 21981 1811 22015
rect 3617 21981 3651 22015
rect 3985 21981 4019 22015
rect 6285 21981 6319 22015
rect 6929 21981 6963 22015
rect 8769 21981 8803 22015
rect 10517 21981 10551 22015
rect 12541 21981 12575 22015
rect 14381 21981 14415 22015
rect 15209 21981 15243 22015
rect 20361 21981 20395 22015
rect 25789 21981 25823 22015
rect 28801 21977 28835 22011
rect 29285 21981 29319 22015
rect 30573 21981 30607 22015
rect 32597 21981 32631 22015
rect 32873 21981 32907 22015
rect 33977 21981 34011 22015
rect 34529 21981 34563 22015
rect 35817 21981 35851 22015
rect 37657 21981 37691 22015
rect 37933 21981 37967 22015
rect 38945 21981 38979 22015
rect 48605 21981 48639 22015
rect 49065 21981 49099 22015
rect 5825 21913 5859 21947
rect 8585 21913 8619 21947
rect 17417 21913 17451 21947
rect 19533 21913 19567 21947
rect 21281 21913 21315 21947
rect 24961 21913 24995 21947
rect 26065 21913 26099 21947
rect 31401 21913 31435 21947
rect 34989 21913 35023 21947
rect 3433 21845 3467 21879
rect 6101 21845 6135 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 14933 21845 14967 21879
rect 18889 21845 18923 21879
rect 19625 21845 19659 21879
rect 22109 21845 22143 21879
rect 23305 21845 23339 21879
rect 23673 21845 23707 21879
rect 25053 21845 25087 21879
rect 27997 21845 28031 21879
rect 30113 21845 30147 21879
rect 30481 21845 30515 21879
rect 31493 21845 31527 21879
rect 34069 21845 34103 21879
rect 35081 21845 35115 21879
rect 35633 21845 35667 21879
rect 36277 21845 36311 21879
rect 37473 21845 37507 21879
rect 38761 21845 38795 21879
rect 49249 21845 49283 21879
rect 9413 21641 9447 21675
rect 10333 21641 10367 21675
rect 10977 21641 11011 21675
rect 11161 21641 11195 21675
rect 16037 21641 16071 21675
rect 20821 21641 20855 21675
rect 21005 21641 21039 21675
rect 23029 21641 23063 21675
rect 25973 21641 26007 21675
rect 26709 21641 26743 21675
rect 27629 21641 27663 21675
rect 27721 21641 27755 21675
rect 7941 21573 7975 21607
rect 13369 21573 13403 21607
rect 23673 21573 23707 21607
rect 28733 21573 28767 21607
rect 31033 21573 31067 21607
rect 33977 21573 34011 21607
rect 35449 21573 35483 21607
rect 1593 21505 1627 21539
rect 3433 21505 3467 21539
rect 5641 21505 5675 21539
rect 7021 21505 7055 21539
rect 7665 21505 7699 21539
rect 10241 21505 10275 21539
rect 12173 21505 12207 21539
rect 13093 21505 13127 21539
rect 15945 21505 15979 21539
rect 16865 21505 16899 21539
rect 21281 21505 21315 21539
rect 22385 21505 22419 21539
rect 22477 21505 22511 21539
rect 23397 21505 23431 21539
rect 26065 21505 26099 21539
rect 31125 21505 31159 21539
rect 32413 21505 32447 21539
rect 33241 21505 33275 21539
rect 34529 21505 34563 21539
rect 47961 21505 47995 21539
rect 2053 21437 2087 21471
rect 4169 21437 4203 21471
rect 5733 21437 5767 21471
rect 5917 21437 5951 21471
rect 10517 21437 10551 21471
rect 12265 21437 12299 21471
rect 12449 21437 12483 21471
rect 16221 21437 16255 21471
rect 17325 21437 17359 21471
rect 18705 21437 18739 21471
rect 18981 21437 19015 21471
rect 22661 21437 22695 21471
rect 25145 21437 25179 21471
rect 26249 21437 26283 21471
rect 27813 21437 27847 21471
rect 28457 21437 28491 21471
rect 31217 21437 31251 21471
rect 49157 21437 49191 21471
rect 6561 21369 6595 21403
rect 15577 21369 15611 21403
rect 22017 21369 22051 21403
rect 31861 21369 31895 21403
rect 33517 21369 33551 21403
rect 34621 21369 34655 21403
rect 5273 21301 5307 21335
rect 6469 21301 6503 21335
rect 7113 21301 7147 21335
rect 9873 21301 9907 21335
rect 11345 21301 11379 21335
rect 11805 21301 11839 21335
rect 14841 21301 14875 21335
rect 15301 21301 15335 21335
rect 20453 21301 20487 21335
rect 25605 21301 25639 21335
rect 27261 21301 27295 21335
rect 30205 21301 30239 21335
rect 30665 21301 30699 21335
rect 31769 21301 31803 21335
rect 32505 21301 32539 21335
rect 33057 21301 33091 21335
rect 34069 21301 34103 21335
rect 34897 21301 34931 21335
rect 47593 21301 47627 21335
rect 3433 21097 3467 21131
rect 5089 21097 5123 21131
rect 7665 21097 7699 21131
rect 13737 21097 13771 21131
rect 14565 21097 14599 21131
rect 34253 21097 34287 21131
rect 49433 21097 49467 21131
rect 3617 21029 3651 21063
rect 21649 21029 21683 21063
rect 25697 21029 25731 21063
rect 32505 21029 32539 21063
rect 4261 20961 4295 20995
rect 5733 20961 5767 20995
rect 8401 20961 8435 20995
rect 9689 20961 9723 20995
rect 10977 20961 11011 20995
rect 12633 20961 12667 20995
rect 14289 20961 14323 20995
rect 15117 20961 15151 20995
rect 16221 20961 16255 20995
rect 16405 20961 16439 20995
rect 17417 20961 17451 20995
rect 17601 20961 17635 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 19717 20961 19751 20995
rect 22753 20961 22787 20995
rect 23765 20961 23799 20995
rect 23857 20961 23891 20995
rect 25329 20961 25363 20995
rect 26065 20961 26099 20995
rect 26341 20961 26375 20995
rect 28549 20961 28583 20995
rect 29745 20961 29779 20995
rect 30021 20961 30055 20995
rect 33149 20961 33183 20995
rect 33517 20961 33551 20995
rect 33609 20961 33643 20995
rect 1777 20893 1811 20927
rect 3985 20893 4019 20927
rect 5457 20893 5491 20927
rect 8217 20893 8251 20927
rect 8309 20893 8343 20927
rect 9321 20893 9355 20927
rect 11989 20893 12023 20927
rect 16129 20893 16163 20927
rect 18521 20893 18555 20927
rect 19441 20893 19475 20927
rect 22569 20893 22603 20927
rect 28273 20893 28307 20927
rect 31125 20893 31159 20927
rect 32689 20893 32723 20927
rect 32965 20893 32999 20927
rect 2789 20825 2823 20859
rect 11345 20825 11379 20859
rect 15025 20825 15059 20859
rect 21833 20825 21867 20859
rect 22477 20825 22511 20859
rect 25053 20825 25087 20859
rect 31861 20825 31895 20859
rect 32045 20825 32079 20859
rect 7205 20757 7239 20791
rect 7573 20757 7607 20791
rect 7849 20757 7883 20791
rect 11437 20757 11471 20791
rect 13921 20757 13955 20791
rect 14933 20757 14967 20791
rect 15761 20757 15795 20791
rect 16957 20757 16991 20791
rect 17325 20757 17359 20791
rect 18153 20757 18187 20791
rect 21189 20757 21223 20791
rect 22109 20757 22143 20791
rect 23305 20757 23339 20791
rect 23673 20757 23707 20791
rect 24685 20757 24719 20791
rect 25145 20757 25179 20791
rect 27813 20757 27847 20791
rect 31217 20757 31251 20791
rect 34069 20757 34103 20791
rect 5641 20553 5675 20587
rect 12909 20553 12943 20587
rect 13001 20553 13035 20587
rect 16129 20553 16163 20587
rect 17509 20553 17543 20587
rect 18521 20553 18555 20587
rect 18889 20553 18923 20587
rect 23397 20553 23431 20587
rect 24041 20553 24075 20587
rect 26525 20553 26559 20587
rect 27169 20553 27203 20587
rect 27629 20553 27663 20587
rect 30941 20553 30975 20587
rect 32873 20553 32907 20587
rect 8769 20485 8803 20519
rect 11805 20485 11839 20519
rect 14013 20485 14047 20519
rect 22017 20485 22051 20519
rect 22753 20485 22787 20519
rect 26433 20485 26467 20519
rect 31033 20485 31067 20519
rect 1777 20417 1811 20451
rect 3433 20417 3467 20451
rect 5733 20417 5767 20451
rect 6561 20417 6595 20451
rect 13737 20417 13771 20451
rect 16037 20417 16071 20451
rect 17417 20417 17451 20451
rect 19717 20417 19751 20451
rect 24317 20417 24351 20451
rect 26709 20417 26743 20451
rect 27537 20417 27571 20451
rect 32689 20417 32723 20451
rect 2053 20349 2087 20383
rect 3893 20349 3927 20383
rect 5917 20349 5951 20383
rect 7021 20349 7055 20383
rect 9413 20349 9447 20383
rect 9689 20349 9723 20383
rect 13185 20349 13219 20383
rect 16865 20349 16899 20383
rect 17693 20349 17727 20383
rect 18981 20349 19015 20383
rect 19073 20349 19107 20383
rect 19993 20349 20027 20383
rect 24593 20349 24627 20383
rect 26065 20349 26099 20383
rect 27721 20349 27755 20383
rect 28365 20349 28399 20383
rect 28641 20349 28675 20383
rect 31125 20349 31159 20383
rect 15485 20281 15519 20315
rect 17049 20281 17083 20315
rect 32321 20281 32355 20315
rect 5273 20213 5307 20247
rect 8309 20213 8343 20247
rect 8861 20213 8895 20247
rect 11161 20213 11195 20247
rect 11897 20213 11931 20247
rect 12541 20213 12575 20247
rect 13461 20213 13495 20247
rect 13645 20213 13679 20247
rect 16681 20213 16715 20247
rect 18153 20213 18187 20247
rect 21465 20213 21499 20247
rect 30113 20213 30147 20247
rect 30573 20213 30607 20247
rect 31585 20213 31619 20247
rect 31769 20213 31803 20247
rect 32137 20213 32171 20247
rect 32505 20213 32539 20247
rect 3525 20009 3559 20043
rect 3985 20009 4019 20043
rect 4169 20009 4203 20043
rect 6285 20009 6319 20043
rect 10885 20009 10919 20043
rect 13001 20009 13035 20043
rect 18705 20009 18739 20043
rect 27629 20009 27663 20043
rect 29745 20009 29779 20043
rect 30205 20009 30239 20043
rect 31861 20009 31895 20043
rect 14289 19941 14323 19975
rect 14473 19941 14507 19975
rect 16773 19941 16807 19975
rect 17233 19941 17267 19975
rect 4537 19873 4571 19907
rect 6745 19873 6779 19907
rect 9137 19873 9171 19907
rect 11345 19873 11379 19907
rect 11437 19873 11471 19907
rect 12357 19873 12391 19907
rect 13461 19873 13495 19907
rect 13645 19873 13679 19907
rect 14841 19873 14875 19907
rect 17877 19873 17911 19907
rect 20545 19873 20579 19907
rect 22017 19873 22051 19907
rect 23857 19873 23891 19907
rect 25329 19873 25363 19907
rect 28641 19873 28675 19907
rect 31309 19873 31343 19907
rect 1777 19805 1811 19839
rect 12173 19805 12207 19839
rect 14565 19805 14599 19839
rect 17693 19805 17727 19839
rect 18889 19805 18923 19839
rect 20269 19805 20303 19839
rect 22569 19805 22603 19839
rect 23765 19805 23799 19839
rect 25881 19805 25915 19839
rect 28365 19805 28399 19839
rect 29929 19805 29963 19839
rect 31217 19805 31251 19839
rect 2789 19737 2823 19771
rect 4813 19737 4847 19771
rect 7021 19737 7055 19771
rect 9413 19737 9447 19771
rect 13369 19737 13403 19771
rect 16957 19737 16991 19771
rect 19625 19737 19659 19771
rect 26157 19737 26191 19771
rect 3433 19669 3467 19703
rect 3893 19669 3927 19703
rect 8493 19669 8527 19703
rect 11805 19669 11839 19703
rect 12265 19669 12299 19703
rect 13829 19669 13863 19703
rect 16313 19669 16347 19703
rect 17601 19669 17635 19703
rect 18429 19669 18463 19703
rect 19717 19669 19751 19703
rect 22661 19669 22695 19703
rect 23305 19669 23339 19703
rect 23673 19669 23707 19703
rect 24685 19669 24719 19703
rect 25053 19669 25087 19703
rect 25145 19669 25179 19703
rect 27905 19669 27939 19703
rect 30389 19669 30423 19703
rect 30757 19669 30791 19703
rect 31125 19669 31159 19703
rect 5273 19465 5307 19499
rect 5733 19465 5767 19499
rect 10425 19465 10459 19499
rect 14841 19465 14875 19499
rect 17233 19465 17267 19499
rect 17877 19465 17911 19499
rect 19073 19465 19107 19499
rect 21465 19465 21499 19499
rect 22385 19465 22419 19499
rect 26433 19465 26467 19499
rect 27721 19465 27755 19499
rect 30481 19465 30515 19499
rect 4353 19397 4387 19431
rect 9321 19397 9355 19431
rect 18337 19397 18371 19431
rect 22477 19397 22511 19431
rect 24041 19397 24075 19431
rect 1777 19329 1811 19363
rect 2789 19329 2823 19363
rect 3617 19329 3651 19363
rect 5641 19329 5675 19363
rect 6561 19329 6595 19363
rect 7481 19329 7515 19363
rect 8585 19329 8619 19363
rect 10333 19329 10367 19363
rect 10793 19329 10827 19363
rect 10885 19329 10919 19363
rect 11713 19329 11747 19363
rect 14749 19329 14783 19363
rect 15669 19329 15703 19363
rect 17417 19329 17451 19363
rect 18245 19329 18279 19363
rect 19257 19329 19291 19363
rect 24133 19329 24167 19363
rect 24961 19329 24995 19363
rect 30665 19329 30699 19363
rect 31125 19329 31159 19363
rect 5917 19261 5951 19295
rect 10977 19261 11011 19295
rect 11989 19261 12023 19295
rect 14933 19261 14967 19295
rect 18429 19261 18463 19295
rect 19717 19261 19751 19295
rect 22661 19261 22695 19295
rect 24317 19261 24351 19295
rect 25789 19261 25823 19295
rect 26985 19261 27019 19295
rect 27445 19261 27479 19295
rect 27905 19261 27939 19295
rect 28273 19261 28307 19295
rect 10149 19193 10183 19227
rect 13737 19193 13771 19227
rect 13829 19193 13863 19227
rect 14381 19193 14415 19227
rect 15853 19193 15887 19227
rect 23305 19193 23339 19227
rect 13461 19125 13495 19159
rect 14013 19125 14047 19159
rect 14197 19125 14231 19159
rect 15209 19125 15243 19159
rect 15393 19125 15427 19159
rect 16037 19125 16071 19159
rect 16221 19125 16255 19159
rect 16405 19125 16439 19159
rect 16681 19125 16715 19159
rect 16865 19125 16899 19159
rect 17049 19125 17083 19159
rect 17509 19125 17543 19159
rect 17693 19125 17727 19159
rect 19980 19125 20014 19159
rect 22017 19125 22051 19159
rect 23121 19125 23155 19159
rect 23673 19125 23707 19159
rect 27261 19125 27295 19159
rect 28530 19125 28564 19159
rect 30021 19125 30055 19159
rect 30941 19125 30975 19159
rect 3893 18921 3927 18955
rect 11621 18921 11655 18955
rect 14657 18921 14691 18955
rect 14933 18921 14967 18955
rect 22937 18921 22971 18955
rect 27169 18921 27203 18955
rect 8585 18853 8619 18887
rect 14197 18853 14231 18887
rect 23397 18853 23431 18887
rect 2053 18785 2087 18819
rect 3985 18785 4019 18819
rect 6837 18785 6871 18819
rect 10057 18785 10091 18819
rect 11161 18785 11195 18819
rect 12173 18785 12207 18819
rect 13553 18785 13587 18819
rect 13921 18785 13955 18819
rect 15209 18785 15243 18819
rect 17509 18785 17543 18819
rect 18613 18785 18647 18819
rect 18705 18785 18739 18819
rect 20361 18785 20395 18819
rect 21189 18785 21223 18819
rect 21465 18785 21499 18819
rect 24593 18785 24627 18819
rect 25421 18785 25455 18819
rect 30297 18785 30331 18819
rect 1777 18717 1811 18751
rect 4629 18717 4663 18751
rect 9873 18717 9907 18751
rect 10977 18717 11011 18751
rect 14565 18717 14599 18751
rect 19625 18717 19659 18751
rect 23581 18717 23615 18751
rect 25053 18717 25087 18751
rect 27629 18717 27663 18751
rect 27905 18717 27939 18751
rect 30205 18717 30239 18751
rect 4905 18649 4939 18683
rect 7113 18649 7147 18683
rect 9137 18649 9171 18683
rect 12817 18649 12851 18683
rect 15485 18649 15519 18683
rect 25697 18649 25731 18683
rect 30757 18649 30791 18683
rect 3341 18581 3375 18615
rect 3617 18581 3651 18615
rect 6377 18581 6411 18615
rect 9413 18581 9447 18615
rect 9781 18581 9815 18615
rect 10609 18581 10643 18615
rect 11989 18581 12023 18615
rect 12081 18581 12115 18615
rect 15117 18581 15151 18615
rect 16957 18581 16991 18615
rect 18153 18581 18187 18615
rect 18521 18581 18555 18615
rect 19349 18581 19383 18615
rect 20821 18581 20855 18615
rect 23949 18581 23983 18615
rect 24133 18581 24167 18615
rect 29745 18581 29779 18615
rect 30113 18581 30147 18615
rect 15393 18377 15427 18411
rect 16313 18377 16347 18411
rect 17325 18377 17359 18411
rect 20729 18377 20763 18411
rect 24869 18377 24903 18411
rect 27169 18377 27203 18411
rect 30665 18377 30699 18411
rect 31309 18377 31343 18411
rect 7757 18309 7791 18343
rect 14473 18309 14507 18343
rect 18153 18309 18187 18343
rect 22017 18309 22051 18343
rect 22569 18309 22603 18343
rect 22845 18309 22879 18343
rect 25329 18309 25363 18343
rect 26065 18309 26099 18343
rect 28365 18309 28399 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 5641 18241 5675 18275
rect 6745 18241 6779 18275
rect 8493 18241 8527 18275
rect 9229 18241 9263 18275
rect 10793 18241 10827 18275
rect 11713 18241 11747 18275
rect 12357 18241 12391 18275
rect 13185 18241 13219 18275
rect 13645 18241 13679 18275
rect 16497 18241 16531 18275
rect 17233 18241 17267 18275
rect 18337 18241 18371 18275
rect 19901 18241 19935 18275
rect 19993 18241 20027 18275
rect 21097 18241 21131 18275
rect 26525 18241 26559 18275
rect 28089 18241 28123 18275
rect 30757 18241 30791 18275
rect 31493 18241 31527 18275
rect 2053 18173 2087 18207
rect 3893 18173 3927 18207
rect 5733 18173 5767 18207
rect 5917 18173 5951 18207
rect 9873 18173 9907 18207
rect 10885 18173 10919 18207
rect 11069 18173 11103 18207
rect 12449 18173 12483 18207
rect 12541 18173 12575 18207
rect 15485 18173 15519 18207
rect 15669 18173 15703 18207
rect 17509 18173 17543 18207
rect 18889 18173 18923 18207
rect 20085 18173 20119 18207
rect 21189 18173 21223 18207
rect 21373 18173 21407 18207
rect 23121 18173 23155 18207
rect 23397 18173 23431 18207
rect 30849 18173 30883 18207
rect 10425 18105 10459 18139
rect 15025 18105 15059 18139
rect 19533 18105 19567 18139
rect 30297 18105 30331 18139
rect 5273 18037 5307 18071
rect 9689 18037 9723 18071
rect 10057 18037 10091 18071
rect 11989 18037 12023 18071
rect 13369 18037 13403 18071
rect 16037 18037 16071 18071
rect 16865 18037 16899 18071
rect 26709 18037 26743 18071
rect 29837 18037 29871 18071
rect 3617 17833 3651 17867
rect 10609 17833 10643 17867
rect 26617 17833 26651 17867
rect 27334 17833 27368 17867
rect 29101 17833 29135 17867
rect 31953 17833 31987 17867
rect 4445 17765 4479 17799
rect 6653 17765 6687 17799
rect 7849 17765 7883 17799
rect 13737 17765 13771 17799
rect 16037 17765 16071 17799
rect 29745 17765 29779 17799
rect 7389 17697 7423 17731
rect 8401 17697 8435 17731
rect 9873 17697 9907 17731
rect 11161 17697 11195 17731
rect 16313 17697 16347 17731
rect 16589 17697 16623 17731
rect 19441 17697 19475 17731
rect 19717 17697 19751 17731
rect 21281 17697 21315 17731
rect 24869 17697 24903 17731
rect 27077 17697 27111 17731
rect 30205 17697 30239 17731
rect 30297 17697 30331 17731
rect 31493 17697 31527 17731
rect 1777 17629 1811 17663
rect 4905 17629 4939 17663
rect 8217 17629 8251 17663
rect 9137 17629 9171 17663
rect 10977 17629 11011 17663
rect 11989 17629 12023 17663
rect 18337 17629 18371 17663
rect 21741 17629 21775 17663
rect 22293 17629 22327 17663
rect 31309 17629 31343 17663
rect 2513 17561 2547 17595
rect 4261 17561 4295 17595
rect 5181 17561 5215 17595
rect 7205 17561 7239 17595
rect 8309 17561 8343 17595
rect 11069 17561 11103 17595
rect 12265 17561 12299 17595
rect 14381 17561 14415 17595
rect 21097 17561 21131 17595
rect 22569 17561 22603 17595
rect 25145 17561 25179 17595
rect 30113 17561 30147 17595
rect 31401 17561 31435 17595
rect 3433 17493 3467 17527
rect 3801 17493 3835 17527
rect 11621 17493 11655 17527
rect 14473 17493 14507 17527
rect 14933 17493 14967 17527
rect 15117 17493 15151 17527
rect 15393 17493 15427 17527
rect 18061 17493 18095 17527
rect 18705 17493 18739 17527
rect 20729 17493 20763 17527
rect 21189 17493 21223 17527
rect 21925 17493 21959 17527
rect 24041 17493 24075 17527
rect 24409 17493 24443 17527
rect 28825 17493 28859 17527
rect 30941 17493 30975 17527
rect 5273 17289 5307 17323
rect 7297 17289 7331 17323
rect 8033 17289 8067 17323
rect 8493 17289 8527 17323
rect 9505 17289 9539 17323
rect 9965 17289 9999 17323
rect 12541 17289 12575 17323
rect 12909 17289 12943 17323
rect 13737 17289 13771 17323
rect 15025 17289 15059 17323
rect 23673 17289 23707 17323
rect 29837 17289 29871 17323
rect 30573 17289 30607 17323
rect 4445 17221 4479 17255
rect 10977 17221 11011 17255
rect 13001 17221 13035 17255
rect 18429 17221 18463 17255
rect 20361 17221 20395 17255
rect 22477 17221 22511 17255
rect 23765 17221 23799 17255
rect 24317 17221 24351 17255
rect 24961 17221 24995 17255
rect 30849 17221 30883 17255
rect 1777 17153 1811 17187
rect 3617 17153 3651 17187
rect 5641 17153 5675 17187
rect 7205 17153 7239 17187
rect 8401 17153 8435 17187
rect 9137 17153 9171 17187
rect 9873 17153 9907 17187
rect 10793 17153 10827 17187
rect 11805 17153 11839 17187
rect 14105 17153 14139 17187
rect 15209 17153 15243 17187
rect 15669 17153 15703 17187
rect 16313 17153 16347 17187
rect 17233 17153 17267 17187
rect 21097 17153 21131 17187
rect 22385 17153 22419 17187
rect 24685 17153 24719 17187
rect 27813 17153 27847 17187
rect 2053 17085 2087 17119
rect 5733 17085 5767 17119
rect 5825 17085 5859 17119
rect 7389 17085 7423 17119
rect 8677 17085 8711 17119
rect 10057 17085 10091 17119
rect 13093 17085 13127 17119
rect 14197 17085 14231 17119
rect 14381 17085 14415 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 18153 17085 18187 17119
rect 20269 17085 20303 17119
rect 21189 17085 21223 17119
rect 21373 17085 21407 17119
rect 22569 17085 22603 17119
rect 23857 17085 23891 17119
rect 26433 17085 26467 17119
rect 27169 17085 27203 17119
rect 28089 17085 28123 17119
rect 6469 17017 6503 17051
rect 6837 17017 6871 17051
rect 11989 17017 12023 17051
rect 14749 17017 14783 17051
rect 16129 17017 16163 17051
rect 11345 16949 11379 16983
rect 15485 16949 15519 16983
rect 16865 16949 16899 16983
rect 19901 16949 19935 16983
rect 20729 16949 20763 16983
rect 22017 16949 22051 16983
rect 23305 16949 23339 16983
rect 26709 16949 26743 16983
rect 29561 16949 29595 16983
rect 3617 16745 3651 16779
rect 6009 16745 6043 16779
rect 12541 16745 12575 16779
rect 12633 16745 12667 16779
rect 16129 16745 16163 16779
rect 16405 16745 16439 16779
rect 10057 16677 10091 16711
rect 12357 16677 12391 16711
rect 25697 16677 25731 16711
rect 25973 16677 26007 16711
rect 3341 16609 3375 16643
rect 7113 16609 7147 16643
rect 7297 16609 7331 16643
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 10701 16609 10735 16643
rect 11897 16609 11931 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 15485 16609 15519 16643
rect 15669 16609 15703 16643
rect 16773 16609 16807 16643
rect 19717 16609 19751 16643
rect 22477 16609 22511 16643
rect 22569 16609 22603 16643
rect 23765 16609 23799 16643
rect 25145 16609 25179 16643
rect 25329 16609 25363 16643
rect 27077 16609 27111 16643
rect 27169 16609 27203 16643
rect 28273 16609 28307 16643
rect 28457 16609 28491 16643
rect 28917 16609 28951 16643
rect 1777 16541 1811 16575
rect 4077 16541 4111 16575
rect 5181 16541 5215 16575
rect 9413 16541 9447 16575
rect 10517 16541 10551 16575
rect 11621 16541 11655 16575
rect 14565 16541 14599 16575
rect 15393 16541 15427 16575
rect 17601 16541 17635 16575
rect 18245 16541 18279 16575
rect 19441 16541 19475 16575
rect 22385 16541 22419 16575
rect 23581 16541 23615 16575
rect 28181 16541 28215 16575
rect 2513 16473 2547 16507
rect 5917 16473 5951 16507
rect 9229 16473 9263 16507
rect 13369 16473 13403 16507
rect 21465 16473 21499 16507
rect 23673 16473 23707 16507
rect 26985 16473 27019 16507
rect 6653 16405 6687 16439
rect 7021 16405 7055 16439
rect 7849 16405 7883 16439
rect 8217 16405 8251 16439
rect 9781 16405 9815 16439
rect 10425 16405 10459 16439
rect 11253 16405 11287 16439
rect 11713 16405 11747 16439
rect 13001 16405 13035 16439
rect 14381 16405 14415 16439
rect 15025 16405 15059 16439
rect 16221 16405 16255 16439
rect 17417 16405 17451 16439
rect 18061 16405 18095 16439
rect 18705 16405 18739 16439
rect 22017 16405 22051 16439
rect 23213 16405 23247 16439
rect 24685 16405 24719 16439
rect 25053 16405 25087 16439
rect 26617 16405 26651 16439
rect 27813 16405 27847 16439
rect 7297 16201 7331 16235
rect 11621 16201 11655 16235
rect 13737 16201 13771 16235
rect 17141 16201 17175 16235
rect 20453 16201 20487 16235
rect 21281 16201 21315 16235
rect 26617 16201 26651 16235
rect 4353 16133 4387 16167
rect 8769 16133 8803 16167
rect 10609 16133 10643 16167
rect 14657 16133 14691 16167
rect 16957 16133 16991 16167
rect 17877 16133 17911 16167
rect 1777 16065 1811 16099
rect 3525 16065 3559 16099
rect 5641 16065 5675 16099
rect 5733 16065 5767 16099
rect 7665 16065 7699 16099
rect 7757 16065 7791 16099
rect 8493 16065 8527 16099
rect 11161 16065 11195 16099
rect 11989 16065 12023 16099
rect 14749 16065 14783 16099
rect 16313 16065 16347 16099
rect 17785 16065 17819 16099
rect 18613 16065 18647 16099
rect 19717 16065 19751 16099
rect 20545 16065 20579 16099
rect 21465 16065 21499 16099
rect 22293 16065 22327 16099
rect 23673 16065 23707 16099
rect 24317 16065 24351 16099
rect 24593 16065 24627 16099
rect 24869 16065 24903 16099
rect 26985 16065 27019 16099
rect 2053 15997 2087 16031
rect 5917 15997 5951 16031
rect 6653 15997 6687 16031
rect 7849 15997 7883 16031
rect 10241 15997 10275 16031
rect 12265 15997 12299 16031
rect 14841 15997 14875 16031
rect 15485 15997 15519 16031
rect 16773 15997 16807 16031
rect 17969 15997 18003 16031
rect 18889 15997 18923 16031
rect 20729 15997 20763 16031
rect 22017 15997 22051 16031
rect 23765 15997 23799 16031
rect 23949 15997 23983 16031
rect 25145 15997 25179 16031
rect 10977 15929 11011 15963
rect 17417 15929 17451 15963
rect 5273 15861 5307 15895
rect 14289 15861 14323 15895
rect 16129 15861 16163 15895
rect 20085 15861 20119 15895
rect 23305 15861 23339 15895
rect 3433 15657 3467 15691
rect 9321 15657 9355 15691
rect 15853 15657 15887 15691
rect 19441 15657 19475 15691
rect 19901 15657 19935 15691
rect 22569 15657 22603 15691
rect 24501 15657 24535 15691
rect 3617 15589 3651 15623
rect 7849 15589 7883 15623
rect 10885 15589 10919 15623
rect 12081 15589 12115 15623
rect 26433 15589 26467 15623
rect 2053 15521 2087 15555
rect 4445 15521 4479 15555
rect 4629 15521 4663 15555
rect 5641 15521 5675 15555
rect 5825 15521 5859 15555
rect 6837 15521 6871 15555
rect 6929 15521 6963 15555
rect 8309 15521 8343 15555
rect 8401 15521 8435 15555
rect 10241 15521 10275 15555
rect 11437 15521 11471 15555
rect 12725 15521 12759 15555
rect 14105 15521 14139 15555
rect 15025 15521 15059 15555
rect 16497 15521 16531 15555
rect 20269 15521 20303 15555
rect 25697 15521 25731 15555
rect 25789 15521 25823 15555
rect 1777 15453 1811 15487
rect 12449 15453 12483 15487
rect 13277 15453 13311 15487
rect 13737 15453 13771 15487
rect 14841 15453 14875 15487
rect 17049 15453 17083 15487
rect 19625 15453 19659 15487
rect 22845 15453 22879 15487
rect 23121 15453 23155 15487
rect 25605 15453 25639 15487
rect 26341 15453 26375 15487
rect 5549 15385 5583 15419
rect 6745 15385 6779 15419
rect 9229 15385 9263 15419
rect 11253 15385 11287 15419
rect 14933 15385 14967 15419
rect 17325 15385 17359 15419
rect 20545 15385 20579 15419
rect 23949 15385 23983 15419
rect 3985 15317 4019 15351
rect 4353 15317 4387 15351
rect 5181 15317 5215 15351
rect 6377 15317 6411 15351
rect 7481 15317 7515 15351
rect 8217 15317 8251 15351
rect 9781 15317 9815 15351
rect 9965 15317 9999 15351
rect 11345 15317 11379 15351
rect 12541 15317 12575 15351
rect 13553 15317 13587 15351
rect 14473 15317 14507 15351
rect 15485 15317 15519 15351
rect 16221 15317 16255 15351
rect 16313 15317 16347 15351
rect 18797 15317 18831 15351
rect 22017 15317 22051 15351
rect 22385 15317 22419 15351
rect 25237 15317 25271 15351
rect 3525 15113 3559 15147
rect 6745 15113 6779 15147
rect 8677 15113 8711 15147
rect 9597 15113 9631 15147
rect 13001 15113 13035 15147
rect 18429 15113 18463 15147
rect 6653 15045 6687 15079
rect 9689 15045 9723 15079
rect 10793 15045 10827 15079
rect 14197 15045 14231 15079
rect 14841 15045 14875 15079
rect 19165 15045 19199 15079
rect 20177 15045 20211 15079
rect 22293 15045 22327 15079
rect 25145 15045 25179 15079
rect 1777 14977 1811 15011
rect 3709 14977 3743 15011
rect 4169 14977 4203 15011
rect 7665 14977 7699 15011
rect 8585 14977 8619 15011
rect 10885 14977 10919 15011
rect 11989 14977 12023 15011
rect 13369 14977 13403 15011
rect 13461 14977 13495 15011
rect 14013 14977 14047 15011
rect 17141 14977 17175 15011
rect 20085 14977 20119 15011
rect 22017 14977 22051 15011
rect 24869 14977 24903 15011
rect 2053 14909 2087 14943
rect 7757 14909 7791 14943
rect 7941 14909 7975 14943
rect 9873 14909 9907 14943
rect 10977 14909 11011 14943
rect 11713 14909 11747 14943
rect 13553 14909 13587 14943
rect 14565 14909 14599 14943
rect 20361 14909 20395 14943
rect 20913 14909 20947 14943
rect 24041 14909 24075 14943
rect 24225 14909 24259 14943
rect 26985 14909 27019 14943
rect 9229 14841 9263 14875
rect 19717 14841 19751 14875
rect 23765 14841 23799 14875
rect 4432 14773 4466 14807
rect 5917 14773 5951 14807
rect 7297 14773 7331 14807
rect 10425 14773 10459 14807
rect 16313 14773 16347 14807
rect 16681 14773 16715 14807
rect 19349 14773 19383 14807
rect 26617 14773 26651 14807
rect 13737 14569 13771 14603
rect 14105 14569 14139 14603
rect 14381 14569 14415 14603
rect 18613 14569 18647 14603
rect 26985 14569 27019 14603
rect 3985 14501 4019 14535
rect 11621 14501 11655 14535
rect 18889 14501 18923 14535
rect 21741 14501 21775 14535
rect 24041 14501 24075 14535
rect 2053 14433 2087 14467
rect 4905 14433 4939 14467
rect 7205 14433 7239 14467
rect 8493 14433 8527 14467
rect 9965 14433 9999 14467
rect 11161 14433 11195 14467
rect 12265 14433 12299 14467
rect 14933 14433 14967 14467
rect 16865 14433 16899 14467
rect 21097 14433 21131 14467
rect 22293 14433 22327 14467
rect 25145 14433 25179 14467
rect 26341 14433 26375 14467
rect 1777 14365 1811 14399
rect 4629 14365 4663 14399
rect 5457 14365 5491 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 9873 14365 9907 14399
rect 10977 14365 11011 14399
rect 11989 14365 12023 14399
rect 14657 14365 14691 14399
rect 19625 14365 19659 14399
rect 20913 14365 20947 14399
rect 21005 14365 21039 14399
rect 26157 14365 26191 14399
rect 5733 14297 5767 14331
rect 17141 14297 17175 14331
rect 21557 14297 21591 14331
rect 22569 14297 22603 14331
rect 24961 14297 24995 14331
rect 25053 14297 25087 14331
rect 26249 14297 26283 14331
rect 26801 14297 26835 14331
rect 3433 14229 3467 14263
rect 3617 14229 3651 14263
rect 4261 14229 4295 14263
rect 4721 14229 4755 14263
rect 7849 14229 7883 14263
rect 9045 14229 9079 14263
rect 9413 14229 9447 14263
rect 9781 14229 9815 14263
rect 10609 14229 10643 14263
rect 11069 14229 11103 14263
rect 16405 14229 16439 14263
rect 19441 14229 19475 14263
rect 20545 14229 20579 14263
rect 24593 14229 24627 14263
rect 25789 14229 25823 14263
rect 3433 14025 3467 14059
rect 4077 14025 4111 14059
rect 5641 14025 5675 14059
rect 6929 14025 6963 14059
rect 7297 14025 7331 14059
rect 8125 14025 8159 14059
rect 11989 14025 12023 14059
rect 13185 14025 13219 14059
rect 14381 14025 14415 14059
rect 14749 14025 14783 14059
rect 15577 14025 15611 14059
rect 18889 14025 18923 14059
rect 20085 14025 20119 14059
rect 23397 14025 23431 14059
rect 24961 14025 24995 14059
rect 4537 13957 4571 13991
rect 5733 13957 5767 13991
rect 8493 13957 8527 13991
rect 8585 13957 8619 13991
rect 11621 13957 11655 13991
rect 13645 13957 13679 13991
rect 16773 13957 16807 13991
rect 25053 13957 25087 13991
rect 25605 13957 25639 13991
rect 25881 13957 25915 13991
rect 1777 13889 1811 13923
rect 3617 13889 3651 13923
rect 4445 13889 4479 13923
rect 7389 13889 7423 13923
rect 12357 13889 12391 13923
rect 13553 13889 13587 13923
rect 15945 13889 15979 13923
rect 19625 13889 19659 13923
rect 20453 13889 20487 13923
rect 20545 13889 20579 13923
rect 21833 13889 21867 13923
rect 22569 13889 22603 13923
rect 22661 13889 22695 13923
rect 23765 13889 23799 13923
rect 2053 13821 2087 13855
rect 4721 13821 4755 13855
rect 5825 13821 5859 13855
rect 6377 13821 6411 13855
rect 7573 13821 7607 13855
rect 8677 13821 8711 13855
rect 9321 13821 9355 13855
rect 9597 13821 9631 13855
rect 11069 13821 11103 13855
rect 12449 13821 12483 13855
rect 12541 13821 12575 13855
rect 13829 13821 13863 13855
rect 14841 13821 14875 13855
rect 14933 13821 14967 13855
rect 16037 13821 16071 13855
rect 16221 13821 16255 13855
rect 17141 13821 17175 13855
rect 17417 13821 17451 13855
rect 20637 13821 20671 13855
rect 22845 13821 22879 13855
rect 23857 13821 23891 13855
rect 24041 13821 24075 13855
rect 25237 13821 25271 13855
rect 26157 13821 26191 13855
rect 6561 13753 6595 13787
rect 19441 13753 19475 13787
rect 22201 13753 22235 13787
rect 25973 13753 26007 13787
rect 5273 13685 5307 13719
rect 24593 13685 24627 13719
rect 6469 13481 6503 13515
rect 13737 13481 13771 13515
rect 16037 13481 16071 13515
rect 18889 13481 18923 13515
rect 20618 13481 20652 13515
rect 22109 13481 22143 13515
rect 23949 13481 23983 13515
rect 8493 13413 8527 13447
rect 11437 13413 11471 13447
rect 11713 13413 11747 13447
rect 22845 13413 22879 13447
rect 24133 13413 24167 13447
rect 2053 13345 2087 13379
rect 4169 13345 4203 13379
rect 6745 13345 6779 13379
rect 9413 13345 9447 13379
rect 10977 13345 11011 13379
rect 11989 13345 12023 13379
rect 14565 13345 14599 13379
rect 16497 13345 16531 13379
rect 17141 13345 17175 13379
rect 20361 13345 20395 13379
rect 23305 13345 23339 13379
rect 23489 13345 23523 13379
rect 1777 13277 1811 13311
rect 9137 13277 9171 13311
rect 10793 13277 10827 13311
rect 14289 13277 14323 13311
rect 22477 13277 22511 13311
rect 3525 13209 3559 13243
rect 4445 13209 4479 13243
rect 7021 13209 7055 13243
rect 12265 13209 12299 13243
rect 17417 13209 17451 13243
rect 23213 13209 23247 13243
rect 24593 13209 24627 13243
rect 25421 13209 25455 13243
rect 3433 13141 3467 13175
rect 3893 13141 3927 13175
rect 5917 13141 5951 13175
rect 6193 13141 6227 13175
rect 10425 13141 10459 13175
rect 10885 13141 10919 13175
rect 19349 13141 19383 13175
rect 19441 13141 19475 13175
rect 3893 12937 3927 12971
rect 7205 12937 7239 12971
rect 7297 12937 7331 12971
rect 12541 12937 12575 12971
rect 13737 12937 13771 12971
rect 14197 12937 14231 12971
rect 17785 12937 17819 12971
rect 18153 12937 18187 12971
rect 21097 12937 21131 12971
rect 22201 12937 22235 12971
rect 24777 12937 24811 12971
rect 4261 12869 4295 12903
rect 5733 12869 5767 12903
rect 10057 12869 10091 12903
rect 11897 12869 11931 12903
rect 15669 12869 15703 12903
rect 16129 12869 16163 12903
rect 16405 12869 16439 12903
rect 18981 12869 19015 12903
rect 1869 12801 1903 12835
rect 2881 12801 2915 12835
rect 4997 12801 5031 12835
rect 5641 12801 5675 12835
rect 6561 12801 6595 12835
rect 10701 12801 10735 12835
rect 12909 12801 12943 12835
rect 14105 12801 14139 12835
rect 14933 12801 14967 12835
rect 18245 12801 18279 12835
rect 21189 12801 21223 12835
rect 23029 12801 23063 12835
rect 1593 12733 1627 12767
rect 4813 12733 4847 12767
rect 5917 12733 5951 12767
rect 7389 12733 7423 12767
rect 8033 12733 8067 12767
rect 8309 12733 8343 12767
rect 13001 12733 13035 12767
rect 13185 12733 13219 12767
rect 14381 12733 14415 12767
rect 16865 12733 16899 12767
rect 18429 12733 18463 12767
rect 19809 12733 19843 12767
rect 21373 12733 21407 12767
rect 23305 12733 23339 12767
rect 4445 12665 4479 12699
rect 10517 12665 10551 12699
rect 11161 12665 11195 12699
rect 3525 12597 3559 12631
rect 5273 12597 5307 12631
rect 6837 12597 6871 12631
rect 11253 12597 11287 12631
rect 11621 12597 11655 12631
rect 20729 12597 20763 12631
rect 25053 12597 25087 12631
rect 3065 12393 3099 12427
rect 3525 12393 3559 12427
rect 4721 12393 4755 12427
rect 7849 12393 7883 12427
rect 11805 12393 11839 12427
rect 14381 12393 14415 12427
rect 18061 12393 18095 12427
rect 21833 12393 21867 12427
rect 4261 12325 4295 12359
rect 5365 12257 5399 12291
rect 8401 12257 8435 12291
rect 9873 12257 9907 12291
rect 11253 12257 11287 12291
rect 12265 12257 12299 12291
rect 12357 12257 12391 12291
rect 13645 12257 13679 12291
rect 16589 12257 16623 12291
rect 19073 12257 19107 12291
rect 20085 12257 20119 12291
rect 22569 12257 22603 12291
rect 1593 12189 1627 12223
rect 1869 12189 1903 12223
rect 4905 12189 4939 12223
rect 7389 12189 7423 12223
rect 8309 12189 8343 12223
rect 11069 12189 11103 12223
rect 13369 12189 13403 12223
rect 14105 12189 14139 12223
rect 15485 12189 15519 12223
rect 16313 12189 16347 12223
rect 18337 12189 18371 12223
rect 19533 12189 19567 12223
rect 22293 12189 22327 12223
rect 2973 12121 3007 12155
rect 4077 12121 4111 12155
rect 5641 12121 5675 12155
rect 9137 12121 9171 12155
rect 10977 12121 11011 12155
rect 12173 12121 12207 12155
rect 13461 12121 13495 12155
rect 14766 12121 14800 12155
rect 20361 12121 20395 12155
rect 8217 12053 8251 12087
rect 10609 12053 10643 12087
rect 13001 12053 13035 12087
rect 15945 12053 15979 12087
rect 18521 12053 18555 12087
rect 18797 12053 18831 12087
rect 19349 12053 19383 12087
rect 24041 12053 24075 12087
rect 24501 12053 24535 12087
rect 2237 11849 2271 11883
rect 4445 11849 4479 11883
rect 5273 11849 5307 11883
rect 5641 11849 5675 11883
rect 6745 11849 6779 11883
rect 12357 11849 12391 11883
rect 14933 11849 14967 11883
rect 17417 11849 17451 11883
rect 18153 11849 18187 11883
rect 18521 11849 18555 11883
rect 18613 11849 18647 11883
rect 19349 11849 19383 11883
rect 3801 11781 3835 11815
rect 5733 11781 5767 11815
rect 12449 11781 12483 11815
rect 16037 11781 16071 11815
rect 19165 11781 19199 11815
rect 21925 11781 21959 11815
rect 22661 11781 22695 11815
rect 1593 11713 1627 11747
rect 2697 11713 2731 11747
rect 4537 11713 4571 11747
rect 7389 11713 7423 11747
rect 9597 11713 9631 11747
rect 10977 11713 11011 11747
rect 13185 11713 13219 11747
rect 15945 11713 15979 11747
rect 17325 11713 17359 11747
rect 4721 11645 4755 11679
rect 5917 11645 5951 11679
rect 7665 11645 7699 11679
rect 10333 11645 10367 11679
rect 12541 11645 12575 11679
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 17509 11645 17543 11679
rect 18705 11645 18739 11679
rect 19717 11645 19751 11679
rect 19993 11645 20027 11679
rect 22385 11645 22419 11679
rect 24133 11645 24167 11679
rect 9137 11577 9171 11611
rect 11621 11577 11655 11611
rect 15577 11577 15611 11611
rect 3341 11509 3375 11543
rect 4077 11509 4111 11543
rect 6377 11509 6411 11543
rect 11989 11509 12023 11543
rect 15301 11509 15335 11543
rect 16957 11509 16991 11543
rect 21465 11509 21499 11543
rect 24501 11509 24535 11543
rect 1501 11305 1535 11339
rect 1685 11305 1719 11339
rect 3893 11305 3927 11339
rect 6561 11305 6595 11339
rect 7481 11305 7515 11339
rect 9137 11305 9171 11339
rect 13277 11305 13311 11339
rect 14381 11305 14415 11339
rect 16497 11305 16531 11339
rect 18889 11305 18923 11339
rect 22661 11305 22695 11339
rect 13553 11237 13587 11271
rect 14105 11237 14139 11271
rect 23029 11237 23063 11271
rect 1961 11169 1995 11203
rect 4169 11169 4203 11203
rect 5089 11169 5123 11203
rect 7021 11169 7055 11203
rect 8309 11169 8343 11203
rect 8401 11169 8435 11203
rect 9597 11169 9631 11203
rect 9689 11169 9723 11203
rect 10977 11169 11011 11203
rect 11805 11169 11839 11203
rect 15025 11169 15059 11203
rect 29745 11169 29779 11203
rect 32045 11169 32079 11203
rect 2605 11101 2639 11135
rect 2881 11101 2915 11135
rect 4813 11101 4847 11135
rect 8217 11101 8251 11135
rect 9505 11101 9539 11135
rect 11529 11101 11563 11135
rect 14749 11101 14783 11135
rect 17141 11101 17175 11135
rect 19533 11101 19567 11135
rect 20913 11101 20947 11135
rect 31769 11101 31803 11135
rect 10701 11033 10735 11067
rect 17417 11033 17451 11067
rect 20269 11033 20303 11067
rect 21189 11033 21223 11067
rect 30021 11033 30055 11067
rect 7849 10965 7883 10999
rect 10333 10965 10367 10999
rect 10793 10965 10827 10999
rect 13829 10965 13863 10999
rect 16773 10965 16807 10999
rect 1777 10761 1811 10795
rect 5825 10761 5859 10795
rect 9873 10761 9907 10795
rect 15577 10761 15611 10795
rect 19257 10761 19291 10795
rect 21925 10761 21959 10795
rect 1685 10693 1719 10727
rect 10701 10693 10735 10727
rect 10793 10693 10827 10727
rect 12357 10693 12391 10727
rect 14841 10693 14875 10727
rect 22017 10693 22051 10727
rect 2421 10625 2455 10659
rect 4721 10625 4755 10659
rect 7021 10625 7055 10659
rect 9505 10625 9539 10659
rect 11621 10625 11655 10659
rect 14749 10625 14783 10659
rect 15945 10625 15979 10659
rect 17509 10625 17543 10659
rect 2053 10557 2087 10591
rect 2145 10557 2179 10591
rect 3433 10557 3467 10591
rect 3709 10557 3743 10591
rect 7481 10557 7515 10591
rect 7757 10557 7791 10591
rect 10057 10557 10091 10591
rect 10885 10557 10919 10591
rect 12081 10557 12115 10591
rect 15025 10557 15059 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 16865 10557 16899 10591
rect 17785 10557 17819 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 1501 10489 1535 10523
rect 10333 10489 10367 10523
rect 14381 10489 14415 10523
rect 21465 10489 21499 10523
rect 5365 10421 5399 10455
rect 6469 10421 6503 10455
rect 6837 10421 6871 10455
rect 13829 10421 13863 10455
rect 1961 10217 1995 10251
rect 3801 10217 3835 10251
rect 9137 10217 9171 10251
rect 10057 10217 10091 10251
rect 16313 10217 16347 10251
rect 18889 10217 18923 10251
rect 21557 10217 21591 10251
rect 6377 10149 6411 10183
rect 6561 10149 6595 10183
rect 1685 10081 1719 10115
rect 2605 10081 2639 10115
rect 2881 10081 2915 10115
rect 4537 10081 4571 10115
rect 6837 10081 6871 10115
rect 9413 10081 9447 10115
rect 10701 10081 10735 10115
rect 13553 10081 13587 10115
rect 14841 10081 14875 10115
rect 19441 10081 19475 10115
rect 2145 10013 2179 10047
rect 4261 10013 4295 10047
rect 5825 10013 5859 10047
rect 11253 10013 11287 10047
rect 14565 10013 14599 10047
rect 17141 10013 17175 10047
rect 7113 9945 7147 9979
rect 10517 9945 10551 9979
rect 11529 9945 11563 9979
rect 17417 9945 17451 9979
rect 19717 9945 19751 9979
rect 21649 9945 21683 9979
rect 1501 9877 1535 9911
rect 5365 9877 5399 9911
rect 8585 9877 8619 9911
rect 10425 9877 10459 9911
rect 13001 9877 13035 9911
rect 14197 9877 14231 9911
rect 16681 9877 16715 9911
rect 16865 9877 16899 9911
rect 21189 9877 21223 9911
rect 1593 9673 1627 9707
rect 6469 9673 6503 9707
rect 16221 9673 16255 9707
rect 1409 9605 1443 9639
rect 3249 9605 3283 9639
rect 5733 9605 5767 9639
rect 5825 9605 5859 9639
rect 10793 9605 10827 9639
rect 11989 9605 12023 9639
rect 13829 9605 13863 9639
rect 13921 9605 13955 9639
rect 14197 9605 14231 9639
rect 17141 9605 17175 9639
rect 19533 9605 19567 9639
rect 28641 9605 28675 9639
rect 2421 9537 2455 9571
rect 3801 9537 3835 9571
rect 6837 9537 6871 9571
rect 10701 9537 10735 9571
rect 19441 9537 19475 9571
rect 20177 9537 20211 9571
rect 27537 9537 27571 9571
rect 1869 9469 1903 9503
rect 2145 9469 2179 9503
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 7113 9469 7147 9503
rect 8125 9469 8159 9503
rect 8401 9469 8435 9503
rect 10885 9469 10919 9503
rect 11713 9469 11747 9503
rect 14473 9469 14507 9503
rect 14749 9469 14783 9503
rect 16865 9469 16899 9503
rect 19717 9469 19751 9503
rect 27997 9469 28031 9503
rect 3617 9401 3651 9435
rect 13461 9401 13495 9435
rect 19073 9401 19107 9435
rect 5365 9333 5399 9367
rect 9873 9333 9907 9367
rect 10333 9333 10367 9367
rect 18613 9333 18647 9367
rect 27813 9333 27847 9367
rect 28457 9333 28491 9367
rect 3525 9129 3559 9163
rect 5273 9129 5307 9163
rect 7205 9129 7239 9163
rect 7849 9129 7883 9163
rect 10149 9129 10183 9163
rect 14289 9129 14323 9163
rect 17785 9129 17819 9163
rect 18153 9129 18187 9163
rect 18797 9129 18831 9163
rect 18981 9129 19015 9163
rect 4537 9061 4571 9095
rect 15393 9061 15427 9095
rect 2513 8993 2547 9027
rect 3433 8993 3467 9027
rect 4629 8993 4663 9027
rect 6193 8993 6227 9027
rect 8401 8993 8435 9027
rect 9413 8993 9447 9027
rect 10793 8993 10827 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 16037 8993 16071 9027
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 5457 8925 5491 8959
rect 5917 8925 5951 8959
rect 7389 8925 7423 8959
rect 8217 8925 8251 8959
rect 11345 8925 11379 8959
rect 11621 8925 11655 8959
rect 10517 8857 10551 8891
rect 13553 8857 13587 8891
rect 14657 8857 14691 8891
rect 16313 8857 16347 8891
rect 1593 8789 1627 8823
rect 3985 8789 4019 8823
rect 8309 8789 8343 8823
rect 9045 8789 9079 8823
rect 10609 8789 10643 8823
rect 12633 8789 12667 8823
rect 7297 8585 7331 8619
rect 10149 8585 10183 8619
rect 12541 8585 12575 8619
rect 14289 8585 14323 8619
rect 15945 8585 15979 8619
rect 5089 8517 5123 8551
rect 5365 8517 5399 8551
rect 11253 8517 11287 8551
rect 16037 8517 16071 8551
rect 1593 8449 1627 8483
rect 2881 8449 2915 8483
rect 3157 8449 3191 8483
rect 4077 8449 4111 8483
rect 4353 8449 4387 8483
rect 4813 8449 4847 8483
rect 6009 8449 6043 8483
rect 7205 8449 7239 8483
rect 7941 8449 7975 8483
rect 8677 8449 8711 8483
rect 10517 8449 10551 8483
rect 11621 8449 11655 8483
rect 13645 8449 13679 8483
rect 14657 8449 14691 8483
rect 1869 8381 1903 8415
rect 8033 8381 8067 8415
rect 8401 8381 8435 8415
rect 9689 8381 9723 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 12633 8381 12667 8415
rect 12817 8381 12851 8415
rect 14749 8381 14783 8415
rect 14933 8381 14967 8415
rect 16221 8381 16255 8415
rect 4629 8313 4663 8347
rect 5825 8313 5859 8347
rect 9873 8313 9907 8347
rect 12173 8313 12207 8347
rect 15577 8313 15611 8347
rect 6377 8245 6411 8279
rect 6745 8245 6779 8279
rect 7757 8245 7791 8279
rect 3433 8041 3467 8075
rect 5181 8041 5215 8075
rect 5365 8041 5399 8075
rect 6377 8041 6411 8075
rect 6561 8041 6595 8075
rect 7573 8041 7607 8075
rect 7757 8041 7791 8075
rect 9597 8041 9631 8075
rect 12449 8041 12483 8075
rect 13001 8041 13035 8075
rect 14197 8041 14231 8075
rect 3525 7973 3559 8007
rect 5733 7973 5767 8007
rect 15209 7973 15243 8007
rect 1593 7905 1627 7939
rect 7113 7905 7147 7939
rect 8769 7905 8803 7939
rect 10241 7905 10275 7939
rect 11253 7905 11287 7939
rect 13645 7905 13679 7939
rect 14841 7905 14875 7939
rect 1869 7837 1903 7871
rect 3065 7837 3099 7871
rect 4169 7837 4203 7871
rect 4813 7837 4847 7871
rect 5457 7837 5491 7871
rect 7849 7837 7883 7871
rect 10057 7837 10091 7871
rect 11529 7837 11563 7871
rect 13461 7837 13495 7871
rect 15025 7837 15059 7871
rect 9965 7769 9999 7803
rect 13369 7769 13403 7803
rect 2881 7701 2915 7735
rect 3985 7701 4019 7735
rect 4629 7701 4663 7735
rect 15853 7701 15887 7735
rect 2881 7497 2915 7531
rect 3617 7497 3651 7531
rect 4629 7497 4663 7531
rect 9137 7497 9171 7531
rect 11897 7497 11931 7531
rect 13461 7497 13495 7531
rect 23949 7497 23983 7531
rect 24317 7429 24351 7463
rect 1593 7361 1627 7395
rect 1869 7361 1903 7395
rect 3065 7361 3099 7395
rect 4169 7361 4203 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 5365 7361 5399 7395
rect 9321 7361 9355 7395
rect 10793 7361 10827 7395
rect 12725 7361 12759 7395
rect 14289 7361 14323 7395
rect 22201 7361 22235 7395
rect 22477 7293 22511 7327
rect 3341 7225 3375 7259
rect 3985 7225 4019 7259
rect 10609 7157 10643 7191
rect 12541 7157 12575 7191
rect 14105 7157 14139 7191
rect 1501 6953 1535 6987
rect 2605 6953 2639 6987
rect 3249 6953 3283 6987
rect 23213 6953 23247 6987
rect 3985 6885 4019 6919
rect 23765 6885 23799 6919
rect 1593 6817 1627 6851
rect 4813 6817 4847 6851
rect 10609 6817 10643 6851
rect 2145 6749 2179 6783
rect 2789 6749 2823 6783
rect 3433 6749 3467 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 22937 6749 22971 6783
rect 1961 6613 1995 6647
rect 4629 6613 4663 6647
rect 23397 6613 23431 6647
rect 3985 6409 4019 6443
rect 22845 6409 22879 6443
rect 1869 6273 1903 6307
rect 3065 6273 3099 6307
rect 3709 6273 3743 6307
rect 4169 6273 4203 6307
rect 22436 6273 22470 6307
rect 1593 6205 1627 6239
rect 22523 6205 22557 6239
rect 3525 6137 3559 6171
rect 2881 6069 2915 6103
rect 3341 5865 3375 5899
rect 3617 5865 3651 5899
rect 18889 5865 18923 5899
rect 21005 5865 21039 5899
rect 2881 5797 2915 5831
rect 19349 5797 19383 5831
rect 21741 5797 21775 5831
rect 1869 5729 1903 5763
rect 15577 5729 15611 5763
rect 17141 5729 17175 5763
rect 27077 5729 27111 5763
rect 1593 5661 1627 5695
rect 3065 5661 3099 5695
rect 15761 5661 15795 5695
rect 20913 5661 20947 5695
rect 17417 5593 17451 5627
rect 24777 5593 24811 5627
rect 24869 5593 24903 5627
rect 25789 5593 25823 5627
rect 27169 5593 27203 5627
rect 28089 5593 28123 5627
rect 16221 5525 16255 5559
rect 21373 5525 21407 5559
rect 2789 5321 2823 5355
rect 2881 5321 2915 5355
rect 3065 5321 3099 5355
rect 22891 5321 22925 5355
rect 28825 5253 28859 5287
rect 1593 5185 1627 5219
rect 1869 5185 1903 5219
rect 15669 5185 15703 5219
rect 17509 5185 17543 5219
rect 22176 5185 22210 5219
rect 22788 5185 22822 5219
rect 15853 5117 15887 5151
rect 17693 5117 17727 5151
rect 28733 5117 28767 5151
rect 29745 5117 29779 5151
rect 3249 5049 3283 5083
rect 16313 4981 16347 5015
rect 18153 4981 18187 5015
rect 22247 4981 22281 5015
rect 2881 4777 2915 4811
rect 19533 4777 19567 4811
rect 20269 4777 20303 4811
rect 24731 4777 24765 4811
rect 3525 4709 3559 4743
rect 1593 4641 1627 4675
rect 1869 4641 1903 4675
rect 25881 4641 25915 4675
rect 3065 4573 3099 4607
rect 3341 4573 3375 4607
rect 19441 4573 19475 4607
rect 24628 4573 24662 4607
rect 25973 4505 26007 4539
rect 26893 4505 26927 4539
rect 19901 4437 19935 4471
rect 1409 4233 1443 4267
rect 1869 4097 1903 4131
rect 2513 4097 2547 4131
rect 2973 4097 3007 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 15209 4097 15243 4131
rect 4077 3961 4111 3995
rect 3617 3893 3651 3927
rect 15025 3893 15059 3927
rect 3985 3689 4019 3723
rect 12081 3689 12115 3723
rect 2973 3621 3007 3655
rect 1593 3553 1627 3587
rect 4629 3553 4663 3587
rect 1869 3485 1903 3519
rect 3157 3485 3191 3519
rect 3433 3485 3467 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 11529 3485 11563 3519
rect 35725 3485 35759 3519
rect 37841 3485 37875 3519
rect 36921 3417 36955 3451
rect 39037 3417 39071 3451
rect 11621 3349 11655 3383
rect 3985 3145 4019 3179
rect 14013 3145 14047 3179
rect 25513 3145 25547 3179
rect 28181 3145 28215 3179
rect 33517 3145 33551 3179
rect 10793 3077 10827 3111
rect 12633 3077 12667 3111
rect 13921 3077 13955 3111
rect 15577 3077 15611 3111
rect 1593 3009 1627 3043
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 4169 3009 4203 3043
rect 4629 3009 4663 3043
rect 5273 3009 5307 3043
rect 6561 3009 6595 3043
rect 8769 3009 8803 3043
rect 17049 3009 17083 3043
rect 18337 3009 18371 3043
rect 20545 3009 20579 3043
rect 25697 3009 25731 3043
rect 28365 3009 28399 3043
rect 31033 3009 31067 3043
rect 33701 3009 33735 3043
rect 35265 3009 35299 3043
rect 37473 3009 37507 3043
rect 1869 2941 1903 2975
rect 7205 2941 7239 2975
rect 9045 2941 9079 2975
rect 10517 2941 10551 2975
rect 36461 2941 36495 2975
rect 38577 2941 38611 2975
rect 15761 2873 15795 2907
rect 30849 2873 30883 2907
rect 12725 2805 12759 2839
rect 16865 2805 16899 2839
rect 18153 2805 18187 2839
rect 20361 2805 20395 2839
rect 2881 2601 2915 2635
rect 26249 2601 26283 2635
rect 28917 2601 28951 2635
rect 31585 2601 31619 2635
rect 34253 2601 34287 2635
rect 3525 2533 3559 2567
rect 1593 2465 1627 2499
rect 3801 2465 3835 2499
rect 4629 2465 4663 2499
rect 7297 2465 7331 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 15301 2465 15335 2499
rect 17969 2465 18003 2499
rect 20545 2465 20579 2499
rect 23121 2465 23155 2499
rect 36369 2465 36403 2499
rect 3065 2397 3099 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 9597 2397 9631 2431
rect 12357 2397 12391 2431
rect 15025 2397 15059 2431
rect 17509 2397 17543 2431
rect 20085 2397 20119 2431
rect 22661 2397 22695 2431
rect 25605 2397 25639 2431
rect 28273 2397 28307 2431
rect 30941 2397 30975 2431
rect 33609 2397 33643 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
rect 3341 2329 3375 2363
rect 1823 2261 1857 2295
rect 25329 2261 25363 2295
rect 27905 2261 27939 2295
rect 30665 2261 30699 2295
rect 33333 2261 33367 2295
<< metal1 >>
rect 9674 25576 9680 25628
rect 9732 25616 9738 25628
rect 21818 25616 21824 25628
rect 9732 25588 21824 25616
rect 9732 25576 9738 25588
rect 21818 25576 21824 25588
rect 21876 25576 21882 25628
rect 4798 25508 4804 25560
rect 4856 25548 4862 25560
rect 21174 25548 21180 25560
rect 4856 25520 21180 25548
rect 4856 25508 4862 25520
rect 21174 25508 21180 25520
rect 21232 25508 21238 25560
rect 10042 25440 10048 25492
rect 10100 25480 10106 25492
rect 28442 25480 28448 25492
rect 10100 25452 28448 25480
rect 10100 25440 10106 25452
rect 28442 25440 28448 25452
rect 28500 25440 28506 25492
rect 12066 25372 12072 25424
rect 12124 25412 12130 25424
rect 33962 25412 33968 25424
rect 12124 25384 33968 25412
rect 12124 25372 12130 25384
rect 33962 25372 33968 25384
rect 34020 25372 34026 25424
rect 12342 25304 12348 25356
rect 12400 25344 12406 25356
rect 26418 25344 26424 25356
rect 12400 25316 26424 25344
rect 12400 25304 12406 25316
rect 26418 25304 26424 25316
rect 26476 25304 26482 25356
rect 17770 25236 17776 25288
rect 17828 25276 17834 25288
rect 34330 25276 34336 25288
rect 17828 25248 34336 25276
rect 17828 25236 17834 25248
rect 34330 25236 34336 25248
rect 34388 25236 34394 25288
rect 15378 25168 15384 25220
rect 15436 25208 15442 25220
rect 33594 25208 33600 25220
rect 15436 25180 33600 25208
rect 15436 25168 15442 25180
rect 33594 25168 33600 25180
rect 33652 25168 33658 25220
rect 10594 25100 10600 25152
rect 10652 25140 10658 25152
rect 30374 25140 30380 25152
rect 10652 25112 30380 25140
rect 10652 25100 10658 25112
rect 30374 25100 30380 25112
rect 30432 25100 30438 25152
rect 4062 25032 4068 25084
rect 4120 25072 4126 25084
rect 8478 25072 8484 25084
rect 4120 25044 8484 25072
rect 4120 25032 4126 25044
rect 8478 25032 8484 25044
rect 8536 25032 8542 25084
rect 12710 25032 12716 25084
rect 12768 25072 12774 25084
rect 33410 25072 33416 25084
rect 12768 25044 33416 25072
rect 12768 25032 12774 25044
rect 33410 25032 33416 25044
rect 33468 25032 33474 25084
rect 15010 24964 15016 25016
rect 15068 25004 15074 25016
rect 30006 25004 30012 25016
rect 15068 24976 30012 25004
rect 15068 24964 15074 24976
rect 30006 24964 30012 24976
rect 30064 24964 30070 25016
rect 30558 24964 30564 25016
rect 30616 25004 30622 25016
rect 32858 25004 32864 25016
rect 30616 24976 32864 25004
rect 30616 24964 30622 24976
rect 32858 24964 32864 24976
rect 32916 24964 32922 25016
rect 14826 24896 14832 24948
rect 14884 24936 14890 24948
rect 39298 24936 39304 24948
rect 14884 24908 39304 24936
rect 14884 24896 14890 24908
rect 39298 24896 39304 24908
rect 39356 24896 39362 24948
rect 10778 24828 10784 24880
rect 10836 24868 10842 24880
rect 36538 24868 36544 24880
rect 10836 24840 36544 24868
rect 10836 24828 10842 24840
rect 36538 24828 36544 24840
rect 36596 24828 36602 24880
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 8294 24800 8300 24812
rect 4120 24772 8300 24800
rect 4120 24760 4126 24772
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 11698 24760 11704 24812
rect 11756 24800 11762 24812
rect 21910 24800 21916 24812
rect 11756 24772 21916 24800
rect 11756 24760 11762 24772
rect 21910 24760 21916 24772
rect 21968 24760 21974 24812
rect 22646 24760 22652 24812
rect 22704 24800 22710 24812
rect 28534 24800 28540 24812
rect 22704 24772 28540 24800
rect 22704 24760 22710 24772
rect 28534 24760 28540 24772
rect 28592 24760 28598 24812
rect 28626 24760 28632 24812
rect 28684 24800 28690 24812
rect 32306 24800 32312 24812
rect 28684 24772 32312 24800
rect 28684 24760 28690 24772
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 4246 24692 4252 24744
rect 4304 24732 4310 24744
rect 4304 24704 17080 24732
rect 4304 24692 4310 24704
rect 6454 24624 6460 24676
rect 6512 24664 6518 24676
rect 13630 24664 13636 24676
rect 6512 24636 13636 24664
rect 6512 24624 6518 24636
rect 13630 24624 13636 24636
rect 13688 24624 13694 24676
rect 17052 24596 17080 24704
rect 25038 24692 25044 24744
rect 25096 24732 25102 24744
rect 30558 24732 30564 24744
rect 25096 24704 30564 24732
rect 25096 24692 25102 24704
rect 30558 24692 30564 24704
rect 30616 24692 30622 24744
rect 35526 24732 35532 24744
rect 31726 24704 35532 24732
rect 17126 24624 17132 24676
rect 17184 24664 17190 24676
rect 18598 24664 18604 24676
rect 17184 24636 18604 24664
rect 17184 24624 17190 24636
rect 18598 24624 18604 24636
rect 18656 24664 18662 24676
rect 25958 24664 25964 24676
rect 18656 24636 25964 24664
rect 18656 24624 18662 24636
rect 25958 24624 25964 24636
rect 26016 24624 26022 24676
rect 27522 24624 27528 24676
rect 27580 24664 27586 24676
rect 31294 24664 31300 24676
rect 27580 24636 31300 24664
rect 27580 24624 27586 24636
rect 31294 24624 31300 24636
rect 31352 24624 31358 24676
rect 24118 24596 24124 24608
rect 17052 24568 24124 24596
rect 24118 24556 24124 24568
rect 24176 24556 24182 24608
rect 25222 24556 25228 24608
rect 25280 24596 25286 24608
rect 28994 24596 29000 24608
rect 25280 24568 29000 24596
rect 25280 24556 25286 24568
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 29086 24556 29092 24608
rect 29144 24596 29150 24608
rect 31726 24596 31754 24704
rect 35526 24692 35532 24704
rect 35584 24692 35590 24744
rect 29144 24568 31754 24596
rect 29144 24556 29150 24568
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 5258 24392 5264 24404
rect 2832 24364 5264 24392
rect 2832 24352 2838 24364
rect 5258 24352 5264 24364
rect 5316 24352 5322 24404
rect 9125 24395 9183 24401
rect 9125 24361 9137 24395
rect 9171 24392 9183 24395
rect 16482 24392 16488 24404
rect 9171 24364 16488 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 18966 24392 18972 24404
rect 16776 24364 18972 24392
rect 566 24284 572 24336
rect 624 24324 630 24336
rect 624 24296 3924 24324
rect 624 24284 630 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 1026 24148 1032 24200
rect 1084 24188 1090 24200
rect 3896 24197 3924 24296
rect 9306 24284 9312 24336
rect 9364 24284 9370 24336
rect 14734 24324 14740 24336
rect 9692 24296 14740 24324
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 7374 24256 7380 24268
rect 5859 24228 7380 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 7374 24216 7380 24228
rect 7432 24216 7438 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9324 24256 9352 24284
rect 8251 24228 9352 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 2041 24191 2099 24197
rect 2041 24188 2053 24191
rect 1084 24160 2053 24188
rect 1084 24148 1090 24160
rect 2041 24157 2053 24160
rect 2087 24157 2099 24191
rect 2041 24151 2099 24157
rect 3881 24191 3939 24197
rect 3881 24157 3893 24191
rect 3927 24188 3939 24191
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 3927 24160 4169 24188
rect 3927 24157 3939 24160
rect 3881 24151 3939 24157
rect 4157 24157 4169 24160
rect 4203 24188 4215 24191
rect 4246 24188 4252 24200
rect 4203 24160 4252 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4246 24148 4252 24160
rect 4304 24148 4310 24200
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 6457 24191 6515 24197
rect 6457 24157 6469 24191
rect 6503 24188 6515 24191
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 6503 24160 6745 24188
rect 6503 24157 6515 24160
rect 6457 24151 6515 24157
rect 6733 24157 6745 24160
rect 6779 24188 6791 24191
rect 6822 24188 6828 24200
rect 6779 24160 6828 24188
rect 6779 24157 6791 24160
rect 6733 24151 6791 24157
rect 658 24080 664 24132
rect 716 24120 722 24132
rect 4632 24120 4660 24151
rect 6822 24148 6828 24160
rect 6880 24148 6886 24200
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24188 7343 24191
rect 8570 24188 8576 24200
rect 7331 24160 8576 24188
rect 7331 24157 7343 24160
rect 7285 24151 7343 24157
rect 8570 24148 8576 24160
rect 8628 24148 8634 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9692 24188 9720 24296
rect 14734 24284 14740 24296
rect 14792 24284 14798 24336
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 13541 24259 13599 24265
rect 11011 24228 12020 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 9355 24160 9720 24188
rect 9953 24191 10011 24197
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10042 24188 10048 24200
rect 9999 24160 10048 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 10042 24148 10048 24160
rect 10100 24148 10106 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 716 24092 4660 24120
rect 716 24080 722 24092
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 1673 24055 1731 24061
rect 1673 24052 1685 24055
rect 1627 24024 1685 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 1673 24021 1685 24024
rect 1719 24052 1731 24055
rect 3694 24052 3700 24064
rect 1719 24024 3700 24052
rect 1719 24021 1731 24024
rect 1673 24015 1731 24021
rect 3694 24012 3700 24024
rect 3752 24012 3758 24064
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 6270 24052 6276 24064
rect 4019 24024 6276 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 6270 24012 6276 24024
rect 6328 24012 6334 24064
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 9674 24052 9680 24064
rect 6595 24024 9680 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 9674 24012 9680 24024
rect 9732 24012 9738 24064
rect 11698 24012 11704 24064
rect 11756 24012 11762 24064
rect 11900 24052 11928 24151
rect 11992 24120 12020 24228
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 14366 24256 14372 24268
rect 13587 24228 14372 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 14366 24216 14372 24228
rect 14424 24216 14430 24268
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 16776 24256 16804 24364
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 19058 24352 19064 24404
rect 19116 24392 19122 24404
rect 19116 24364 26648 24392
rect 19116 24352 19122 24364
rect 23845 24327 23903 24333
rect 23845 24293 23857 24327
rect 23891 24324 23903 24327
rect 23891 24296 26464 24324
rect 23891 24293 23903 24296
rect 23845 24287 23903 24293
rect 16163 24228 16804 24256
rect 16853 24259 16911 24265
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 18690 24256 18696 24268
rect 16899 24228 18696 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 22094 24216 22100 24268
rect 22152 24256 22158 24268
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 22152 24228 22477 24256
rect 22152 24216 22158 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 25038 24216 25044 24268
rect 25096 24216 25102 24268
rect 25222 24216 25228 24268
rect 25280 24216 25286 24268
rect 26329 24259 26387 24265
rect 26329 24225 26341 24259
rect 26375 24225 26387 24259
rect 26329 24219 26387 24225
rect 12434 24148 12440 24200
rect 12492 24148 12498 24200
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24188 14519 24191
rect 14550 24188 14556 24200
rect 14507 24160 14556 24188
rect 14507 24157 14519 24160
rect 14461 24151 14519 24157
rect 14550 24148 14556 24160
rect 14608 24148 14614 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 16574 24188 16580 24200
rect 15151 24160 16580 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 18414 24148 18420 24200
rect 18472 24188 18478 24200
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 18472 24160 19625 24188
rect 18472 24148 18478 24160
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19886 24148 19892 24200
rect 19944 24188 19950 24200
rect 20073 24191 20131 24197
rect 20073 24188 20085 24191
rect 19944 24160 20085 24188
rect 19944 24148 19950 24160
rect 20073 24157 20085 24160
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21968 24160 22017 24188
rect 21968 24148 21974 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 23566 24148 23572 24200
rect 23624 24188 23630 24200
rect 24029 24191 24087 24197
rect 24029 24188 24041 24191
rect 23624 24160 24041 24188
rect 23624 24148 23630 24160
rect 24029 24157 24041 24160
rect 24075 24188 24087 24191
rect 24762 24188 24768 24200
rect 24075 24160 24768 24188
rect 24075 24157 24087 24160
rect 24029 24151 24087 24157
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 13814 24120 13820 24132
rect 11992 24092 13820 24120
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 15286 24120 15292 24132
rect 13924 24092 15292 24120
rect 13924 24052 13952 24092
rect 15286 24080 15292 24092
rect 15344 24080 15350 24132
rect 17126 24080 17132 24132
rect 17184 24080 17190 24132
rect 18506 24120 18512 24132
rect 18354 24092 18512 24120
rect 18506 24080 18512 24092
rect 18564 24120 18570 24132
rect 19061 24123 19119 24129
rect 19061 24120 19073 24123
rect 18564 24092 19073 24120
rect 18564 24080 18570 24092
rect 19061 24089 19073 24092
rect 19107 24120 19119 24123
rect 19518 24120 19524 24132
rect 19107 24092 19524 24120
rect 19107 24089 19119 24092
rect 19061 24083 19119 24089
rect 19518 24080 19524 24092
rect 19576 24080 19582 24132
rect 23934 24080 23940 24132
rect 23992 24120 23998 24132
rect 23992 24092 25820 24120
rect 23992 24080 23998 24092
rect 11900 24024 13952 24052
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 17034 24012 17040 24064
rect 17092 24052 17098 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 17092 24024 18613 24052
rect 17092 24012 17098 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 18601 24015 18659 24021
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 20162 24052 20168 24064
rect 19475 24024 20168 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 24578 24012 24584 24064
rect 24636 24012 24642 24064
rect 24946 24012 24952 24064
rect 25004 24012 25010 24064
rect 25792 24061 25820 24092
rect 25958 24080 25964 24132
rect 26016 24120 26022 24132
rect 26344 24120 26372 24219
rect 26436 24188 26464 24296
rect 26620 24256 26648 24364
rect 26970 24352 26976 24404
rect 27028 24392 27034 24404
rect 29454 24392 29460 24404
rect 27028 24364 29460 24392
rect 27028 24352 27034 24364
rect 29454 24352 29460 24364
rect 29512 24352 29518 24404
rect 29546 24352 29552 24404
rect 29604 24392 29610 24404
rect 31018 24392 31024 24404
rect 29604 24364 31024 24392
rect 29604 24352 29610 24364
rect 31018 24352 31024 24364
rect 31076 24352 31082 24404
rect 31294 24352 31300 24404
rect 31352 24392 31358 24404
rect 34790 24392 34796 24404
rect 31352 24364 34796 24392
rect 31352 24352 31358 24364
rect 34790 24352 34796 24364
rect 34848 24352 34854 24404
rect 37921 24395 37979 24401
rect 37921 24392 37933 24395
rect 35360 24364 37933 24392
rect 27338 24284 27344 24336
rect 27396 24324 27402 24336
rect 30742 24324 30748 24336
rect 27396 24296 30748 24324
rect 27396 24284 27402 24296
rect 30742 24284 30748 24296
rect 30800 24284 30806 24336
rect 33778 24284 33784 24336
rect 33836 24324 33842 24336
rect 33836 24296 34836 24324
rect 33836 24284 33842 24296
rect 27709 24259 27767 24265
rect 27709 24256 27721 24259
rect 26620 24228 27721 24256
rect 27709 24225 27721 24228
rect 27755 24225 27767 24259
rect 27709 24219 27767 24225
rect 29733 24259 29791 24265
rect 29733 24225 29745 24259
rect 29779 24256 29791 24259
rect 31665 24259 31723 24265
rect 31665 24256 31677 24259
rect 29779 24228 31677 24256
rect 29779 24225 29791 24228
rect 29733 24219 29791 24225
rect 31665 24225 31677 24228
rect 31711 24225 31723 24259
rect 34808 24256 34836 24296
rect 35360 24256 35388 24364
rect 37921 24361 37933 24364
rect 37967 24361 37979 24395
rect 37921 24355 37979 24361
rect 41506 24352 41512 24404
rect 41564 24392 41570 24404
rect 42429 24395 42487 24401
rect 42429 24392 42441 24395
rect 41564 24364 42441 24392
rect 41564 24352 41570 24364
rect 42429 24361 42441 24364
rect 42475 24392 42487 24395
rect 42610 24392 42616 24404
rect 42475 24364 42616 24392
rect 42475 24361 42487 24364
rect 42429 24355 42487 24361
rect 42610 24352 42616 24364
rect 42668 24352 42674 24404
rect 44726 24352 44732 24404
rect 44784 24352 44790 24404
rect 46845 24395 46903 24401
rect 46845 24392 46857 24395
rect 44836 24364 46857 24392
rect 35618 24284 35624 24336
rect 35676 24324 35682 24336
rect 36909 24327 36967 24333
rect 36909 24324 36921 24327
rect 35676 24296 36921 24324
rect 35676 24284 35682 24296
rect 36909 24293 36921 24296
rect 36955 24293 36967 24327
rect 36909 24287 36967 24293
rect 37090 24284 37096 24336
rect 37148 24324 37154 24336
rect 39393 24327 39451 24333
rect 39393 24324 39405 24327
rect 37148 24296 39405 24324
rect 37148 24284 37154 24296
rect 39393 24293 39405 24296
rect 39439 24293 39451 24327
rect 39393 24287 39451 24293
rect 43438 24284 43444 24336
rect 43496 24324 43502 24336
rect 44836 24324 44864 24364
rect 46845 24361 46857 24364
rect 46891 24361 46903 24395
rect 46845 24355 46903 24361
rect 43496 24296 44864 24324
rect 43496 24284 43502 24296
rect 44910 24284 44916 24336
rect 44968 24324 44974 24336
rect 47949 24327 48007 24333
rect 47949 24324 47961 24327
rect 44968 24296 47961 24324
rect 44968 24284 44974 24296
rect 47949 24293 47961 24296
rect 47995 24293 48007 24327
rect 47949 24287 48007 24293
rect 31665 24219 31723 24225
rect 32324 24228 34468 24256
rect 27617 24191 27675 24197
rect 27617 24188 27629 24191
rect 26436 24160 27629 24188
rect 27617 24157 27629 24160
rect 27663 24157 27675 24191
rect 27617 24151 27675 24157
rect 27982 24148 27988 24200
rect 28040 24188 28046 24200
rect 28442 24188 28448 24200
rect 28040 24160 28448 24188
rect 28040 24148 28046 24160
rect 28442 24148 28448 24160
rect 28500 24188 28506 24200
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 28500 24160 28549 24188
rect 28500 24148 28506 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 30009 24191 30067 24197
rect 30009 24188 30021 24191
rect 28537 24151 28595 24157
rect 28644 24160 30021 24188
rect 26016 24092 26372 24120
rect 26016 24080 26022 24092
rect 26418 24080 26424 24132
rect 26476 24120 26482 24132
rect 28644 24120 28672 24160
rect 30009 24157 30021 24160
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 31018 24148 31024 24200
rect 31076 24188 31082 24200
rect 31386 24188 31392 24200
rect 31076 24160 31392 24188
rect 31076 24148 31082 24160
rect 31386 24148 31392 24160
rect 31444 24148 31450 24200
rect 32324 24197 32352 24228
rect 32309 24191 32367 24197
rect 32309 24188 32321 24191
rect 31726 24160 32321 24188
rect 26476 24092 28672 24120
rect 26476 24080 26482 24092
rect 29914 24080 29920 24132
rect 29972 24120 29978 24132
rect 31726 24120 31754 24160
rect 32309 24157 32321 24160
rect 32355 24157 32367 24191
rect 32309 24151 32367 24157
rect 33318 24148 33324 24200
rect 33376 24188 33382 24200
rect 33413 24191 33471 24197
rect 33413 24188 33425 24191
rect 33376 24160 33425 24188
rect 33376 24148 33382 24160
rect 33413 24157 33425 24160
rect 33459 24157 33471 24191
rect 33413 24151 33471 24157
rect 29972 24092 31754 24120
rect 29972 24080 29978 24092
rect 32030 24080 32036 24132
rect 32088 24120 32094 24132
rect 34333 24123 34391 24129
rect 34333 24120 34345 24123
rect 32088 24092 34345 24120
rect 32088 24080 32094 24092
rect 34333 24089 34345 24092
rect 34379 24089 34391 24123
rect 34440 24120 34468 24228
rect 34808 24228 35388 24256
rect 34808 24188 34836 24228
rect 35526 24216 35532 24268
rect 35584 24256 35590 24268
rect 47670 24256 47676 24268
rect 35584 24228 47676 24256
rect 35584 24216 35590 24228
rect 47670 24216 47676 24228
rect 47728 24216 47734 24268
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34808 24160 34897 24188
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 35066 24148 35072 24200
rect 35124 24188 35130 24200
rect 35989 24191 36047 24197
rect 35989 24188 36001 24191
rect 35124 24160 36001 24188
rect 35124 24148 35130 24160
rect 35989 24157 36001 24160
rect 36035 24157 36047 24191
rect 35989 24151 36047 24157
rect 35618 24120 35624 24132
rect 34440 24092 35624 24120
rect 34333 24083 34391 24089
rect 35618 24080 35624 24092
rect 35676 24080 35682 24132
rect 36004 24120 36032 24151
rect 36354 24148 36360 24200
rect 36412 24188 36418 24200
rect 37645 24191 37703 24197
rect 37645 24188 37657 24191
rect 36412 24160 37657 24188
rect 36412 24148 36418 24160
rect 37645 24157 37657 24160
rect 37691 24188 37703 24191
rect 37691 24160 38240 24188
rect 37691 24157 37703 24160
rect 37645 24151 37703 24157
rect 38105 24123 38163 24129
rect 38105 24120 38117 24123
rect 36004 24092 38117 24120
rect 38105 24089 38117 24092
rect 38151 24089 38163 24123
rect 38212 24120 38240 24160
rect 38470 24148 38476 24200
rect 38528 24148 38534 24200
rect 38930 24148 38936 24200
rect 38988 24188 38994 24200
rect 39942 24188 39948 24200
rect 38988 24160 39948 24188
rect 38988 24148 38994 24160
rect 39942 24148 39948 24160
rect 40000 24188 40006 24200
rect 40037 24191 40095 24197
rect 40037 24188 40049 24191
rect 40000 24160 40049 24188
rect 40000 24148 40006 24160
rect 40037 24157 40049 24160
rect 40083 24157 40095 24191
rect 40037 24151 40095 24157
rect 40218 24148 40224 24200
rect 40276 24188 40282 24200
rect 41141 24191 41199 24197
rect 41141 24188 41153 24191
rect 40276 24160 41153 24188
rect 40276 24148 40282 24160
rect 41141 24157 41153 24160
rect 41187 24188 41199 24191
rect 42061 24191 42119 24197
rect 42061 24188 42073 24191
rect 41187 24160 42073 24188
rect 41187 24157 41199 24160
rect 41141 24151 41199 24157
rect 42061 24157 42073 24160
rect 42107 24157 42119 24191
rect 42061 24151 42119 24157
rect 44174 24148 44180 24200
rect 44232 24188 44238 24200
rect 44361 24191 44419 24197
rect 44361 24188 44373 24191
rect 44232 24160 44373 24188
rect 44232 24148 44238 24160
rect 44361 24157 44373 24160
rect 44407 24157 44419 24191
rect 44361 24151 44419 24157
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44784 24160 45201 24188
rect 44784 24148 44790 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45922 24188 45928 24200
rect 45612 24160 45928 24188
rect 45612 24148 45618 24160
rect 45922 24148 45928 24160
rect 45980 24148 45986 24200
rect 46014 24148 46020 24200
rect 46072 24188 46078 24200
rect 46661 24191 46719 24197
rect 46661 24188 46673 24191
rect 46072 24160 46673 24188
rect 46072 24148 46078 24160
rect 46661 24157 46673 24160
rect 46707 24188 46719 24191
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 46707 24160 47225 24188
rect 46707 24157 46719 24160
rect 46661 24151 46719 24157
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 47765 24191 47823 24197
rect 47765 24188 47777 24191
rect 47360 24160 47777 24188
rect 47360 24148 47366 24160
rect 47765 24157 47777 24160
rect 47811 24157 47823 24191
rect 47765 24151 47823 24157
rect 48590 24148 48596 24200
rect 48648 24148 48654 24200
rect 39577 24123 39635 24129
rect 39577 24120 39589 24123
rect 38212 24092 39589 24120
rect 38105 24083 38163 24089
rect 39577 24089 39589 24092
rect 39623 24089 39635 24123
rect 39577 24083 39635 24089
rect 43346 24080 43352 24132
rect 43404 24120 43410 24132
rect 43404 24092 45554 24120
rect 43404 24080 43410 24092
rect 25777 24055 25835 24061
rect 25777 24021 25789 24055
rect 25823 24021 25835 24055
rect 25777 24015 25835 24021
rect 25866 24012 25872 24064
rect 25924 24052 25930 24064
rect 26145 24055 26203 24061
rect 26145 24052 26157 24055
rect 25924 24024 26157 24052
rect 25924 24012 25930 24024
rect 26145 24021 26157 24024
rect 26191 24021 26203 24055
rect 26145 24015 26203 24021
rect 26234 24012 26240 24064
rect 26292 24012 26298 24064
rect 26326 24012 26332 24064
rect 26384 24052 26390 24064
rect 27157 24055 27215 24061
rect 27157 24052 27169 24055
rect 26384 24024 27169 24052
rect 26384 24012 26390 24024
rect 27157 24021 27169 24024
rect 27203 24021 27215 24055
rect 27157 24015 27215 24021
rect 27338 24012 27344 24064
rect 27396 24052 27402 24064
rect 27525 24055 27583 24061
rect 27525 24052 27537 24055
rect 27396 24024 27537 24052
rect 27396 24012 27402 24024
rect 27525 24021 27537 24024
rect 27571 24021 27583 24055
rect 27525 24015 27583 24021
rect 28261 24055 28319 24061
rect 28261 24021 28273 24055
rect 28307 24052 28319 24055
rect 28350 24052 28356 24064
rect 28307 24024 28356 24052
rect 28307 24021 28319 24024
rect 28261 24015 28319 24021
rect 28350 24012 28356 24024
rect 28408 24012 28414 24064
rect 29178 24012 29184 24064
rect 29236 24012 29242 24064
rect 30650 24012 30656 24064
rect 30708 24052 30714 24064
rect 32953 24055 33011 24061
rect 32953 24052 32965 24055
rect 30708 24024 32965 24052
rect 30708 24012 30714 24024
rect 32953 24021 32965 24024
rect 32999 24021 33011 24055
rect 32953 24015 33011 24021
rect 33502 24012 33508 24064
rect 33560 24052 33566 24064
rect 34057 24055 34115 24061
rect 34057 24052 34069 24055
rect 33560 24024 34069 24052
rect 33560 24012 33566 24024
rect 34057 24021 34069 24024
rect 34103 24021 34115 24055
rect 34057 24015 34115 24021
rect 34146 24012 34152 24064
rect 34204 24052 34210 24064
rect 35529 24055 35587 24061
rect 35529 24052 35541 24055
rect 34204 24024 35541 24052
rect 34204 24012 34210 24024
rect 35529 24021 35541 24024
rect 35575 24021 35587 24055
rect 35529 24015 35587 24021
rect 35986 24012 35992 24064
rect 36044 24052 36050 24064
rect 36633 24055 36691 24061
rect 36633 24052 36645 24055
rect 36044 24024 36645 24052
rect 36044 24012 36050 24024
rect 36633 24021 36645 24024
rect 36679 24021 36691 24055
rect 36633 24015 36691 24021
rect 37366 24012 37372 24064
rect 37424 24052 37430 24064
rect 37461 24055 37519 24061
rect 37461 24052 37473 24055
rect 37424 24024 37473 24052
rect 37424 24012 37430 24024
rect 37461 24021 37473 24024
rect 37507 24021 37519 24055
rect 37461 24015 37519 24021
rect 38470 24012 38476 24064
rect 38528 24052 38534 24064
rect 39117 24055 39175 24061
rect 39117 24052 39129 24055
rect 38528 24024 39129 24052
rect 38528 24012 38534 24024
rect 39117 24021 39129 24024
rect 39163 24021 39175 24055
rect 39117 24015 39175 24021
rect 40678 24012 40684 24064
rect 40736 24012 40742 24064
rect 41414 24012 41420 24064
rect 41472 24052 41478 24064
rect 41785 24055 41843 24061
rect 41785 24052 41797 24055
rect 41472 24024 41797 24052
rect 41472 24012 41478 24024
rect 41785 24021 41797 24024
rect 41831 24021 41843 24055
rect 41785 24015 41843 24021
rect 42794 24012 42800 24064
rect 42852 24052 42858 24064
rect 44177 24055 44235 24061
rect 44177 24052 44189 24055
rect 42852 24024 44189 24052
rect 42852 24012 42858 24024
rect 44177 24021 44189 24024
rect 44223 24021 44235 24055
rect 44177 24015 44235 24021
rect 45370 24012 45376 24064
rect 45428 24012 45434 24064
rect 45526 24052 45554 24092
rect 46109 24055 46167 24061
rect 46109 24052 46121 24055
rect 45526 24024 46121 24052
rect 46109 24021 46121 24024
rect 46155 24021 46167 24055
rect 46109 24015 46167 24021
rect 48682 24012 48688 24064
rect 48740 24052 48746 24064
rect 49237 24055 49295 24061
rect 49237 24052 49249 24055
rect 48740 24024 49249 24052
rect 48740 24012 48746 24024
rect 49237 24021 49249 24024
rect 49283 24021 49295 24055
rect 49237 24015 49295 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 1765 23851 1823 23857
rect 1765 23817 1777 23851
rect 1811 23848 1823 23851
rect 1811 23820 5672 23848
rect 1811 23817 1823 23820
rect 1765 23811 1823 23817
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4154 23780 4160 23792
rect 4019 23752 4160 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 5644 23780 5672 23820
rect 6454 23808 6460 23860
rect 6512 23808 6518 23860
rect 9766 23848 9772 23860
rect 6564 23820 9772 23848
rect 6564 23780 6592 23820
rect 9766 23808 9772 23820
rect 9824 23808 9830 23860
rect 12345 23851 12403 23857
rect 12345 23817 12357 23851
rect 12391 23848 12403 23851
rect 23934 23848 23940 23860
rect 12391 23820 23940 23848
rect 12391 23817 12403 23820
rect 12345 23811 12403 23817
rect 23934 23808 23940 23820
rect 23992 23808 23998 23860
rect 24213 23851 24271 23857
rect 24213 23817 24225 23851
rect 24259 23848 24271 23851
rect 24946 23848 24952 23860
rect 24259 23820 24952 23848
rect 24259 23817 24271 23820
rect 24213 23811 24271 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 28442 23808 28448 23860
rect 28500 23848 28506 23860
rect 28500 23820 29132 23848
rect 28500 23808 28506 23820
rect 5644 23752 6592 23780
rect 7193 23783 7251 23789
rect 7193 23749 7205 23783
rect 7239 23780 7251 23783
rect 7374 23780 7380 23792
rect 7239 23752 7380 23780
rect 7239 23749 7251 23752
rect 7193 23743 7251 23749
rect 7374 23740 7380 23752
rect 7432 23740 7438 23792
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9950 23780 9956 23792
rect 9171 23752 9956 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 12526 23780 12532 23792
rect 11011 23752 12532 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 15746 23780 15752 23792
rect 14323 23752 15752 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 17126 23780 17132 23792
rect 16040 23752 17132 23780
rect 750 23672 756 23724
rect 808 23712 814 23724
rect 2133 23715 2191 23721
rect 2133 23712 2145 23715
rect 808 23684 2145 23712
rect 808 23672 814 23684
rect 2133 23681 2145 23684
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 2976 23644 3004 23675
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 7101 23715 7159 23721
rect 7101 23712 7113 23715
rect 6604 23684 7113 23712
rect 6604 23672 6610 23684
rect 7101 23681 7113 23684
rect 7147 23681 7159 23715
rect 7101 23675 7159 23681
rect 7650 23672 7656 23724
rect 7708 23712 7714 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7708 23684 7941 23712
rect 7708 23672 7714 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 9858 23672 9864 23724
rect 9916 23672 9922 23724
rect 11790 23672 11796 23724
rect 11848 23712 11854 23724
rect 12253 23715 12311 23721
rect 12253 23712 12265 23715
rect 11848 23684 12265 23712
rect 11848 23672 11854 23684
rect 12253 23681 12265 23684
rect 12299 23681 12311 23715
rect 12253 23675 12311 23681
rect 13262 23672 13268 23724
rect 13320 23672 13326 23724
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23712 15163 23715
rect 16040 23712 16068 23752
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 17865 23783 17923 23789
rect 17865 23749 17877 23783
rect 17911 23780 17923 23783
rect 19242 23780 19248 23792
rect 17911 23752 19248 23780
rect 17911 23749 17923 23752
rect 17865 23743 17923 23749
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 19518 23740 19524 23792
rect 19576 23740 19582 23792
rect 21174 23740 21180 23792
rect 21232 23740 21238 23792
rect 23658 23780 23664 23792
rect 23506 23752 23664 23780
rect 23658 23740 23664 23752
rect 23716 23740 23722 23792
rect 26418 23780 26424 23792
rect 26358 23752 26424 23780
rect 26418 23740 26424 23752
rect 26476 23780 26482 23792
rect 29104 23780 29132 23820
rect 29178 23808 29184 23860
rect 29236 23848 29242 23860
rect 29236 23820 34376 23848
rect 29236 23808 29242 23820
rect 26476 23752 27922 23780
rect 29104 23752 29684 23780
rect 26476 23740 26482 23752
rect 15151 23684 16068 23712
rect 15151 23681 15163 23684
rect 15105 23675 15163 23681
rect 16942 23672 16948 23724
rect 17000 23712 17006 23724
rect 17037 23715 17095 23721
rect 17037 23712 17049 23715
rect 17000 23684 17049 23712
rect 17000 23672 17006 23684
rect 17037 23681 17049 23684
rect 17083 23712 17095 23715
rect 17494 23712 17500 23724
rect 17083 23684 17500 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 18690 23672 18696 23724
rect 18748 23672 18754 23724
rect 20438 23672 20444 23724
rect 20496 23712 20502 23724
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 20496 23684 21005 23712
rect 20496 23672 20502 23684
rect 20993 23681 21005 23684
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 29454 23672 29460 23724
rect 29512 23712 29518 23724
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 29512 23684 29561 23712
rect 29512 23672 29518 23684
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29656 23712 29684 23752
rect 30650 23740 30656 23792
rect 30708 23740 30714 23792
rect 30742 23740 30748 23792
rect 30800 23780 30806 23792
rect 32030 23780 32036 23792
rect 30800 23752 32036 23780
rect 30800 23740 30806 23752
rect 31496 23721 31524 23752
rect 32030 23740 32036 23752
rect 32088 23740 32094 23792
rect 33502 23740 33508 23792
rect 33560 23740 33566 23792
rect 33686 23740 33692 23792
rect 33744 23740 33750 23792
rect 31481 23715 31539 23721
rect 29656 23684 31432 23712
rect 29549 23675 29607 23681
rect 3970 23644 3976 23656
rect 2976 23616 3976 23644
rect 3970 23604 3976 23616
rect 4028 23604 4034 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6270 23604 6276 23656
rect 6328 23644 6334 23656
rect 7377 23647 7435 23653
rect 6328 23616 7328 23644
rect 6328 23604 6334 23616
rect 842 23536 848 23588
rect 900 23576 906 23588
rect 6733 23579 6791 23585
rect 6733 23576 6745 23579
rect 900 23548 2360 23576
rect 900 23536 906 23548
rect 1578 23468 1584 23520
rect 1636 23468 1642 23520
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 2225 23511 2283 23517
rect 2225 23508 2237 23511
rect 1820 23480 2237 23508
rect 1820 23468 1826 23480
rect 2225 23477 2237 23480
rect 2271 23477 2283 23511
rect 2332 23508 2360 23548
rect 2746 23548 6745 23576
rect 2746 23508 2774 23548
rect 6733 23545 6745 23548
rect 6779 23545 6791 23579
rect 7300 23576 7328 23616
rect 7377 23613 7389 23647
rect 7423 23644 7435 23647
rect 7558 23644 7564 23656
rect 7423 23616 7564 23644
rect 7423 23613 7435 23616
rect 7377 23607 7435 23613
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 12529 23647 12587 23653
rect 12529 23613 12541 23647
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 16117 23647 16175 23653
rect 16117 23613 16129 23647
rect 16163 23644 16175 23647
rect 18322 23644 18328 23656
rect 16163 23616 18328 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 12544 23576 12572 23607
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 18969 23647 19027 23653
rect 18969 23613 18981 23647
rect 19015 23644 19027 23647
rect 19058 23644 19064 23656
rect 19015 23616 19064 23644
rect 19015 23613 19027 23616
rect 18969 23607 19027 23613
rect 19058 23604 19064 23616
rect 19116 23604 19122 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 20088 23616 22017 23644
rect 17034 23576 17040 23588
rect 7300 23548 12434 23576
rect 12544 23548 17040 23576
rect 6733 23539 6791 23545
rect 2332 23480 2774 23508
rect 2225 23471 2283 23477
rect 3786 23468 3792 23520
rect 3844 23508 3850 23520
rect 9674 23508 9680 23520
rect 3844 23480 9680 23508
rect 3844 23468 3850 23480
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 11514 23468 11520 23520
rect 11572 23468 11578 23520
rect 11882 23468 11888 23520
rect 11940 23468 11946 23520
rect 12406 23508 12434 23548
rect 17034 23536 17040 23548
rect 17092 23536 17098 23588
rect 20088 23520 20116 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22278 23604 22284 23656
rect 22336 23604 22342 23656
rect 24394 23604 24400 23656
rect 24452 23644 24458 23656
rect 24857 23647 24915 23653
rect 24857 23644 24869 23647
rect 24452 23616 24869 23644
rect 24452 23604 24458 23616
rect 24857 23613 24869 23616
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23644 25191 23647
rect 25866 23644 25872 23656
rect 25179 23616 25872 23644
rect 25179 23613 25191 23616
rect 25133 23607 25191 23613
rect 25866 23604 25872 23616
rect 25924 23604 25930 23656
rect 27154 23604 27160 23656
rect 27212 23604 27218 23656
rect 27430 23604 27436 23656
rect 27488 23604 27494 23656
rect 31404 23644 31432 23684
rect 31481 23681 31493 23715
rect 31527 23712 31539 23715
rect 32214 23712 32220 23724
rect 31527 23684 31561 23712
rect 31726 23684 32220 23712
rect 31527 23681 31539 23684
rect 31481 23675 31539 23681
rect 31726 23644 31754 23684
rect 32214 23672 32220 23684
rect 32272 23672 32278 23724
rect 32306 23672 32312 23724
rect 32364 23672 32370 23724
rect 34348 23721 34376 23820
rect 34790 23808 34796 23860
rect 34848 23848 34854 23860
rect 36633 23851 36691 23857
rect 36633 23848 36645 23851
rect 34848 23820 36645 23848
rect 34848 23808 34854 23820
rect 36633 23817 36645 23820
rect 36679 23817 36691 23851
rect 36633 23811 36691 23817
rect 39298 23808 39304 23860
rect 39356 23808 39362 23860
rect 39942 23808 39948 23860
rect 40000 23848 40006 23860
rect 41049 23851 41107 23857
rect 41049 23848 41061 23851
rect 40000 23820 41061 23848
rect 40000 23808 40006 23820
rect 41049 23817 41061 23820
rect 41095 23817 41107 23851
rect 41049 23811 41107 23817
rect 45922 23808 45928 23860
rect 45980 23848 45986 23860
rect 46293 23851 46351 23857
rect 46293 23848 46305 23851
rect 45980 23820 46305 23848
rect 45980 23808 45986 23820
rect 46293 23817 46305 23820
rect 46339 23817 46351 23851
rect 46293 23811 46351 23817
rect 47302 23808 47308 23860
rect 47360 23848 47366 23860
rect 47581 23851 47639 23857
rect 47581 23848 47593 23851
rect 47360 23820 47593 23848
rect 47360 23808 47366 23820
rect 47581 23817 47593 23820
rect 47627 23817 47639 23851
rect 47581 23811 47639 23817
rect 47670 23808 47676 23860
rect 47728 23848 47734 23860
rect 48133 23851 48191 23857
rect 48133 23848 48145 23851
rect 47728 23820 48145 23848
rect 47728 23808 47734 23820
rect 48133 23817 48145 23820
rect 48179 23817 48191 23851
rect 48133 23811 48191 23817
rect 35986 23740 35992 23792
rect 36044 23740 36050 23792
rect 36170 23740 36176 23792
rect 36228 23740 36234 23792
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 36832 23752 37933 23780
rect 36832 23724 36860 23752
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 38470 23740 38476 23792
rect 38528 23740 38534 23792
rect 38654 23740 38660 23792
rect 38712 23740 38718 23792
rect 39209 23783 39267 23789
rect 39209 23749 39221 23783
rect 39255 23780 39267 23783
rect 40678 23780 40684 23792
rect 39255 23752 40684 23780
rect 39255 23749 39267 23752
rect 39209 23743 39267 23749
rect 40678 23740 40684 23752
rect 40736 23740 40742 23792
rect 43257 23783 43315 23789
rect 43257 23780 43269 23783
rect 41432 23752 43269 23780
rect 34333 23715 34391 23721
rect 34333 23681 34345 23715
rect 34379 23681 34391 23715
rect 34333 23675 34391 23681
rect 34514 23672 34520 23724
rect 34572 23712 34578 23724
rect 34793 23715 34851 23721
rect 34793 23712 34805 23715
rect 34572 23684 34805 23712
rect 34572 23672 34578 23684
rect 34793 23681 34805 23684
rect 34839 23681 34851 23715
rect 34793 23675 34851 23681
rect 36814 23672 36820 23724
rect 36872 23672 36878 23724
rect 37090 23672 37096 23724
rect 37148 23712 37154 23724
rect 37645 23715 37703 23721
rect 37645 23712 37657 23715
rect 37148 23684 37657 23712
rect 37148 23672 37154 23684
rect 37645 23681 37657 23684
rect 37691 23681 37703 23715
rect 37645 23675 37703 23681
rect 39574 23672 39580 23724
rect 39632 23712 39638 23724
rect 41432 23721 41460 23752
rect 43257 23749 43269 23752
rect 43303 23749 43315 23783
rect 43257 23743 43315 23749
rect 44082 23740 44088 23792
rect 44140 23780 44146 23792
rect 46201 23783 46259 23789
rect 46201 23780 46213 23783
rect 44140 23752 46213 23780
rect 44140 23740 44146 23752
rect 39945 23715 40003 23721
rect 39945 23712 39957 23715
rect 39632 23684 39957 23712
rect 39632 23672 39638 23684
rect 39945 23681 39957 23684
rect 39991 23712 40003 23715
rect 40865 23715 40923 23721
rect 40865 23712 40877 23715
rect 39991 23684 40877 23712
rect 39991 23681 40003 23684
rect 39945 23675 40003 23681
rect 40865 23681 40877 23684
rect 40911 23681 40923 23715
rect 40865 23675 40923 23681
rect 41417 23715 41475 23721
rect 41417 23681 41429 23715
rect 41463 23681 41475 23715
rect 41417 23675 41475 23681
rect 42610 23672 42616 23724
rect 42668 23672 42674 23724
rect 43717 23715 43775 23721
rect 43717 23681 43729 23715
rect 43763 23681 43775 23715
rect 43717 23675 43775 23681
rect 28460 23616 30880 23644
rect 31404 23616 31754 23644
rect 42061 23647 42119 23653
rect 26326 23536 26332 23588
rect 26384 23576 26390 23588
rect 26384 23548 26740 23576
rect 26384 23536 26390 23548
rect 14274 23508 14280 23520
rect 12406 23480 14280 23508
rect 14274 23468 14280 23480
rect 14332 23468 14338 23520
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 17678 23508 17684 23520
rect 16632 23480 17684 23508
rect 16632 23468 16638 23480
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 20070 23508 20076 23520
rect 18748 23480 20076 23508
rect 18748 23468 18754 23480
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20441 23511 20499 23517
rect 20441 23477 20453 23511
rect 20487 23508 20499 23511
rect 20530 23508 20536 23520
rect 20487 23480 20536 23508
rect 20487 23477 20499 23480
rect 20441 23471 20499 23477
rect 20530 23468 20536 23480
rect 20588 23468 20594 23520
rect 21634 23468 21640 23520
rect 21692 23468 21698 23520
rect 23750 23468 23756 23520
rect 23808 23468 23814 23520
rect 26602 23468 26608 23520
rect 26660 23468 26666 23520
rect 26712 23508 26740 23548
rect 28460 23508 28488 23616
rect 28534 23536 28540 23588
rect 28592 23576 28598 23588
rect 29365 23579 29423 23585
rect 29365 23576 29377 23579
rect 28592 23548 29377 23576
rect 28592 23536 28598 23548
rect 29365 23545 29377 23548
rect 29411 23545 29423 23579
rect 29365 23539 29423 23545
rect 29454 23536 29460 23588
rect 29512 23576 29518 23588
rect 30193 23579 30251 23585
rect 30193 23576 30205 23579
rect 29512 23548 30205 23576
rect 29512 23536 29518 23548
rect 30193 23545 30205 23548
rect 30239 23545 30251 23579
rect 30193 23539 30251 23545
rect 26712 23480 28488 23508
rect 28902 23468 28908 23520
rect 28960 23468 28966 23520
rect 29917 23511 29975 23517
rect 29917 23477 29929 23511
rect 29963 23508 29975 23511
rect 30098 23508 30104 23520
rect 29963 23480 30104 23508
rect 29963 23477 29975 23480
rect 29917 23471 29975 23477
rect 30098 23468 30104 23480
rect 30156 23468 30162 23520
rect 30374 23468 30380 23520
rect 30432 23508 30438 23520
rect 30745 23511 30803 23517
rect 30745 23508 30757 23511
rect 30432 23480 30757 23508
rect 30432 23468 30438 23480
rect 30745 23477 30757 23480
rect 30791 23477 30803 23511
rect 30852 23508 30880 23616
rect 42061 23613 42073 23647
rect 42107 23644 42119 23647
rect 43732 23644 43760 23675
rect 43806 23672 43812 23724
rect 43864 23712 43870 23724
rect 44634 23712 44640 23724
rect 43864 23684 44640 23712
rect 43864 23672 43870 23684
rect 44634 23672 44640 23684
rect 44692 23712 44698 23724
rect 45572 23721 45600 23752
rect 46201 23749 46213 23752
rect 46247 23749 46259 23783
rect 46201 23743 46259 23749
rect 44821 23715 44879 23721
rect 44821 23712 44833 23715
rect 44692 23684 44833 23712
rect 44692 23672 44698 23684
rect 44821 23681 44833 23684
rect 44867 23681 44879 23715
rect 44821 23675 44879 23681
rect 45557 23715 45615 23721
rect 45557 23681 45569 23715
rect 45603 23712 45615 23715
rect 45603 23684 45637 23712
rect 45603 23681 45615 23684
rect 45557 23675 45615 23681
rect 46658 23672 46664 23724
rect 46716 23712 46722 23724
rect 46753 23715 46811 23721
rect 46753 23712 46765 23715
rect 46716 23684 46765 23712
rect 46716 23672 46722 23684
rect 46753 23681 46765 23684
rect 46799 23712 46811 23715
rect 47305 23715 47363 23721
rect 47305 23712 47317 23715
rect 46799 23684 47317 23712
rect 46799 23681 46811 23684
rect 46753 23675 46811 23681
rect 47305 23681 47317 23684
rect 47351 23681 47363 23715
rect 47305 23675 47363 23681
rect 47762 23672 47768 23724
rect 47820 23712 47826 23724
rect 47949 23715 48007 23721
rect 47949 23712 47961 23715
rect 47820 23684 47961 23712
rect 47820 23672 47826 23684
rect 47949 23681 47961 23684
rect 47995 23712 48007 23715
rect 48314 23712 48320 23724
rect 47995 23684 48320 23712
rect 47995 23681 48007 23684
rect 47949 23675 48007 23681
rect 48314 23672 48320 23684
rect 48372 23672 48378 23724
rect 48682 23672 48688 23724
rect 48740 23672 48746 23724
rect 42107 23616 43760 23644
rect 42107 23613 42119 23616
rect 42061 23607 42119 23613
rect 31018 23536 31024 23588
rect 31076 23576 31082 23588
rect 37461 23579 37519 23585
rect 37461 23576 37473 23579
rect 31076 23548 37473 23576
rect 31076 23536 31082 23548
rect 37461 23545 37473 23548
rect 37507 23545 37519 23579
rect 44910 23576 44916 23588
rect 37461 23539 37519 23545
rect 37752 23548 44916 23576
rect 31297 23511 31355 23517
rect 31297 23508 31309 23511
rect 30852 23480 31309 23508
rect 30745 23471 30803 23477
rect 31297 23477 31309 23480
rect 31343 23477 31355 23511
rect 31297 23471 31355 23477
rect 31846 23468 31852 23520
rect 31904 23468 31910 23520
rect 32766 23468 32772 23520
rect 32824 23508 32830 23520
rect 32953 23511 33011 23517
rect 32953 23508 32965 23511
rect 32824 23480 32965 23508
rect 32824 23468 32830 23480
rect 32953 23477 32965 23480
rect 32999 23477 33011 23511
rect 32953 23471 33011 23477
rect 34054 23468 34060 23520
rect 34112 23508 34118 23520
rect 34149 23511 34207 23517
rect 34149 23508 34161 23511
rect 34112 23480 34161 23508
rect 34112 23468 34118 23480
rect 34149 23477 34161 23480
rect 34195 23477 34207 23511
rect 34149 23471 34207 23477
rect 35434 23468 35440 23520
rect 35492 23468 35498 23520
rect 36998 23468 37004 23520
rect 37056 23508 37062 23520
rect 37752 23508 37780 23548
rect 44910 23536 44916 23548
rect 44968 23536 44974 23588
rect 37056 23480 37780 23508
rect 37056 23468 37062 23480
rect 40586 23468 40592 23520
rect 40644 23468 40650 23520
rect 44358 23468 44364 23520
rect 44416 23468 44422 23520
rect 45002 23468 45008 23520
rect 45060 23468 45066 23520
rect 45738 23468 45744 23520
rect 45796 23468 45802 23520
rect 46934 23468 46940 23520
rect 46992 23468 46998 23520
rect 48682 23468 48688 23520
rect 48740 23508 48746 23520
rect 49329 23511 49387 23517
rect 49329 23508 49341 23511
rect 48740 23480 49341 23508
rect 48740 23468 48746 23480
rect 49329 23477 49341 23480
rect 49375 23477 49387 23511
rect 49329 23471 49387 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 3602 23264 3608 23316
rect 3660 23264 3666 23316
rect 3694 23264 3700 23316
rect 3752 23304 3758 23316
rect 3789 23307 3847 23313
rect 3789 23304 3801 23307
rect 3752 23276 3801 23304
rect 3752 23264 3758 23276
rect 3789 23273 3801 23276
rect 3835 23273 3847 23307
rect 3789 23267 3847 23273
rect 7742 23264 7748 23316
rect 7800 23304 7806 23316
rect 11057 23307 11115 23313
rect 11057 23304 11069 23307
rect 7800 23276 11069 23304
rect 7800 23264 7806 23276
rect 11057 23273 11069 23276
rect 11103 23304 11115 23307
rect 11774 23307 11832 23313
rect 11774 23304 11786 23307
rect 11103 23276 11786 23304
rect 11103 23273 11115 23276
rect 11057 23267 11115 23273
rect 11774 23273 11786 23276
rect 11820 23273 11832 23307
rect 11774 23267 11832 23273
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 13633 23307 13691 23313
rect 13633 23304 13645 23307
rect 12308 23276 13645 23304
rect 12308 23264 12314 23276
rect 13633 23273 13645 23276
rect 13679 23304 13691 23307
rect 13814 23304 13820 23316
rect 13679 23276 13820 23304
rect 13679 23273 13691 23276
rect 13633 23267 13691 23273
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 13909 23307 13967 23313
rect 13909 23273 13921 23307
rect 13955 23304 13967 23307
rect 19429 23307 19487 23313
rect 13955 23276 19380 23304
rect 13955 23273 13967 23276
rect 13909 23267 13967 23273
rect 8754 23236 8760 23248
rect 2746 23208 8760 23236
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 2746 23100 2774 23208
rect 8754 23196 8760 23208
rect 8812 23196 8818 23248
rect 13832 23236 13860 23264
rect 14921 23239 14979 23245
rect 14921 23236 14933 23239
rect 13832 23208 14933 23236
rect 14921 23205 14933 23208
rect 14967 23205 14979 23239
rect 14921 23199 14979 23205
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 19058 23236 19064 23248
rect 18923 23208 19064 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 19058 23196 19064 23208
rect 19116 23196 19122 23248
rect 19352 23236 19380 23276
rect 19429 23273 19441 23307
rect 19475 23304 19487 23307
rect 23290 23304 23296 23316
rect 19475 23276 23296 23304
rect 19475 23273 19487 23276
rect 19429 23267 19487 23273
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 23842 23264 23848 23316
rect 23900 23304 23906 23316
rect 25777 23307 25835 23313
rect 25777 23304 25789 23307
rect 23900 23276 25789 23304
rect 23900 23264 23906 23276
rect 25777 23273 25789 23276
rect 25823 23273 25835 23307
rect 28534 23304 28540 23316
rect 25777 23267 25835 23273
rect 25884 23276 26372 23304
rect 19352 23208 20208 23236
rect 3421 23171 3479 23177
rect 3421 23137 3433 23171
rect 3467 23168 3479 23171
rect 4062 23168 4068 23180
rect 3467 23140 4068 23168
rect 3467 23137 3479 23140
rect 3421 23131 3479 23137
rect 4062 23128 4068 23140
rect 4120 23128 4126 23180
rect 4801 23171 4859 23177
rect 4801 23137 4813 23171
rect 4847 23168 4859 23171
rect 4982 23168 4988 23180
rect 4847 23140 4988 23168
rect 4847 23137 4859 23140
rect 4801 23131 4859 23137
rect 4982 23128 4988 23140
rect 5040 23128 5046 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 12434 23168 12440 23180
rect 11563 23140 12440 23168
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 13262 23128 13268 23180
rect 13320 23168 13326 23180
rect 15838 23168 15844 23180
rect 13320 23140 15844 23168
rect 13320 23128 13326 23140
rect 15838 23128 15844 23140
rect 15896 23128 15902 23180
rect 16485 23171 16543 23177
rect 16485 23137 16497 23171
rect 16531 23168 16543 23171
rect 17402 23168 17408 23180
rect 16531 23140 17408 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 20070 23128 20076 23180
rect 20128 23128 20134 23180
rect 20180 23168 20208 23208
rect 23750 23196 23756 23248
rect 23808 23236 23814 23248
rect 25884 23236 25912 23276
rect 23808 23208 25912 23236
rect 23808 23196 23814 23208
rect 20714 23168 20720 23180
rect 20180 23140 20720 23168
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 22557 23171 22615 23177
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 23768 23168 23796 23196
rect 22603 23140 23796 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 26344 23177 26372 23276
rect 27080 23276 28540 23304
rect 26329 23171 26387 23177
rect 26329 23137 26341 23171
rect 26375 23137 26387 23171
rect 26329 23131 26387 23137
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 1811 23072 2774 23100
rect 4816 23072 5365 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 4816 23044 4844 23072
rect 5353 23069 5365 23072
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 7190 23060 7196 23112
rect 7248 23060 7254 23112
rect 8938 23060 8944 23112
rect 8996 23100 9002 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 8996 23072 9321 23100
rect 8996 23060 9002 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 13096 23072 14504 23100
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 4065 23035 4123 23041
rect 4065 23001 4077 23035
rect 4111 23032 4123 23035
rect 4522 23032 4528 23044
rect 4111 23004 4528 23032
rect 4111 23001 4123 23004
rect 4065 22995 4123 23001
rect 4522 22992 4528 23004
rect 4580 22992 4586 23044
rect 4798 22992 4804 23044
rect 4856 22992 4862 23044
rect 9490 22992 9496 23044
rect 9548 23032 9554 23044
rect 9585 23035 9643 23041
rect 9585 23032 9597 23035
rect 9548 23004 9597 23032
rect 9548 22992 9554 23004
rect 9585 23001 9597 23004
rect 9631 23001 9643 23035
rect 12250 23032 12256 23044
rect 9585 22995 9643 23001
rect 9968 23004 10074 23032
rect 11532 23004 12256 23032
rect 4154 22924 4160 22976
rect 4212 22924 4218 22976
rect 4617 22967 4675 22973
rect 4617 22933 4629 22967
rect 4663 22964 4675 22967
rect 7098 22964 7104 22976
rect 4663 22936 7104 22964
rect 4663 22933 4675 22936
rect 4617 22927 4675 22933
rect 7098 22924 7104 22936
rect 7156 22924 7162 22976
rect 9030 22924 9036 22976
rect 9088 22964 9094 22976
rect 9968 22964 9996 23004
rect 11532 22976 11560 23004
rect 12250 22992 12256 23004
rect 12308 22992 12314 23044
rect 11514 22964 11520 22976
rect 9088 22936 11520 22964
rect 9088 22924 9094 22936
rect 11514 22924 11520 22936
rect 11572 22924 11578 22976
rect 11974 22924 11980 22976
rect 12032 22964 12038 22976
rect 12618 22964 12624 22976
rect 12032 22936 12624 22964
rect 12032 22924 12038 22936
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 13096 22964 13124 23072
rect 13630 22992 13636 23044
rect 13688 23032 13694 23044
rect 14366 23032 14372 23044
rect 13688 23004 14372 23032
rect 13688 22992 13694 23004
rect 14366 22992 14372 23004
rect 14424 22992 14430 23044
rect 14476 23032 14504 23072
rect 15470 23060 15476 23112
rect 15528 23060 15534 23112
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 16908 23072 17141 23100
rect 16908 23060 16914 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 18506 23060 18512 23112
rect 18564 23060 18570 23112
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23100 19671 23103
rect 19794 23100 19800 23112
rect 19659 23072 19800 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 19794 23060 19800 23072
rect 19852 23060 19858 23112
rect 21726 23060 21732 23112
rect 21784 23100 21790 23112
rect 22281 23103 22339 23109
rect 22281 23100 22293 23103
rect 21784 23072 22293 23100
rect 21784 23060 21790 23072
rect 22281 23069 22293 23072
rect 22327 23069 22339 23103
rect 22281 23063 22339 23069
rect 23658 23060 23664 23112
rect 23716 23060 23722 23112
rect 26237 23103 26295 23109
rect 26237 23069 26249 23103
rect 26283 23100 26295 23103
rect 27080 23100 27108 23276
rect 28534 23264 28540 23276
rect 28592 23264 28598 23316
rect 28994 23264 29000 23316
rect 29052 23264 29058 23316
rect 29365 23307 29423 23313
rect 29365 23273 29377 23307
rect 29411 23304 29423 23307
rect 29454 23304 29460 23316
rect 29411 23276 29460 23304
rect 29411 23273 29423 23276
rect 29365 23267 29423 23273
rect 29454 23264 29460 23276
rect 29512 23264 29518 23316
rect 29822 23264 29828 23316
rect 29880 23304 29886 23316
rect 30098 23304 30104 23316
rect 29880 23276 30104 23304
rect 29880 23264 29886 23276
rect 30098 23264 30104 23276
rect 30156 23304 30162 23316
rect 31846 23304 31852 23316
rect 30156 23276 31852 23304
rect 30156 23264 30162 23276
rect 31846 23264 31852 23276
rect 31904 23264 31910 23316
rect 32214 23264 32220 23316
rect 32272 23304 32278 23316
rect 33597 23307 33655 23313
rect 33597 23304 33609 23307
rect 32272 23276 33609 23304
rect 32272 23264 32278 23276
rect 33597 23273 33609 23276
rect 33643 23273 33655 23307
rect 33597 23267 33655 23273
rect 33870 23264 33876 23316
rect 33928 23304 33934 23316
rect 34149 23307 34207 23313
rect 34149 23304 34161 23307
rect 33928 23276 34161 23304
rect 33928 23264 33934 23276
rect 34149 23273 34161 23276
rect 34195 23273 34207 23307
rect 34149 23267 34207 23273
rect 38562 23264 38568 23316
rect 38620 23304 38626 23316
rect 39577 23307 39635 23313
rect 39577 23304 39589 23307
rect 38620 23276 39589 23304
rect 38620 23264 38626 23276
rect 39577 23273 39589 23276
rect 39623 23273 39635 23307
rect 39577 23267 39635 23273
rect 43993 23307 44051 23313
rect 43993 23273 44005 23307
rect 44039 23304 44051 23307
rect 44174 23304 44180 23316
rect 44039 23276 44180 23304
rect 44039 23273 44051 23276
rect 43993 23267 44051 23273
rect 44174 23264 44180 23276
rect 44232 23264 44238 23316
rect 44634 23264 44640 23316
rect 44692 23264 44698 23316
rect 48590 23264 48596 23316
rect 48648 23304 48654 23316
rect 49329 23307 49387 23313
rect 49329 23304 49341 23307
rect 48648 23276 49341 23304
rect 48648 23264 48654 23276
rect 49329 23273 49341 23276
rect 49375 23273 49387 23307
rect 49329 23267 49387 23273
rect 29012 23236 29040 23264
rect 29012 23208 29868 23236
rect 27246 23128 27252 23180
rect 27304 23128 27310 23180
rect 27525 23171 27583 23177
rect 27525 23137 27537 23171
rect 27571 23168 27583 23171
rect 28902 23168 28908 23180
rect 27571 23140 28908 23168
rect 27571 23137 27583 23140
rect 27525 23131 27583 23137
rect 28902 23128 28908 23140
rect 28960 23168 28966 23180
rect 29840 23168 29868 23208
rect 32490 23196 32496 23248
rect 32548 23236 32554 23248
rect 37090 23236 37096 23248
rect 32548 23208 37096 23236
rect 32548 23196 32554 23208
rect 37090 23196 37096 23208
rect 37148 23196 37154 23248
rect 30009 23171 30067 23177
rect 30009 23168 30021 23171
rect 28960 23140 29500 23168
rect 29840 23140 30021 23168
rect 28960 23128 28966 23140
rect 29362 23100 29368 23112
rect 26283 23072 27108 23100
rect 28658 23072 29368 23100
rect 26283 23069 26295 23072
rect 26237 23063 26295 23069
rect 29362 23060 29368 23072
rect 29420 23060 29426 23112
rect 16942 23032 16948 23044
rect 14476 23004 16948 23032
rect 16942 22992 16948 23004
rect 17000 22992 17006 23044
rect 17034 22992 17040 23044
rect 17092 23032 17098 23044
rect 17405 23035 17463 23041
rect 17405 23032 17417 23035
rect 17092 23004 17417 23032
rect 17092 22992 17098 23004
rect 17405 23001 17417 23004
rect 17451 23001 17463 23035
rect 17405 22995 17463 23001
rect 20346 22992 20352 23044
rect 20404 22992 20410 23044
rect 21634 23032 21640 23044
rect 21574 23004 21640 23032
rect 21634 22992 21640 23004
rect 21692 22992 21698 23044
rect 25041 23035 25099 23041
rect 25041 23001 25053 23035
rect 25087 23032 25099 23035
rect 29472 23032 29500 23140
rect 30009 23137 30021 23140
rect 30055 23137 30067 23171
rect 30009 23131 30067 23137
rect 30742 23128 30748 23180
rect 30800 23168 30806 23180
rect 31481 23171 31539 23177
rect 31481 23168 31493 23171
rect 30800 23140 31493 23168
rect 30800 23128 30806 23140
rect 31481 23137 31493 23140
rect 31527 23137 31539 23171
rect 31481 23131 31539 23137
rect 31938 23128 31944 23180
rect 31996 23168 32002 23180
rect 36814 23168 36820 23180
rect 31996 23140 36820 23168
rect 31996 23128 32002 23140
rect 36814 23128 36820 23140
rect 36872 23128 36878 23180
rect 40037 23171 40095 23177
rect 40037 23137 40049 23171
rect 40083 23168 40095 23171
rect 40586 23168 40592 23180
rect 40083 23140 40592 23168
rect 40083 23137 40095 23140
rect 40037 23131 40095 23137
rect 40586 23128 40592 23140
rect 40644 23128 40650 23180
rect 47489 23171 47547 23177
rect 47489 23137 47501 23171
rect 47535 23168 47547 23171
rect 47535 23140 48544 23168
rect 47535 23137 47547 23140
rect 47489 23131 47547 23137
rect 48516 23112 48544 23140
rect 29730 23060 29736 23112
rect 29788 23060 29794 23112
rect 32125 23103 32183 23109
rect 32125 23069 32137 23103
rect 32171 23100 32183 23103
rect 32398 23100 32404 23112
rect 32171 23072 32404 23100
rect 32171 23069 32183 23072
rect 32125 23063 32183 23069
rect 32398 23060 32404 23072
rect 32456 23060 32462 23112
rect 32674 23060 32680 23112
rect 32732 23100 32738 23112
rect 32732 23072 33088 23100
rect 32732 23060 32738 23072
rect 29914 23032 29920 23044
rect 25087 23004 27476 23032
rect 25087 23001 25099 23004
rect 25041 22995 25099 23001
rect 12860 22936 13124 22964
rect 12860 22924 12866 22936
rect 14458 22924 14464 22976
rect 14516 22924 14522 22976
rect 17218 22924 17224 22976
rect 17276 22964 17282 22976
rect 21821 22967 21879 22973
rect 21821 22964 21833 22967
rect 17276 22936 21833 22964
rect 17276 22924 17282 22936
rect 21821 22933 21833 22936
rect 21867 22964 21879 22967
rect 22278 22964 22284 22976
rect 21867 22936 22284 22964
rect 21867 22933 21879 22936
rect 21821 22927 21879 22933
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 23382 22924 23388 22976
rect 23440 22964 23446 22976
rect 24029 22967 24087 22973
rect 24029 22964 24041 22967
rect 23440 22936 24041 22964
rect 23440 22924 23446 22936
rect 24029 22933 24041 22936
rect 24075 22933 24087 22967
rect 24029 22927 24087 22933
rect 24118 22924 24124 22976
rect 24176 22964 24182 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 24176 22936 24593 22964
rect 24176 22924 24182 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 24670 22924 24676 22976
rect 24728 22964 24734 22976
rect 24949 22967 25007 22973
rect 24949 22964 24961 22967
rect 24728 22936 24961 22964
rect 24728 22924 24734 22936
rect 24949 22933 24961 22936
rect 24995 22933 25007 22967
rect 24949 22927 25007 22933
rect 25866 22924 25872 22976
rect 25924 22964 25930 22976
rect 26145 22967 26203 22973
rect 26145 22964 26157 22967
rect 25924 22936 26157 22964
rect 25924 22924 25930 22936
rect 26145 22933 26157 22936
rect 26191 22964 26203 22967
rect 26786 22964 26792 22976
rect 26191 22936 26792 22964
rect 26191 22933 26203 22936
rect 26145 22927 26203 22933
rect 26786 22924 26792 22936
rect 26844 22924 26850 22976
rect 26881 22967 26939 22973
rect 26881 22933 26893 22967
rect 26927 22964 26939 22967
rect 26970 22964 26976 22976
rect 26927 22936 26976 22964
rect 26927 22933 26939 22936
rect 26881 22927 26939 22933
rect 26970 22924 26976 22936
rect 27028 22924 27034 22976
rect 27448 22964 27476 23004
rect 28920 23004 29408 23032
rect 29472 23004 29920 23032
rect 28920 22964 28948 23004
rect 27448 22936 28948 22964
rect 29380 22964 29408 23004
rect 29914 22992 29920 23004
rect 29972 22992 29978 23044
rect 31478 23032 31484 23044
rect 31234 23004 31484 23032
rect 31478 22992 31484 23004
rect 31536 22992 31542 23044
rect 33060 23032 33088 23072
rect 33134 23060 33140 23112
rect 33192 23100 33198 23112
rect 33870 23100 33876 23112
rect 33192 23072 33876 23100
rect 33192 23060 33198 23072
rect 33870 23060 33876 23072
rect 33928 23060 33934 23112
rect 34057 23103 34115 23109
rect 34057 23069 34069 23103
rect 34103 23100 34115 23103
rect 34146 23100 34152 23112
rect 34103 23072 34152 23100
rect 34103 23069 34115 23072
rect 34057 23063 34115 23069
rect 34146 23060 34152 23072
rect 34204 23060 34210 23112
rect 34977 23103 35035 23109
rect 34977 23069 34989 23103
rect 35023 23100 35035 23103
rect 35434 23100 35440 23112
rect 35023 23072 35440 23100
rect 35023 23069 35035 23072
rect 34977 23063 35035 23069
rect 35434 23060 35440 23072
rect 35492 23060 35498 23112
rect 35710 23060 35716 23112
rect 35768 23100 35774 23112
rect 38933 23103 38991 23109
rect 38933 23100 38945 23103
rect 35768 23072 38945 23100
rect 35768 23060 35774 23072
rect 38933 23069 38945 23072
rect 38979 23100 38991 23103
rect 39209 23103 39267 23109
rect 39209 23100 39221 23103
rect 38979 23072 39221 23100
rect 38979 23069 38991 23072
rect 38933 23063 38991 23069
rect 39209 23069 39221 23072
rect 39255 23069 39267 23103
rect 39209 23063 39267 23069
rect 40310 23060 40316 23112
rect 40368 23060 40374 23112
rect 42889 23103 42947 23109
rect 42889 23069 42901 23103
rect 42935 23100 42947 23103
rect 43254 23100 43260 23112
rect 42935 23072 43260 23100
rect 42935 23069 42947 23072
rect 42889 23063 42947 23069
rect 43254 23060 43260 23072
rect 43312 23060 43318 23112
rect 43349 23103 43407 23109
rect 43349 23069 43361 23103
rect 43395 23100 43407 23103
rect 44358 23100 44364 23112
rect 43395 23072 44364 23100
rect 43395 23069 43407 23072
rect 43349 23063 43407 23069
rect 44358 23060 44364 23072
rect 44416 23060 44422 23112
rect 46201 23103 46259 23109
rect 46201 23069 46213 23103
rect 46247 23069 46259 23103
rect 46201 23063 46259 23069
rect 47673 23103 47731 23109
rect 47673 23069 47685 23103
rect 47719 23100 47731 23103
rect 47854 23100 47860 23112
rect 47719 23072 47860 23100
rect 47719 23069 47731 23072
rect 47673 23063 47731 23069
rect 33413 23035 33471 23041
rect 33413 23032 33425 23035
rect 33060 23004 33425 23032
rect 33413 23001 33425 23004
rect 33459 23001 33471 23035
rect 33413 22995 33471 23001
rect 31941 22967 31999 22973
rect 31941 22964 31953 22967
rect 29380 22936 31953 22964
rect 31941 22933 31953 22936
rect 31987 22933 31999 22967
rect 31941 22927 31999 22933
rect 32030 22924 32036 22976
rect 32088 22964 32094 22976
rect 32401 22967 32459 22973
rect 32401 22964 32413 22967
rect 32088 22936 32413 22964
rect 32088 22924 32094 22936
rect 32401 22933 32413 22936
rect 32447 22933 32459 22967
rect 32401 22927 32459 22933
rect 32582 22924 32588 22976
rect 32640 22924 32646 22976
rect 32950 22924 32956 22976
rect 33008 22924 33014 22976
rect 33428 22964 33456 22995
rect 33502 22992 33508 23044
rect 33560 23032 33566 23044
rect 35161 23035 35219 23041
rect 35161 23032 35173 23035
rect 33560 23004 35173 23032
rect 33560 22992 33566 23004
rect 35161 23001 35173 23004
rect 35207 23001 35219 23035
rect 35161 22995 35219 23001
rect 35618 22992 35624 23044
rect 35676 22992 35682 23044
rect 36541 23035 36599 23041
rect 36541 23001 36553 23035
rect 36587 23032 36599 23035
rect 46216 23032 46244 23063
rect 47854 23060 47860 23072
rect 47912 23100 47918 23112
rect 47949 23103 48007 23109
rect 47949 23100 47961 23103
rect 47912 23072 47961 23100
rect 47912 23060 47918 23072
rect 47949 23069 47961 23072
rect 47995 23069 48007 23103
rect 47949 23063 48007 23069
rect 48498 23060 48504 23112
rect 48556 23100 48562 23112
rect 48685 23103 48743 23109
rect 48685 23100 48697 23103
rect 48556 23072 48697 23100
rect 48556 23060 48562 23072
rect 48685 23069 48697 23072
rect 48731 23069 48743 23103
rect 48685 23063 48743 23069
rect 48406 23032 48412 23044
rect 36587 23004 42748 23032
rect 46216 23004 48412 23032
rect 36587 23001 36599 23004
rect 36541 22995 36599 23001
rect 36081 22967 36139 22973
rect 36081 22964 36093 22967
rect 33428 22936 36093 22964
rect 36081 22933 36093 22936
rect 36127 22964 36139 22967
rect 37458 22964 37464 22976
rect 36127 22936 37464 22964
rect 36127 22933 36139 22936
rect 36081 22927 36139 22933
rect 37458 22924 37464 22936
rect 37516 22964 37522 22976
rect 37829 22967 37887 22973
rect 37829 22964 37841 22967
rect 37516 22936 37841 22964
rect 37516 22924 37522 22936
rect 37829 22933 37841 22936
rect 37875 22933 37887 22967
rect 37829 22927 37887 22933
rect 38746 22924 38752 22976
rect 38804 22924 38810 22976
rect 42720 22973 42748 23004
rect 48406 22992 48412 23004
rect 48464 22992 48470 23044
rect 42705 22967 42763 22973
rect 42705 22933 42717 22967
rect 42751 22933 42763 22967
rect 42705 22927 42763 22933
rect 46842 22924 46848 22976
rect 46900 22924 46906 22976
rect 47486 22924 47492 22976
rect 47544 22964 47550 22976
rect 48133 22967 48191 22973
rect 48133 22964 48145 22967
rect 47544 22936 48145 22964
rect 47544 22924 47550 22936
rect 48133 22933 48145 22936
rect 48179 22933 48191 22967
rect 48133 22927 48191 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 14458 22760 14464 22772
rect 2746 22732 14464 22760
rect 2746 22692 2774 22732
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 18598 22720 18604 22772
rect 18656 22720 18662 22772
rect 20346 22720 20352 22772
rect 20404 22760 20410 22772
rect 21453 22763 21511 22769
rect 21453 22760 21465 22763
rect 20404 22732 21465 22760
rect 20404 22720 20410 22732
rect 21453 22729 21465 22732
rect 21499 22760 21511 22763
rect 25130 22760 25136 22772
rect 21499 22732 25136 22760
rect 21499 22729 21511 22732
rect 21453 22723 21511 22729
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 25777 22763 25835 22769
rect 25777 22729 25789 22763
rect 25823 22760 25835 22763
rect 26326 22760 26332 22772
rect 25823 22732 26332 22760
rect 25823 22729 25835 22732
rect 25777 22723 25835 22729
rect 26326 22720 26332 22732
rect 26384 22720 26390 22772
rect 26418 22720 26424 22772
rect 26476 22720 26482 22772
rect 27522 22720 27528 22772
rect 27580 22760 27586 22772
rect 27617 22763 27675 22769
rect 27617 22760 27629 22763
rect 27580 22732 27629 22760
rect 27580 22720 27586 22732
rect 27617 22729 27629 22732
rect 27663 22729 27675 22763
rect 30742 22760 30748 22772
rect 27617 22723 27675 22729
rect 28644 22732 30748 22760
rect 1780 22664 2774 22692
rect 4816 22664 6500 22692
rect 1780 22633 1808 22664
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22593 1823 22627
rect 1765 22587 1823 22593
rect 3786 22584 3792 22636
rect 3844 22584 3850 22636
rect 4816 22633 4844 22664
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 6362 22624 6368 22636
rect 4801 22587 4859 22593
rect 5000 22596 6368 22624
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3326 22516 3332 22568
rect 3384 22556 3390 22568
rect 3881 22559 3939 22565
rect 3881 22556 3893 22559
rect 3384 22528 3893 22556
rect 3384 22516 3390 22528
rect 3881 22525 3893 22528
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22556 4123 22559
rect 5000 22556 5028 22596
rect 6362 22584 6368 22596
rect 6420 22584 6426 22636
rect 4111 22528 5028 22556
rect 4111 22525 4123 22528
rect 4065 22519 4123 22525
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 6472 22556 6500 22664
rect 7006 22652 7012 22704
rect 7064 22692 7070 22704
rect 7064 22664 7972 22692
rect 7064 22652 7070 22664
rect 6822 22584 6828 22636
rect 6880 22624 6886 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 6880 22596 7113 22624
rect 6880 22584 6886 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22624 7251 22627
rect 7834 22624 7840 22636
rect 7239 22596 7840 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 7944 22633 7972 22664
rect 10686 22652 10692 22704
rect 10744 22652 10750 22704
rect 10962 22652 10968 22704
rect 11020 22692 11026 22704
rect 12802 22692 12808 22704
rect 11020 22664 12808 22692
rect 11020 22652 11026 22664
rect 12802 22652 12808 22664
rect 12860 22652 12866 22704
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 16666 22652 16672 22704
rect 16724 22692 16730 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16724 22664 17141 22692
rect 16724 22652 16730 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 18506 22692 18512 22704
rect 18354 22664 18512 22692
rect 17129 22655 17187 22661
rect 18506 22652 18512 22664
rect 18564 22652 18570 22704
rect 20070 22692 20076 22704
rect 19720 22664 20076 22692
rect 7929 22627 7987 22633
rect 7929 22593 7941 22627
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 9766 22584 9772 22636
rect 9824 22584 9830 22636
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 12250 22624 12256 22636
rect 11839 22596 12256 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 13814 22584 13820 22636
rect 13872 22624 13878 22636
rect 14553 22627 14611 22633
rect 14553 22624 14565 22627
rect 13872 22596 14565 22624
rect 13872 22584 13878 22596
rect 14553 22593 14565 22596
rect 14599 22593 14611 22627
rect 14553 22587 14611 22593
rect 15010 22584 15016 22636
rect 15068 22584 15074 22636
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19720 22633 19748 22664
rect 20070 22652 20076 22664
rect 20128 22652 20134 22704
rect 21634 22692 21640 22704
rect 21206 22664 21640 22692
rect 21634 22652 21640 22664
rect 21692 22692 21698 22704
rect 22189 22695 22247 22701
rect 22189 22692 22201 22695
rect 21692 22664 22201 22692
rect 21692 22652 21698 22664
rect 22189 22661 22201 22664
rect 22235 22692 22247 22695
rect 23658 22692 23664 22704
rect 22235 22664 23664 22692
rect 22235 22661 22247 22664
rect 22189 22655 22247 22661
rect 23658 22652 23664 22664
rect 23716 22692 23722 22704
rect 23716 22664 23874 22692
rect 23716 22652 23722 22664
rect 24670 22652 24676 22704
rect 24728 22692 24734 22704
rect 26513 22695 26571 22701
rect 26513 22692 26525 22695
rect 24728 22664 26525 22692
rect 24728 22652 24734 22664
rect 26513 22661 26525 22664
rect 26559 22692 26571 22695
rect 26602 22692 26608 22704
rect 26559 22664 26608 22692
rect 26559 22661 26571 22664
rect 26513 22655 26571 22661
rect 26602 22652 26608 22664
rect 26660 22652 26666 22704
rect 26786 22652 26792 22704
rect 26844 22692 26850 22704
rect 28350 22692 28356 22704
rect 26844 22664 28356 22692
rect 26844 22652 26850 22664
rect 19705 22627 19763 22633
rect 19705 22624 19717 22627
rect 19484 22596 19717 22624
rect 19484 22584 19490 22596
rect 19705 22593 19717 22596
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22624 22523 22627
rect 22830 22624 22836 22636
rect 22511 22596 22836 22624
rect 22511 22593 22523 22596
rect 22465 22587 22523 22593
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 25498 22584 25504 22636
rect 25556 22624 25562 22636
rect 25685 22627 25743 22633
rect 25685 22624 25697 22627
rect 25556 22596 25697 22624
rect 25556 22584 25562 22596
rect 25685 22593 25697 22596
rect 25731 22624 25743 22627
rect 26970 22624 26976 22636
rect 25731 22596 26976 22624
rect 25731 22593 25743 22596
rect 25685 22587 25743 22593
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 27540 22633 27568 22664
rect 28350 22652 28356 22664
rect 28408 22692 28414 22704
rect 28534 22692 28540 22704
rect 28408 22664 28540 22692
rect 28408 22652 28414 22664
rect 28534 22652 28540 22664
rect 28592 22652 28598 22704
rect 28644 22701 28672 22732
rect 30742 22720 30748 22732
rect 30800 22720 30806 22772
rect 31018 22720 31024 22772
rect 31076 22720 31082 22772
rect 32950 22760 32956 22772
rect 31128 22732 32956 22760
rect 28629 22695 28687 22701
rect 28629 22661 28641 22695
rect 28675 22661 28687 22695
rect 28629 22655 28687 22661
rect 29362 22652 29368 22704
rect 29420 22652 29426 22704
rect 30834 22652 30840 22704
rect 30892 22692 30898 22704
rect 31128 22692 31156 22732
rect 32950 22720 32956 22732
rect 33008 22720 33014 22772
rect 33229 22763 33287 22769
rect 33229 22729 33241 22763
rect 33275 22760 33287 22763
rect 33410 22760 33416 22772
rect 33275 22732 33416 22760
rect 33275 22729 33287 22732
rect 33229 22723 33287 22729
rect 33410 22720 33416 22732
rect 33468 22720 33474 22772
rect 34514 22720 34520 22772
rect 34572 22760 34578 22772
rect 36817 22763 36875 22769
rect 36817 22760 36829 22763
rect 34572 22732 36829 22760
rect 34572 22720 34578 22732
rect 36817 22729 36829 22732
rect 36863 22729 36875 22763
rect 36817 22723 36875 22729
rect 37458 22720 37464 22772
rect 37516 22720 37522 22772
rect 40862 22720 40868 22772
rect 40920 22760 40926 22772
rect 40920 22732 41414 22760
rect 40920 22720 40926 22732
rect 30892 22664 31156 22692
rect 30892 22652 30898 22664
rect 31386 22652 31392 22704
rect 31444 22692 31450 22704
rect 33781 22695 33839 22701
rect 33781 22692 33793 22695
rect 31444 22664 33793 22692
rect 31444 22652 31450 22664
rect 33781 22661 33793 22664
rect 33827 22661 33839 22695
rect 33781 22655 33839 22661
rect 36538 22652 36544 22704
rect 36596 22652 36602 22704
rect 37476 22692 37504 22720
rect 41386 22692 41414 22732
rect 43254 22720 43260 22772
rect 43312 22720 43318 22772
rect 47762 22720 47768 22772
rect 47820 22720 47826 22772
rect 41785 22695 41843 22701
rect 41785 22692 41797 22695
rect 37476 22664 38594 22692
rect 41386 22664 41797 22692
rect 27525 22627 27583 22633
rect 27525 22593 27537 22627
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 27632 22596 28396 22624
rect 6472 22528 6868 22556
rect 3694 22448 3700 22500
rect 3752 22488 3758 22500
rect 4614 22488 4620 22500
rect 3752 22460 4620 22488
rect 3752 22448 3758 22460
rect 4614 22448 4620 22460
rect 4672 22448 4678 22500
rect 5718 22448 5724 22500
rect 5776 22488 5782 22500
rect 6733 22491 6791 22497
rect 6733 22488 6745 22491
rect 5776 22460 6745 22488
rect 5776 22448 5782 22460
rect 6733 22457 6745 22460
rect 6779 22457 6791 22491
rect 6840 22488 6868 22528
rect 7282 22516 7288 22568
rect 7340 22516 7346 22568
rect 8662 22516 8668 22568
rect 8720 22516 8726 22568
rect 8754 22516 8760 22568
rect 8812 22556 8818 22568
rect 11974 22556 11980 22568
rect 8812 22528 11980 22556
rect 8812 22516 8818 22528
rect 11974 22516 11980 22528
rect 12032 22516 12038 22568
rect 12434 22516 12440 22568
rect 12492 22516 12498 22568
rect 12713 22559 12771 22565
rect 12713 22556 12725 22559
rect 12544 22528 12725 22556
rect 9582 22488 9588 22500
rect 6840 22460 9588 22488
rect 6733 22451 6791 22457
rect 9582 22448 9588 22460
rect 9640 22448 9646 22500
rect 10870 22448 10876 22500
rect 10928 22488 10934 22500
rect 12544 22488 12572 22528
rect 12713 22525 12725 22528
rect 12759 22556 12771 22559
rect 13262 22556 13268 22568
rect 12759 22528 13268 22556
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 13262 22516 13268 22528
rect 13320 22516 13326 22568
rect 16850 22516 16856 22568
rect 16908 22516 16914 22568
rect 18598 22516 18604 22568
rect 18656 22556 18662 22568
rect 19981 22559 20039 22565
rect 19981 22556 19993 22559
rect 18656 22528 19993 22556
rect 18656 22516 18662 22528
rect 19981 22525 19993 22528
rect 20027 22556 20039 22559
rect 20530 22556 20536 22568
rect 20027 22528 20536 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 21726 22516 21732 22568
rect 21784 22556 21790 22568
rect 21913 22559 21971 22565
rect 21913 22556 21925 22559
rect 21784 22528 21925 22556
rect 21784 22516 21790 22528
rect 21913 22525 21925 22528
rect 21959 22556 21971 22559
rect 23109 22559 23167 22565
rect 23109 22556 23121 22559
rect 21959 22528 23121 22556
rect 21959 22525 21971 22528
rect 21913 22519 21971 22525
rect 23109 22525 23121 22528
rect 23155 22525 23167 22559
rect 23109 22519 23167 22525
rect 23382 22516 23388 22568
rect 23440 22516 23446 22568
rect 23750 22516 23756 22568
rect 23808 22556 23814 22568
rect 24026 22556 24032 22568
rect 23808 22528 24032 22556
rect 23808 22516 23814 22528
rect 24026 22516 24032 22528
rect 24084 22516 24090 22568
rect 25869 22559 25927 22565
rect 25869 22525 25881 22559
rect 25915 22525 25927 22559
rect 25869 22519 25927 22525
rect 25884 22488 25912 22519
rect 27246 22516 27252 22568
rect 27304 22556 27310 22568
rect 27632 22556 27660 22596
rect 28368 22568 28396 22596
rect 29914 22584 29920 22636
rect 29972 22624 29978 22636
rect 30929 22627 30987 22633
rect 29972 22596 30236 22624
rect 29972 22584 29978 22596
rect 27304 22528 27660 22556
rect 27709 22559 27767 22565
rect 27304 22516 27310 22528
rect 27709 22525 27721 22559
rect 27755 22525 27767 22559
rect 27709 22519 27767 22525
rect 10928 22460 12572 22488
rect 24872 22460 25912 22488
rect 10928 22448 10934 22460
rect 3421 22423 3479 22429
rect 3421 22389 3433 22423
rect 3467 22420 3479 22423
rect 5350 22420 5356 22432
rect 3467 22392 5356 22420
rect 3467 22389 3479 22392
rect 3421 22383 3479 22389
rect 5350 22380 5356 22392
rect 5408 22380 5414 22432
rect 6457 22423 6515 22429
rect 6457 22389 6469 22423
rect 6503 22420 6515 22423
rect 11330 22420 11336 22432
rect 6503 22392 11336 22420
rect 6503 22389 6515 22392
rect 6457 22383 6515 22389
rect 11330 22380 11336 22392
rect 11388 22380 11394 22432
rect 11882 22380 11888 22432
rect 11940 22380 11946 22432
rect 13446 22380 13452 22432
rect 13504 22420 13510 22432
rect 14185 22423 14243 22429
rect 14185 22420 14197 22423
rect 13504 22392 14197 22420
rect 13504 22380 13510 22392
rect 14185 22389 14197 22392
rect 14231 22389 14243 22423
rect 14185 22383 14243 22389
rect 19061 22423 19119 22429
rect 19061 22389 19073 22423
rect 19107 22420 19119 22423
rect 19150 22420 19156 22432
rect 19107 22392 19156 22420
rect 19107 22389 19119 22392
rect 19061 22383 19119 22389
rect 19150 22380 19156 22392
rect 19208 22380 19214 22432
rect 20162 22380 20168 22432
rect 20220 22420 20226 22432
rect 20346 22420 20352 22432
rect 20220 22392 20352 22420
rect 20220 22380 20226 22392
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 20714 22380 20720 22432
rect 20772 22420 20778 22432
rect 23566 22420 23572 22432
rect 20772 22392 23572 22420
rect 20772 22380 20778 22392
rect 23566 22380 23572 22392
rect 23624 22380 23630 22432
rect 23934 22380 23940 22432
rect 23992 22420 23998 22432
rect 24872 22429 24900 22460
rect 26050 22448 26056 22500
rect 26108 22488 26114 22500
rect 27157 22491 27215 22497
rect 27157 22488 27169 22491
rect 26108 22460 27169 22488
rect 26108 22448 26114 22460
rect 27157 22457 27169 22460
rect 27203 22457 27215 22491
rect 27157 22451 27215 22457
rect 27522 22448 27528 22500
rect 27580 22488 27586 22500
rect 27724 22488 27752 22519
rect 28350 22516 28356 22568
rect 28408 22516 28414 22568
rect 28994 22516 29000 22568
rect 29052 22556 29058 22568
rect 30101 22559 30159 22565
rect 30101 22556 30113 22559
rect 29052 22528 30113 22556
rect 29052 22516 29058 22528
rect 30101 22525 30113 22528
rect 30147 22525 30159 22559
rect 30208 22556 30236 22596
rect 30929 22593 30941 22627
rect 30975 22624 30987 22627
rect 31018 22624 31024 22636
rect 30975 22596 31024 22624
rect 30975 22593 30987 22596
rect 30929 22587 30987 22593
rect 31018 22584 31024 22596
rect 31076 22584 31082 22636
rect 31754 22584 31760 22636
rect 31812 22624 31818 22636
rect 31849 22627 31907 22633
rect 31849 22624 31861 22627
rect 31812 22596 31861 22624
rect 31812 22584 31818 22596
rect 31849 22593 31861 22596
rect 31895 22624 31907 22627
rect 32214 22624 32220 22636
rect 31895 22596 32220 22624
rect 31895 22593 31907 22596
rect 31849 22587 31907 22593
rect 32214 22584 32220 22596
rect 32272 22584 32278 22636
rect 32401 22627 32459 22633
rect 32401 22593 32413 22627
rect 32447 22624 32459 22627
rect 32490 22624 32496 22636
rect 32447 22596 32496 22624
rect 32447 22593 32459 22596
rect 32401 22587 32459 22593
rect 32490 22584 32496 22596
rect 32548 22584 32554 22636
rect 33137 22627 33195 22633
rect 33137 22593 33149 22627
rect 33183 22624 33195 22627
rect 33410 22624 33416 22636
rect 33183 22596 33416 22624
rect 33183 22593 33195 22596
rect 33137 22587 33195 22593
rect 33410 22584 33416 22596
rect 33468 22584 33474 22636
rect 34238 22584 34244 22636
rect 34296 22584 34302 22636
rect 34514 22584 34520 22636
rect 34572 22584 34578 22636
rect 34698 22584 34704 22636
rect 34756 22624 34762 22636
rect 35621 22627 35679 22633
rect 35621 22624 35633 22627
rect 34756 22596 35633 22624
rect 34756 22584 34762 22596
rect 35621 22593 35633 22596
rect 35667 22593 35679 22627
rect 35621 22587 35679 22593
rect 35710 22584 35716 22636
rect 35768 22624 35774 22636
rect 36357 22627 36415 22633
rect 36357 22624 36369 22627
rect 35768 22596 36369 22624
rect 35768 22584 35774 22596
rect 36357 22593 36369 22596
rect 36403 22593 36415 22627
rect 36357 22587 36415 22593
rect 37369 22627 37427 22633
rect 37369 22593 37381 22627
rect 37415 22624 37427 22627
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37415 22596 37841 22624
rect 37415 22593 37427 22596
rect 37369 22587 37427 22593
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 40865 22627 40923 22633
rect 40865 22593 40877 22627
rect 40911 22624 40923 22627
rect 41414 22624 41420 22636
rect 40911 22596 41420 22624
rect 40911 22593 40923 22596
rect 40865 22587 40923 22593
rect 31113 22559 31171 22565
rect 31113 22556 31125 22559
rect 30208 22528 31125 22556
rect 30101 22519 30159 22525
rect 31113 22525 31125 22528
rect 31159 22525 31171 22559
rect 33597 22559 33655 22565
rect 33597 22556 33609 22559
rect 31113 22519 31171 22525
rect 31220 22528 33609 22556
rect 27580 22460 27752 22488
rect 27580 22448 27586 22460
rect 29638 22448 29644 22500
rect 29696 22488 29702 22500
rect 29696 22460 30512 22488
rect 29696 22448 29702 22460
rect 24857 22423 24915 22429
rect 24857 22420 24869 22423
rect 23992 22392 24869 22420
rect 23992 22380 23998 22392
rect 24857 22389 24869 22392
rect 24903 22389 24915 22423
rect 24857 22383 24915 22389
rect 25314 22380 25320 22432
rect 25372 22380 25378 22432
rect 25682 22380 25688 22432
rect 25740 22420 25746 22432
rect 28258 22420 28264 22432
rect 25740 22392 28264 22420
rect 25740 22380 25746 22392
rect 28258 22380 28264 22392
rect 28316 22380 28322 22432
rect 28350 22380 28356 22432
rect 28408 22420 28414 22432
rect 29822 22420 29828 22432
rect 28408 22392 29828 22420
rect 28408 22380 28414 22392
rect 29822 22380 29828 22392
rect 29880 22380 29886 22432
rect 30484 22420 30512 22460
rect 30558 22448 30564 22500
rect 30616 22448 30622 22500
rect 31220 22420 31248 22528
rect 33597 22525 33609 22528
rect 33643 22525 33655 22559
rect 33597 22519 33655 22525
rect 31665 22491 31723 22497
rect 31665 22457 31677 22491
rect 31711 22488 31723 22491
rect 31846 22488 31852 22500
rect 31711 22460 31852 22488
rect 31711 22457 31723 22460
rect 31665 22451 31723 22457
rect 31846 22448 31852 22460
rect 31904 22488 31910 22500
rect 32030 22488 32036 22500
rect 31904 22460 32036 22488
rect 31904 22448 31910 22460
rect 32030 22448 32036 22460
rect 32088 22488 32094 22500
rect 37384 22488 37412 22587
rect 41414 22584 41420 22596
rect 41472 22584 41478 22636
rect 41524 22633 41552 22664
rect 41785 22661 41797 22664
rect 41831 22661 41843 22695
rect 41785 22655 41843 22661
rect 47673 22695 47731 22701
rect 47673 22661 47685 22695
rect 47719 22692 47731 22695
rect 47719 22664 49096 22692
rect 47719 22661 47731 22664
rect 47673 22655 47731 22661
rect 49068 22636 49096 22664
rect 41509 22627 41567 22633
rect 41509 22593 41521 22627
rect 41555 22593 41567 22627
rect 41509 22587 41567 22593
rect 42613 22627 42671 22633
rect 42613 22593 42625 22627
rect 42659 22624 42671 22627
rect 42794 22624 42800 22636
rect 42659 22596 42800 22624
rect 42659 22593 42671 22596
rect 42613 22587 42671 22593
rect 42794 22584 42800 22596
rect 42852 22584 42858 22636
rect 43901 22627 43959 22633
rect 43901 22593 43913 22627
rect 43947 22624 43959 22627
rect 46842 22624 46848 22636
rect 43947 22596 46848 22624
rect 43947 22593 43959 22596
rect 43901 22587 43959 22593
rect 46842 22584 46848 22596
rect 46900 22584 46906 22636
rect 48041 22627 48099 22633
rect 48041 22593 48053 22627
rect 48087 22624 48099 22627
rect 48314 22624 48320 22636
rect 48087 22596 48320 22624
rect 48087 22593 48099 22596
rect 48041 22587 48099 22593
rect 48314 22584 48320 22596
rect 48372 22584 48378 22636
rect 49050 22584 49056 22636
rect 49108 22584 49114 22636
rect 38105 22559 38163 22565
rect 38105 22525 38117 22559
rect 38151 22556 38163 22559
rect 44545 22559 44603 22565
rect 44545 22556 44557 22559
rect 38151 22528 44557 22556
rect 38151 22525 38163 22528
rect 38105 22519 38163 22525
rect 44545 22525 44557 22528
rect 44591 22525 44603 22559
rect 44545 22519 44603 22525
rect 32088 22460 37412 22488
rect 32088 22448 32094 22460
rect 30484 22392 31248 22420
rect 32122 22380 32128 22432
rect 32180 22420 32186 22432
rect 32493 22423 32551 22429
rect 32493 22420 32505 22423
rect 32180 22392 32505 22420
rect 32180 22380 32186 22392
rect 32493 22389 32505 22392
rect 32539 22389 32551 22423
rect 32493 22383 32551 22389
rect 34514 22380 34520 22432
rect 34572 22420 34578 22432
rect 35713 22423 35771 22429
rect 35713 22420 35725 22423
rect 34572 22392 35725 22420
rect 34572 22380 34578 22392
rect 35713 22389 35725 22392
rect 35759 22389 35771 22423
rect 35713 22383 35771 22389
rect 39574 22380 39580 22432
rect 39632 22380 39638 22432
rect 40678 22380 40684 22432
rect 40736 22380 40742 22432
rect 41322 22380 41328 22432
rect 41380 22380 41386 22432
rect 48498 22380 48504 22432
rect 48556 22380 48562 22432
rect 49234 22380 49240 22432
rect 49292 22380 49298 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 3694 22216 3700 22228
rect 2280 22188 3700 22216
rect 2280 22176 2286 22188
rect 3694 22176 3700 22188
rect 3752 22176 3758 22228
rect 11882 22216 11888 22228
rect 5552 22188 11888 22216
rect 3418 22108 3424 22160
rect 3476 22148 3482 22160
rect 4154 22148 4160 22160
rect 3476 22120 4160 22148
rect 3476 22108 3482 22120
rect 4154 22108 4160 22120
rect 4212 22108 4218 22160
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 4062 22040 4068 22092
rect 4120 22080 4126 22092
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 4120 22052 4445 22080
rect 4120 22040 4126 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4433 22043 4491 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 3605 22015 3663 22021
rect 1811 21984 2774 22012
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 2746 21944 2774 21984
rect 3605 21981 3617 22015
rect 3651 22012 3663 22015
rect 3786 22012 3792 22024
rect 3651 21984 3792 22012
rect 3651 21981 3663 21984
rect 3605 21975 3663 21981
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 22012 4031 22015
rect 4246 22012 4252 22024
rect 4019 21984 4252 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 5552 21944 5580 22188
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 11974 22176 11980 22228
rect 12032 22216 12038 22228
rect 14461 22219 14519 22225
rect 14461 22216 14473 22219
rect 12032 22188 14473 22216
rect 12032 22176 12038 22188
rect 14461 22185 14473 22188
rect 14507 22185 14519 22219
rect 14461 22179 14519 22185
rect 14550 22176 14556 22228
rect 14608 22176 14614 22228
rect 16390 22176 16396 22228
rect 16448 22216 16454 22228
rect 23382 22216 23388 22228
rect 16448 22188 23388 22216
rect 16448 22176 16454 22188
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 26050 22216 26056 22228
rect 23768 22188 26056 22216
rect 6730 22108 6736 22160
rect 6788 22148 6794 22160
rect 6788 22120 7328 22148
rect 6788 22108 6794 22120
rect 7300 22089 7328 22120
rect 9030 22108 9036 22160
rect 9088 22108 9094 22160
rect 11054 22148 11060 22160
rect 9784 22120 11060 22148
rect 9784 22089 9812 22120
rect 11054 22108 11060 22120
rect 11112 22108 11118 22160
rect 11330 22108 11336 22160
rect 11388 22148 11394 22160
rect 14568 22148 14596 22176
rect 11388 22120 14596 22148
rect 11388 22108 11394 22120
rect 18506 22108 18512 22160
rect 18564 22148 18570 22160
rect 19058 22148 19064 22160
rect 18564 22120 19064 22148
rect 18564 22108 18570 22120
rect 19058 22108 19064 22120
rect 19116 22108 19122 22160
rect 20073 22151 20131 22157
rect 20073 22117 20085 22151
rect 20119 22148 20131 22151
rect 21726 22148 21732 22160
rect 20119 22120 21732 22148
rect 20119 22117 20131 22120
rect 20073 22111 20131 22117
rect 21726 22108 21732 22120
rect 21784 22108 21790 22160
rect 21818 22108 21824 22160
rect 21876 22148 21882 22160
rect 22278 22148 22284 22160
rect 21876 22120 22284 22148
rect 21876 22108 21882 22120
rect 22278 22108 22284 22120
rect 22336 22108 22342 22160
rect 7285 22083 7343 22089
rect 2746 21916 5580 21944
rect 5644 22052 7052 22080
rect 3421 21879 3479 21885
rect 3421 21845 3433 21879
rect 3467 21876 3479 21879
rect 5644 21876 5672 22052
rect 6273 22015 6331 22021
rect 6273 21981 6285 22015
rect 6319 22012 6331 22015
rect 6638 22012 6644 22024
rect 6319 21984 6644 22012
rect 6319 21981 6331 21984
rect 6273 21975 6331 21981
rect 6638 21972 6644 21984
rect 6696 21972 6702 22024
rect 6914 21972 6920 22024
rect 6972 21972 6978 22024
rect 7024 22012 7052 22052
rect 7285 22049 7297 22083
rect 7331 22049 7343 22083
rect 9769 22083 9827 22089
rect 7285 22043 7343 22049
rect 8680 22052 9076 22080
rect 8386 22012 8392 22024
rect 7024 21984 8392 22012
rect 8386 21972 8392 21984
rect 8444 21972 8450 22024
rect 8680 22012 8708 22052
rect 8496 21984 8708 22012
rect 5813 21947 5871 21953
rect 5813 21913 5825 21947
rect 5859 21944 5871 21947
rect 8496 21944 8524 21984
rect 8754 21972 8760 22024
rect 8812 21972 8818 22024
rect 9048 22012 9076 22052
rect 9769 22049 9781 22083
rect 9815 22080 9827 22083
rect 9953 22083 10011 22089
rect 9815 22052 9849 22080
rect 9815 22049 9827 22052
rect 9769 22043 9827 22049
rect 9953 22049 9965 22083
rect 9999 22080 10011 22083
rect 10042 22080 10048 22092
rect 9999 22052 10048 22080
rect 9999 22049 10011 22052
rect 9953 22043 10011 22049
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 11238 22040 11244 22092
rect 11296 22040 11302 22092
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 15102 22040 15108 22092
rect 15160 22080 15166 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 15160 22052 15669 22080
rect 15160 22040 15166 22052
rect 15657 22049 15669 22052
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 17129 22083 17187 22089
rect 17129 22049 17141 22083
rect 17175 22080 17187 22083
rect 19426 22080 19432 22092
rect 17175 22052 19432 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 22649 22083 22707 22089
rect 22649 22049 22661 22083
rect 22695 22080 22707 22083
rect 23566 22080 23572 22092
rect 22695 22052 23572 22080
rect 22695 22049 22707 22052
rect 22649 22043 22707 22049
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 23768 22089 23796 22188
rect 26050 22176 26056 22188
rect 26108 22176 26114 22228
rect 26234 22176 26240 22228
rect 26292 22216 26298 22228
rect 27522 22216 27528 22228
rect 26292 22188 27528 22216
rect 26292 22176 26298 22188
rect 27522 22176 27528 22188
rect 27580 22176 27586 22228
rect 28629 22219 28687 22225
rect 28629 22216 28641 22219
rect 27632 22188 28641 22216
rect 24302 22108 24308 22160
rect 24360 22148 24366 22160
rect 24581 22151 24639 22157
rect 24581 22148 24593 22151
rect 24360 22120 24593 22148
rect 24360 22108 24366 22120
rect 24581 22117 24593 22120
rect 24627 22117 24639 22151
rect 24581 22111 24639 22117
rect 25240 22120 25912 22148
rect 23753 22083 23811 22089
rect 23753 22049 23765 22083
rect 23799 22049 23811 22083
rect 23753 22043 23811 22049
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 24762 22080 24768 22092
rect 23983 22052 24768 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 24762 22040 24768 22052
rect 24820 22040 24826 22092
rect 25240 22089 25268 22120
rect 25225 22083 25283 22089
rect 25225 22049 25237 22083
rect 25271 22080 25283 22083
rect 25884 22080 25912 22120
rect 27246 22108 27252 22160
rect 27304 22148 27310 22160
rect 27632 22148 27660 22188
rect 28629 22185 28641 22188
rect 28675 22185 28687 22219
rect 28629 22179 28687 22185
rect 29641 22219 29699 22225
rect 29641 22185 29653 22219
rect 29687 22216 29699 22219
rect 29822 22216 29828 22228
rect 29687 22188 29828 22216
rect 29687 22185 29699 22188
rect 29641 22179 29699 22185
rect 29822 22176 29828 22188
rect 29880 22176 29886 22228
rect 31938 22216 31944 22228
rect 29932 22188 31944 22216
rect 27304 22120 27660 22148
rect 27304 22108 27310 22120
rect 28258 22108 28264 22160
rect 28316 22148 28322 22160
rect 29932 22148 29960 22188
rect 31938 22176 31944 22188
rect 31996 22176 32002 22228
rect 35434 22216 35440 22228
rect 32048 22188 35440 22216
rect 28316 22120 29960 22148
rect 30668 22120 30880 22148
rect 28316 22108 28322 22120
rect 26050 22080 26056 22092
rect 25271 22052 25305 22080
rect 25884 22052 26056 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 26050 22040 26056 22052
rect 26108 22040 26114 22092
rect 28442 22040 28448 22092
rect 28500 22080 28506 22092
rect 28500 22052 28994 22080
rect 28500 22040 28506 22052
rect 10410 22012 10416 22024
rect 9048 21984 10416 22012
rect 10410 21972 10416 21984
rect 10468 21972 10474 22024
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 14369 22015 14427 22021
rect 12575 21984 12609 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 14369 21981 14381 22015
rect 14415 22012 14427 22015
rect 14550 22012 14556 22024
rect 14415 21984 14556 22012
rect 14415 21981 14427 21984
rect 14369 21975 14427 21981
rect 5859 21916 8524 21944
rect 8573 21947 8631 21953
rect 5859 21913 5871 21916
rect 5813 21907 5871 21913
rect 8573 21913 8585 21947
rect 8619 21944 8631 21947
rect 12544 21944 12572 21975
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 15194 21972 15200 22024
rect 15252 22012 15258 22024
rect 15378 22012 15384 22024
rect 15252 21984 15384 22012
rect 15252 21972 15258 21984
rect 15378 21972 15384 21984
rect 15436 21972 15442 22024
rect 18506 21972 18512 22024
rect 18564 21972 18570 22024
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 18932 21984 20208 22012
rect 18932 21972 18938 21984
rect 12710 21944 12716 21956
rect 8619 21916 12716 21944
rect 8619 21913 8631 21916
rect 8573 21907 8631 21913
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 17405 21947 17463 21953
rect 17405 21913 17417 21947
rect 17451 21944 17463 21947
rect 17494 21944 17500 21956
rect 17451 21916 17500 21944
rect 17451 21913 17463 21916
rect 17405 21907 17463 21913
rect 17494 21904 17500 21916
rect 17552 21904 17558 21956
rect 19521 21947 19579 21953
rect 19521 21944 19533 21947
rect 18708 21916 19533 21944
rect 3467 21848 5672 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 6086 21836 6092 21888
rect 6144 21836 6150 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9677 21879 9735 21885
rect 9677 21845 9689 21879
rect 9723 21876 9735 21879
rect 9950 21876 9956 21888
rect 9723 21848 9956 21876
rect 9723 21845 9735 21848
rect 9677 21839 9735 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 10502 21836 10508 21888
rect 10560 21876 10566 21888
rect 10778 21876 10784 21888
rect 10560 21848 10784 21876
rect 10560 21836 10566 21848
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 11514 21836 11520 21888
rect 11572 21876 11578 21888
rect 14642 21876 14648 21888
rect 11572 21848 14648 21876
rect 11572 21836 11578 21848
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 14918 21836 14924 21888
rect 14976 21876 14982 21888
rect 18708 21876 18736 21916
rect 19521 21913 19533 21916
rect 19567 21913 19579 21947
rect 19521 21907 19579 21913
rect 14976 21848 18736 21876
rect 14976 21836 14982 21848
rect 18782 21836 18788 21888
rect 18840 21876 18846 21888
rect 18877 21879 18935 21885
rect 18877 21876 18889 21879
rect 18840 21848 18889 21876
rect 18840 21836 18846 21848
rect 18877 21845 18889 21848
rect 18923 21845 18935 21879
rect 18877 21839 18935 21845
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 19613 21879 19671 21885
rect 19613 21876 19625 21879
rect 19392 21848 19625 21876
rect 19392 21836 19398 21848
rect 19613 21845 19625 21848
rect 19659 21845 19671 21879
rect 20180 21876 20208 21984
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 24670 22012 24676 22024
rect 22848 21984 24676 22012
rect 20254 21904 20260 21956
rect 20312 21944 20318 21956
rect 21269 21947 21327 21953
rect 21269 21944 21281 21947
rect 20312 21916 21281 21944
rect 20312 21904 20318 21916
rect 21269 21913 21281 21916
rect 21315 21913 21327 21947
rect 22848 21944 22876 21984
rect 24670 21972 24676 21984
rect 24728 21972 24734 22024
rect 25774 21972 25780 22024
rect 25832 21972 25838 22024
rect 28626 21972 28632 22024
rect 28684 22008 28690 22024
rect 28789 22011 28847 22017
rect 28789 22008 28801 22011
rect 28684 21980 28801 22008
rect 28684 21972 28690 21980
rect 28789 21977 28801 21980
rect 28835 21977 28847 22011
rect 28966 22012 28994 22052
rect 29178 22040 29184 22092
rect 29236 22040 29242 22092
rect 30668 22080 30696 22120
rect 30484 22052 30696 22080
rect 29273 22015 29331 22021
rect 28966 22008 29040 22012
rect 29273 22008 29285 22015
rect 28966 21984 29285 22008
rect 29012 21981 29285 21984
rect 29319 21981 29331 22015
rect 29012 21980 29331 21981
rect 28789 21971 28847 21977
rect 29273 21975 29331 21980
rect 29546 21972 29552 22024
rect 29604 22012 29610 22024
rect 30484 22012 30512 22052
rect 30742 22040 30748 22092
rect 30800 22040 30806 22092
rect 30852 22080 30880 22120
rect 31202 22108 31208 22160
rect 31260 22148 31266 22160
rect 32048 22148 32076 22188
rect 35434 22176 35440 22188
rect 35492 22176 35498 22228
rect 42794 22176 42800 22228
rect 42852 22216 42858 22228
rect 49234 22216 49240 22228
rect 42852 22188 49240 22216
rect 42852 22176 42858 22188
rect 49234 22176 49240 22188
rect 49292 22176 49298 22228
rect 31260 22120 32076 22148
rect 31260 22108 31266 22120
rect 32122 22108 32128 22160
rect 32180 22148 32186 22160
rect 32582 22148 32588 22160
rect 32180 22120 32588 22148
rect 32180 22108 32186 22120
rect 32582 22108 32588 22120
rect 32640 22108 32646 22160
rect 32674 22108 32680 22160
rect 32732 22108 32738 22160
rect 37642 22108 37648 22160
rect 37700 22148 37706 22160
rect 37700 22120 38976 22148
rect 37700 22108 37706 22120
rect 31849 22083 31907 22089
rect 31849 22080 31861 22083
rect 30852 22052 31861 22080
rect 31849 22049 31861 22052
rect 31895 22049 31907 22083
rect 31849 22043 31907 22049
rect 32030 22040 32036 22092
rect 32088 22040 32094 22092
rect 32214 22040 32220 22092
rect 32272 22080 32278 22092
rect 32692 22080 32720 22108
rect 38746 22080 38752 22092
rect 32272 22052 32720 22080
rect 33244 22052 38752 22080
rect 32272 22040 32278 22052
rect 29604 21984 30512 22012
rect 30561 22015 30619 22021
rect 29604 21972 29610 21984
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 30607 21984 31892 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 21269 21907 21327 21913
rect 22020 21916 22876 21944
rect 22020 21876 22048 21916
rect 22922 21904 22928 21956
rect 22980 21944 22986 21956
rect 22980 21916 23612 21944
rect 22980 21904 22986 21916
rect 20180 21848 22048 21876
rect 22097 21879 22155 21885
rect 19613 21839 19671 21845
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22186 21876 22192 21888
rect 22143 21848 22192 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 23290 21836 23296 21888
rect 23348 21836 23354 21888
rect 23584 21876 23612 21916
rect 24946 21904 24952 21956
rect 25004 21904 25010 21956
rect 26050 21904 26056 21956
rect 26108 21904 26114 21956
rect 26510 21904 26516 21956
rect 26568 21904 26574 21956
rect 28902 21904 28908 21956
rect 28960 21944 28966 21956
rect 28960 21916 29500 21944
rect 28960 21904 28966 21916
rect 23661 21879 23719 21885
rect 23661 21876 23673 21879
rect 23584 21848 23673 21876
rect 23661 21845 23673 21848
rect 23707 21845 23719 21879
rect 23661 21839 23719 21845
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 25682 21876 25688 21888
rect 25087 21848 25688 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 25682 21836 25688 21848
rect 25740 21836 25746 21888
rect 25958 21836 25964 21888
rect 26016 21876 26022 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 26016 21848 27997 21876
rect 26016 21836 26022 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 27985 21839 28043 21845
rect 28718 21836 28724 21888
rect 28776 21876 28782 21888
rect 29362 21876 29368 21888
rect 28776 21848 29368 21876
rect 28776 21836 28782 21848
rect 29362 21836 29368 21848
rect 29420 21836 29426 21888
rect 29472 21876 29500 21916
rect 29638 21904 29644 21956
rect 29696 21944 29702 21956
rect 29696 21916 30604 21944
rect 29696 21904 29702 21916
rect 30101 21879 30159 21885
rect 30101 21876 30113 21879
rect 29472 21848 30113 21876
rect 30101 21845 30113 21848
rect 30147 21845 30159 21879
rect 30101 21839 30159 21845
rect 30374 21836 30380 21888
rect 30432 21876 30438 21888
rect 30469 21879 30527 21885
rect 30469 21876 30481 21879
rect 30432 21848 30481 21876
rect 30432 21836 30438 21848
rect 30469 21845 30481 21848
rect 30515 21845 30527 21879
rect 30576 21876 30604 21916
rect 31386 21904 31392 21956
rect 31444 21904 31450 21956
rect 31481 21879 31539 21885
rect 31481 21876 31493 21879
rect 30576 21848 31493 21876
rect 30469 21839 30527 21845
rect 31481 21845 31493 21848
rect 31527 21845 31539 21879
rect 31864 21876 31892 21984
rect 32030 21904 32036 21956
rect 32088 21944 32094 21956
rect 32232 21944 32260 22040
rect 32582 21972 32588 22024
rect 32640 21972 32646 22024
rect 32858 21972 32864 22024
rect 32916 21972 32922 22024
rect 32088 21916 32260 21944
rect 32088 21904 32094 21916
rect 33244 21876 33272 22052
rect 38746 22040 38752 22052
rect 38804 22040 38810 22092
rect 38948 22080 38976 22120
rect 48406 22108 48412 22160
rect 48464 22108 48470 22160
rect 39209 22083 39267 22089
rect 39209 22080 39221 22083
rect 38948 22052 39221 22080
rect 33965 22015 34023 22021
rect 33965 21981 33977 22015
rect 34011 22012 34023 22015
rect 34054 22012 34060 22024
rect 34011 21984 34060 22012
rect 34011 21981 34023 21984
rect 33965 21975 34023 21981
rect 34054 21972 34060 21984
rect 34112 21972 34118 22024
rect 34517 22015 34575 22021
rect 34517 21981 34529 22015
rect 34563 22012 34575 22015
rect 35158 22012 35164 22024
rect 34563 21984 35164 22012
rect 34563 21981 34575 21984
rect 34517 21975 34575 21981
rect 35158 21972 35164 21984
rect 35216 21972 35222 22024
rect 35434 21972 35440 22024
rect 35492 22012 35498 22024
rect 35805 22015 35863 22021
rect 35805 22012 35817 22015
rect 35492 21984 35817 22012
rect 35492 21972 35498 21984
rect 35805 21981 35817 21984
rect 35851 21981 35863 22015
rect 35805 21975 35863 21981
rect 37274 21972 37280 22024
rect 37332 22012 37338 22024
rect 38948 22021 38976 22052
rect 39209 22049 39221 22052
rect 39255 22049 39267 22083
rect 39209 22043 39267 22049
rect 37645 22015 37703 22021
rect 37645 22012 37657 22015
rect 37332 21984 37657 22012
rect 37332 21972 37338 21984
rect 37645 21981 37657 21984
rect 37691 22012 37703 22015
rect 37921 22015 37979 22021
rect 37921 22012 37933 22015
rect 37691 21984 37933 22012
rect 37691 21981 37703 21984
rect 37645 21975 37703 21981
rect 37921 21981 37933 21984
rect 37967 21981 37979 22015
rect 37921 21975 37979 21981
rect 38933 22015 38991 22021
rect 38933 21981 38945 22015
rect 38979 21981 38991 22015
rect 38933 21975 38991 21981
rect 48593 22015 48651 22021
rect 48593 21981 48605 22015
rect 48639 22012 48651 22015
rect 48682 22012 48688 22024
rect 48639 21984 48688 22012
rect 48639 21981 48651 21984
rect 48593 21975 48651 21981
rect 48682 21972 48688 21984
rect 48740 21972 48746 22024
rect 49050 21972 49056 22024
rect 49108 21972 49114 22024
rect 34974 21904 34980 21956
rect 35032 21904 35038 21956
rect 36446 21904 36452 21956
rect 36504 21944 36510 21956
rect 40310 21944 40316 21956
rect 36504 21916 40316 21944
rect 36504 21904 36510 21916
rect 40310 21904 40316 21916
rect 40368 21904 40374 21956
rect 31864 21848 33272 21876
rect 31481 21839 31539 21845
rect 33594 21836 33600 21888
rect 33652 21876 33658 21888
rect 34057 21879 34115 21885
rect 34057 21876 34069 21879
rect 33652 21848 34069 21876
rect 33652 21836 33658 21848
rect 34057 21845 34069 21848
rect 34103 21845 34115 21879
rect 34057 21839 34115 21845
rect 35066 21836 35072 21888
rect 35124 21836 35130 21888
rect 35618 21836 35624 21888
rect 35676 21836 35682 21888
rect 36262 21836 36268 21888
rect 36320 21836 36326 21888
rect 37458 21836 37464 21888
rect 37516 21836 37522 21888
rect 37550 21836 37556 21888
rect 37608 21876 37614 21888
rect 38749 21879 38807 21885
rect 38749 21876 38761 21879
rect 37608 21848 38761 21876
rect 37608 21836 37614 21848
rect 38749 21845 38761 21848
rect 38795 21845 38807 21879
rect 38749 21839 38807 21845
rect 49234 21836 49240 21888
rect 49292 21836 49298 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 3418 21632 3424 21684
rect 3476 21672 3482 21684
rect 3602 21672 3608 21684
rect 3476 21644 3608 21672
rect 3476 21632 3482 21644
rect 3602 21632 3608 21644
rect 3660 21632 3666 21684
rect 4246 21632 4252 21684
rect 4304 21672 4310 21684
rect 9214 21672 9220 21684
rect 4304 21644 9220 21672
rect 4304 21632 4310 21644
rect 9214 21632 9220 21644
rect 9272 21632 9278 21684
rect 9398 21632 9404 21684
rect 9456 21632 9462 21684
rect 10321 21675 10379 21681
rect 10321 21641 10333 21675
rect 10367 21672 10379 21675
rect 10686 21672 10692 21684
rect 10367 21644 10692 21672
rect 10367 21641 10379 21644
rect 10321 21635 10379 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 10962 21632 10968 21684
rect 11020 21632 11026 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 15930 21672 15936 21684
rect 11195 21644 15936 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 16022 21632 16028 21684
rect 16080 21632 16086 21684
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 16264 21644 20300 21672
rect 16264 21632 16270 21644
rect 5810 21604 5816 21616
rect 1596 21576 5816 21604
rect 1596 21545 1624 21576
rect 5810 21564 5816 21576
rect 5868 21564 5874 21616
rect 6270 21564 6276 21616
rect 6328 21604 6334 21616
rect 7558 21604 7564 21616
rect 6328 21576 7564 21604
rect 6328 21564 6334 21576
rect 7558 21564 7564 21576
rect 7616 21604 7622 21616
rect 7929 21607 7987 21613
rect 7929 21604 7941 21607
rect 7616 21576 7941 21604
rect 7616 21564 7622 21576
rect 7929 21573 7941 21576
rect 7975 21573 7987 21607
rect 9416 21604 9444 21632
rect 9416 21576 12480 21604
rect 7929 21567 7987 21573
rect 1581 21539 1639 21545
rect 1581 21505 1593 21539
rect 1627 21505 1639 21539
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 1581 21499 1639 21505
rect 1688 21508 3433 21536
rect 1118 21428 1124 21480
rect 1176 21468 1182 21480
rect 1688 21468 1716 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21536 7067 21539
rect 7098 21536 7104 21548
rect 7055 21508 7104 21536
rect 7055 21505 7067 21508
rect 7009 21499 7067 21505
rect 7098 21496 7104 21508
rect 7156 21496 7162 21548
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7576 21508 7665 21536
rect 1176 21440 1716 21468
rect 1176 21428 1182 21440
rect 1946 21428 1952 21480
rect 2004 21468 2010 21480
rect 2041 21471 2099 21477
rect 2041 21468 2053 21471
rect 2004 21440 2053 21468
rect 2004 21428 2010 21440
rect 2041 21437 2053 21440
rect 2087 21437 2099 21471
rect 2041 21431 2099 21437
rect 4154 21428 4160 21480
rect 4212 21428 4218 21480
rect 5534 21428 5540 21480
rect 5592 21468 5598 21480
rect 5721 21471 5779 21477
rect 5721 21468 5733 21471
rect 5592 21440 5733 21468
rect 5592 21428 5598 21440
rect 5721 21437 5733 21440
rect 5767 21437 5779 21471
rect 5721 21431 5779 21437
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6454 21468 6460 21480
rect 5951 21440 6460 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 6454 21428 6460 21440
rect 6512 21428 6518 21480
rect 6178 21360 6184 21412
rect 6236 21400 6242 21412
rect 6549 21403 6607 21409
rect 6549 21400 6561 21403
rect 6236 21372 6561 21400
rect 6236 21360 6242 21372
rect 6549 21369 6561 21372
rect 6595 21369 6607 21403
rect 6549 21363 6607 21369
rect 3326 21292 3332 21344
rect 3384 21332 3390 21344
rect 3602 21332 3608 21344
rect 3384 21304 3608 21332
rect 3384 21292 3390 21304
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 5261 21335 5319 21341
rect 5261 21301 5273 21335
rect 5307 21332 5319 21335
rect 5534 21332 5540 21344
rect 5307 21304 5540 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 6454 21292 6460 21344
rect 6512 21292 6518 21344
rect 7098 21292 7104 21344
rect 7156 21292 7162 21344
rect 7576 21332 7604 21508
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 9030 21496 9036 21548
rect 9088 21536 9094 21548
rect 10134 21536 10140 21548
rect 9088 21508 10140 21536
rect 9088 21496 9094 21508
rect 10134 21496 10140 21508
rect 10192 21496 10198 21548
rect 10229 21539 10287 21545
rect 10229 21505 10241 21539
rect 10275 21505 10287 21539
rect 10229 21499 10287 21505
rect 7926 21428 7932 21480
rect 7984 21468 7990 21480
rect 10244 21468 10272 21499
rect 10318 21496 10324 21548
rect 10376 21536 10382 21548
rect 12161 21539 12219 21545
rect 12161 21536 12173 21539
rect 10376 21508 12173 21536
rect 10376 21496 10382 21508
rect 12161 21505 12173 21508
rect 12207 21505 12219 21539
rect 12161 21499 12219 21505
rect 7984 21440 10272 21468
rect 10505 21471 10563 21477
rect 7984 21428 7990 21440
rect 10505 21437 10517 21471
rect 10551 21468 10563 21471
rect 10870 21468 10876 21480
rect 10551 21440 10876 21468
rect 10551 21437 10563 21440
rect 10505 21431 10563 21437
rect 10870 21428 10876 21440
rect 10928 21428 10934 21480
rect 12452 21477 12480 21576
rect 12710 21564 12716 21616
rect 12768 21604 12774 21616
rect 13357 21607 13415 21613
rect 13357 21604 13369 21607
rect 12768 21576 13369 21604
rect 12768 21564 12774 21576
rect 13357 21573 13369 21576
rect 13403 21604 13415 21607
rect 13446 21604 13452 21616
rect 13403 21576 13452 21604
rect 13403 21573 13415 21576
rect 13357 21567 13415 21573
rect 13446 21564 13452 21576
rect 13504 21564 13510 21616
rect 13814 21564 13820 21616
rect 13872 21564 13878 21616
rect 14642 21564 14648 21616
rect 14700 21604 14706 21616
rect 20272 21604 20300 21644
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 20993 21675 21051 21681
rect 20993 21672 21005 21675
rect 20864 21644 21005 21672
rect 20864 21632 20870 21644
rect 20993 21641 21005 21644
rect 21039 21672 21051 21675
rect 21634 21672 21640 21684
rect 21039 21644 21640 21672
rect 21039 21641 21051 21644
rect 20993 21635 21051 21641
rect 21634 21632 21640 21644
rect 21692 21632 21698 21684
rect 21726 21632 21732 21684
rect 21784 21672 21790 21684
rect 23017 21675 23075 21681
rect 23017 21672 23029 21675
rect 21784 21644 23029 21672
rect 21784 21632 21790 21644
rect 23017 21641 23029 21644
rect 23063 21672 23075 21675
rect 23382 21672 23388 21684
rect 23063 21644 23388 21672
rect 23063 21641 23075 21644
rect 23017 21635 23075 21641
rect 23382 21632 23388 21644
rect 23440 21672 23446 21684
rect 24394 21672 24400 21684
rect 23440 21644 24400 21672
rect 23440 21632 23446 21644
rect 24394 21632 24400 21644
rect 24452 21632 24458 21684
rect 25958 21632 25964 21684
rect 26016 21632 26022 21684
rect 26602 21632 26608 21684
rect 26660 21672 26666 21684
rect 26697 21675 26755 21681
rect 26697 21672 26709 21675
rect 26660 21644 26709 21672
rect 26660 21632 26666 21644
rect 26697 21641 26709 21644
rect 26743 21672 26755 21675
rect 27614 21672 27620 21684
rect 26743 21644 27620 21672
rect 26743 21641 26755 21644
rect 26697 21635 26755 21641
rect 27614 21632 27620 21644
rect 27672 21632 27678 21684
rect 27709 21675 27767 21681
rect 27709 21641 27721 21675
rect 27755 21672 27767 21675
rect 35618 21672 35624 21684
rect 27755 21644 35624 21672
rect 27755 21641 27767 21644
rect 27709 21635 27767 21641
rect 35618 21632 35624 21644
rect 35676 21632 35682 21684
rect 23566 21604 23572 21616
rect 14700 21576 16896 21604
rect 20272 21576 23572 21604
rect 14700 21564 14706 21576
rect 12526 21496 12532 21548
rect 12584 21536 12590 21548
rect 13081 21539 13139 21545
rect 13081 21536 13093 21539
rect 12584 21508 13093 21536
rect 12584 21496 12590 21508
rect 13081 21505 13093 21508
rect 13127 21505 13139 21539
rect 13081 21499 13139 21505
rect 15930 21496 15936 21548
rect 15988 21496 15994 21548
rect 16868 21545 16896 21576
rect 23566 21564 23572 21576
rect 23624 21564 23630 21616
rect 23661 21607 23719 21613
rect 23661 21573 23673 21607
rect 23707 21604 23719 21607
rect 23934 21604 23940 21616
rect 23707 21576 23940 21604
rect 23707 21573 23719 21576
rect 23661 21567 23719 21573
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 28721 21607 28779 21613
rect 28721 21604 28733 21607
rect 27540 21576 28733 21604
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21505 16911 21539
rect 18598 21536 18604 21548
rect 16853 21499 16911 21505
rect 17236 21508 18604 21536
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 12176 21440 12265 21468
rect 10410 21360 10416 21412
rect 10468 21400 10474 21412
rect 12176 21400 12204 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 16209 21471 16267 21477
rect 16209 21437 16221 21471
rect 16255 21468 16267 21471
rect 17236 21468 17264 21508
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 20806 21536 20812 21548
rect 20102 21522 20812 21536
rect 20088 21508 20812 21522
rect 16255 21440 17264 21468
rect 16255 21437 16267 21440
rect 16209 21431 16267 21437
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21468 18751 21471
rect 18739 21440 18828 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 10468 21372 12204 21400
rect 10468 21360 10474 21372
rect 8938 21332 8944 21344
rect 7576 21304 8944 21332
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9861 21335 9919 21341
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 11146 21332 11152 21344
rect 9907 21304 11152 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11514 21332 11520 21344
rect 11379 21304 11520 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 11790 21292 11796 21344
rect 11848 21292 11854 21344
rect 12176 21332 12204 21372
rect 15562 21360 15568 21412
rect 15620 21360 15626 21412
rect 16666 21360 16672 21412
rect 16724 21400 16730 21412
rect 18598 21400 18604 21412
rect 16724 21372 18604 21400
rect 16724 21360 16730 21372
rect 18598 21360 18604 21372
rect 18656 21360 18662 21412
rect 12802 21332 12808 21344
rect 12176 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 13998 21292 14004 21344
rect 14056 21332 14062 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 14056 21304 14841 21332
rect 14056 21292 14062 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 14829 21295 14887 21301
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 15289 21335 15347 21341
rect 15289 21332 15301 21335
rect 15068 21304 15301 21332
rect 15068 21292 15074 21304
rect 15289 21301 15301 21304
rect 15335 21332 15347 21335
rect 18690 21332 18696 21344
rect 15335 21304 18696 21332
rect 15335 21301 15347 21304
rect 15289 21295 15347 21301
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 18800 21332 18828 21440
rect 18966 21428 18972 21480
rect 19024 21428 19030 21480
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 20088 21468 20116 21508
rect 20806 21496 20812 21508
rect 20864 21496 20870 21548
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21536 21327 21539
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 21315 21508 22385 21536
rect 21315 21505 21327 21508
rect 21269 21499 21327 21505
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22462 21496 22468 21548
rect 22520 21496 22526 21548
rect 23382 21496 23388 21548
rect 23440 21496 23446 21548
rect 26053 21539 26111 21545
rect 26053 21505 26065 21539
rect 26099 21536 26111 21539
rect 26510 21536 26516 21548
rect 26099 21508 26516 21536
rect 26099 21505 26111 21508
rect 26053 21499 26111 21505
rect 26510 21496 26516 21508
rect 26568 21496 26574 21548
rect 19116 21440 20116 21468
rect 22649 21471 22707 21477
rect 19116 21428 19122 21440
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 24670 21468 24676 21480
rect 22695 21440 24676 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 24670 21428 24676 21440
rect 24728 21468 24734 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24728 21440 25145 21468
rect 24728 21428 24734 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 26237 21471 26295 21477
rect 26237 21437 26249 21471
rect 26283 21468 26295 21471
rect 27540 21468 27568 21576
rect 28721 21573 28733 21576
rect 28767 21604 28779 21607
rect 28994 21604 29000 21616
rect 28767 21576 29000 21604
rect 28767 21573 28779 21576
rect 28721 21567 28779 21573
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 29178 21564 29184 21616
rect 29236 21564 29242 21616
rect 31021 21607 31079 21613
rect 31021 21573 31033 21607
rect 31067 21604 31079 21607
rect 31754 21604 31760 21616
rect 31067 21576 31760 21604
rect 31067 21573 31079 21576
rect 31021 21567 31079 21573
rect 31036 21536 31064 21567
rect 31754 21564 31760 21576
rect 31812 21564 31818 21616
rect 31846 21564 31852 21616
rect 31904 21604 31910 21616
rect 33965 21607 34023 21613
rect 33965 21604 33977 21607
rect 31904 21576 33977 21604
rect 31904 21564 31910 21576
rect 33965 21573 33977 21576
rect 34011 21573 34023 21607
rect 33965 21567 34023 21573
rect 35434 21564 35440 21616
rect 35492 21564 35498 21616
rect 29932 21508 31064 21536
rect 31113 21539 31171 21545
rect 26283 21440 27568 21468
rect 26283 21437 26295 21440
rect 26237 21431 26295 21437
rect 27798 21428 27804 21480
rect 27856 21428 27862 21480
rect 28350 21428 28356 21480
rect 28408 21468 28414 21480
rect 28445 21471 28503 21477
rect 28445 21468 28457 21471
rect 28408 21440 28457 21468
rect 28408 21428 28414 21440
rect 28445 21437 28457 21440
rect 28491 21437 28503 21471
rect 29932 21468 29960 21508
rect 31113 21505 31125 21539
rect 31159 21536 31171 21539
rect 31159 21508 32352 21536
rect 31159 21505 31171 21508
rect 31113 21499 31171 21505
rect 31205 21471 31263 21477
rect 31205 21468 31217 21471
rect 28445 21431 28503 21437
rect 28533 21440 29960 21468
rect 30208 21440 31217 21468
rect 20254 21360 20260 21412
rect 20312 21400 20318 21412
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 20312 21372 22017 21400
rect 20312 21360 20318 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 22738 21360 22744 21412
rect 22796 21400 22802 21412
rect 25866 21400 25872 21412
rect 22796 21372 23520 21400
rect 22796 21360 22802 21372
rect 19426 21332 19432 21344
rect 18800 21304 19432 21332
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 19702 21292 19708 21344
rect 19760 21332 19766 21344
rect 20441 21335 20499 21341
rect 20441 21332 20453 21335
rect 19760 21304 20453 21332
rect 19760 21292 19766 21304
rect 20441 21301 20453 21304
rect 20487 21301 20499 21335
rect 23492 21332 23520 21372
rect 24688 21372 25872 21400
rect 24688 21332 24716 21372
rect 25866 21360 25872 21372
rect 25924 21360 25930 21412
rect 26050 21360 26056 21412
rect 26108 21400 26114 21412
rect 27890 21400 27896 21412
rect 26108 21372 27896 21400
rect 26108 21360 26114 21372
rect 27890 21360 27896 21372
rect 27948 21360 27954 21412
rect 23492 21304 24716 21332
rect 20441 21295 20499 21301
rect 25222 21292 25228 21344
rect 25280 21332 25286 21344
rect 25593 21335 25651 21341
rect 25593 21332 25605 21335
rect 25280 21304 25605 21332
rect 25280 21292 25286 21304
rect 25593 21301 25605 21304
rect 25639 21301 25651 21335
rect 25593 21295 25651 21301
rect 25682 21292 25688 21344
rect 25740 21332 25746 21344
rect 27249 21335 27307 21341
rect 27249 21332 27261 21335
rect 25740 21304 27261 21332
rect 25740 21292 25746 21304
rect 27249 21301 27261 21304
rect 27295 21301 27307 21335
rect 27249 21295 27307 21301
rect 27614 21292 27620 21344
rect 27672 21332 27678 21344
rect 28533 21332 28561 21440
rect 30208 21344 30236 21440
rect 31205 21437 31217 21440
rect 31251 21437 31263 21471
rect 32122 21468 32128 21480
rect 31205 21431 31263 21437
rect 31312 21440 32128 21468
rect 30374 21360 30380 21412
rect 30432 21400 30438 21412
rect 31312 21400 31340 21440
rect 32122 21428 32128 21440
rect 32180 21428 32186 21480
rect 32324 21468 32352 21508
rect 32398 21496 32404 21548
rect 32456 21496 32462 21548
rect 32766 21496 32772 21548
rect 32824 21536 32830 21548
rect 33229 21539 33287 21545
rect 33229 21536 33241 21539
rect 32824 21508 33241 21536
rect 32824 21496 32830 21508
rect 33229 21505 33241 21508
rect 33275 21505 33287 21539
rect 33229 21499 33287 21505
rect 33410 21496 33416 21548
rect 33468 21536 33474 21548
rect 34517 21539 34575 21545
rect 34517 21536 34529 21539
rect 33468 21508 34529 21536
rect 33468 21496 33474 21508
rect 34517 21505 34529 21508
rect 34563 21505 34575 21539
rect 34517 21499 34575 21505
rect 47578 21496 47584 21548
rect 47636 21536 47642 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47636 21508 47961 21536
rect 47636 21496 47642 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 37366 21468 37372 21480
rect 32324 21440 37372 21468
rect 37366 21428 37372 21440
rect 37424 21428 37430 21480
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 30432 21372 31340 21400
rect 30432 21360 30438 21372
rect 31386 21360 31392 21412
rect 31444 21400 31450 21412
rect 31849 21403 31907 21409
rect 31849 21400 31861 21403
rect 31444 21372 31861 21400
rect 31444 21360 31450 21372
rect 31849 21369 31861 21372
rect 31895 21369 31907 21403
rect 31849 21363 31907 21369
rect 32306 21360 32312 21412
rect 32364 21400 32370 21412
rect 33505 21403 33563 21409
rect 33505 21400 33517 21403
rect 32364 21372 33517 21400
rect 32364 21360 32370 21372
rect 33505 21369 33517 21372
rect 33551 21369 33563 21403
rect 33505 21363 33563 21369
rect 33870 21360 33876 21412
rect 33928 21400 33934 21412
rect 34609 21403 34667 21409
rect 34609 21400 34621 21403
rect 33928 21372 34621 21400
rect 33928 21360 33934 21372
rect 34609 21369 34621 21372
rect 34655 21369 34667 21403
rect 34609 21363 34667 21369
rect 27672 21304 28561 21332
rect 27672 21292 27678 21304
rect 30190 21292 30196 21344
rect 30248 21292 30254 21344
rect 30650 21292 30656 21344
rect 30708 21292 30714 21344
rect 31570 21292 31576 21344
rect 31628 21332 31634 21344
rect 31757 21335 31815 21341
rect 31757 21332 31769 21335
rect 31628 21304 31769 21332
rect 31628 21292 31634 21304
rect 31757 21301 31769 21304
rect 31803 21332 31815 21335
rect 32030 21332 32036 21344
rect 31803 21304 32036 21332
rect 31803 21301 31815 21304
rect 31757 21295 31815 21301
rect 32030 21292 32036 21304
rect 32088 21292 32094 21344
rect 32398 21292 32404 21344
rect 32456 21332 32462 21344
rect 32493 21335 32551 21341
rect 32493 21332 32505 21335
rect 32456 21304 32505 21332
rect 32456 21292 32462 21304
rect 32493 21301 32505 21304
rect 32539 21301 32551 21335
rect 32493 21295 32551 21301
rect 32766 21292 32772 21344
rect 32824 21332 32830 21344
rect 33045 21335 33103 21341
rect 33045 21332 33057 21335
rect 32824 21304 33057 21332
rect 32824 21292 32830 21304
rect 33045 21301 33057 21304
rect 33091 21301 33103 21335
rect 33045 21295 33103 21301
rect 33962 21292 33968 21344
rect 34020 21332 34026 21344
rect 34057 21335 34115 21341
rect 34057 21332 34069 21335
rect 34020 21304 34069 21332
rect 34020 21292 34026 21304
rect 34057 21301 34069 21304
rect 34103 21301 34115 21335
rect 34057 21295 34115 21301
rect 34885 21335 34943 21341
rect 34885 21301 34897 21335
rect 34931 21332 34943 21335
rect 34974 21332 34980 21344
rect 34931 21304 34980 21332
rect 34931 21301 34943 21304
rect 34885 21295 34943 21301
rect 34974 21292 34980 21304
rect 35032 21292 35038 21344
rect 47578 21292 47584 21344
rect 47636 21292 47642 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 5077 21131 5135 21137
rect 5077 21128 5089 21131
rect 3476 21100 5089 21128
rect 3476 21088 3482 21100
rect 5077 21097 5089 21100
rect 5123 21097 5135 21131
rect 5077 21091 5135 21097
rect 5552 21100 7420 21128
rect 3605 21063 3663 21069
rect 3605 21029 3617 21063
rect 3651 21060 3663 21063
rect 4062 21060 4068 21072
rect 3651 21032 4068 21060
rect 3651 21029 3663 21032
rect 3605 21023 3663 21029
rect 4062 21020 4068 21032
rect 4120 21060 4126 21072
rect 5552 21060 5580 21100
rect 4120 21032 5580 21060
rect 4120 21020 4126 21032
rect 4246 20952 4252 21004
rect 4304 20952 4310 21004
rect 5721 20995 5779 21001
rect 5721 20961 5733 20995
rect 5767 20992 5779 20995
rect 7282 20992 7288 21004
rect 5767 20964 7288 20992
rect 5767 20961 5779 20964
rect 5721 20955 5779 20961
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 3326 20884 3332 20936
rect 3384 20924 3390 20936
rect 3973 20927 4031 20933
rect 3973 20924 3985 20927
rect 3384 20896 3985 20924
rect 3384 20884 3390 20896
rect 3973 20893 3985 20896
rect 4019 20893 4031 20927
rect 3973 20887 4031 20893
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 2774 20816 2780 20868
rect 2832 20816 2838 20868
rect 5258 20816 5264 20868
rect 5316 20856 5322 20868
rect 6178 20856 6184 20868
rect 5316 20828 6184 20856
rect 5316 20816 5322 20828
rect 6178 20816 6184 20828
rect 6236 20816 6242 20868
rect 7392 20856 7420 21100
rect 7466 21088 7472 21140
rect 7524 21128 7530 21140
rect 7653 21131 7711 21137
rect 7653 21128 7665 21131
rect 7524 21100 7665 21128
rect 7524 21088 7530 21100
rect 7653 21097 7665 21100
rect 7699 21097 7711 21131
rect 13725 21131 13783 21137
rect 7653 21091 7711 21097
rect 9508 21100 12434 21128
rect 7558 21020 7564 21072
rect 7616 21060 7622 21072
rect 9508 21060 9536 21100
rect 11790 21060 11796 21072
rect 7616 21032 9536 21060
rect 9600 21032 11796 21060
rect 7616 21020 7622 21032
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 8389 20995 8447 21001
rect 8389 20992 8401 20995
rect 7800 20964 8401 20992
rect 7800 20952 7806 20964
rect 8389 20961 8401 20964
rect 8435 20961 8447 20995
rect 9600 20992 9628 21032
rect 11790 21020 11796 21032
rect 11848 21020 11854 21072
rect 12406 21060 12434 21100
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 13814 21128 13820 21140
rect 13771 21100 13820 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 13814 21088 13820 21100
rect 13872 21128 13878 21140
rect 14458 21128 14464 21140
rect 13872 21100 14464 21128
rect 13872 21088 13878 21100
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 14553 21131 14611 21137
rect 14553 21097 14565 21131
rect 14599 21128 14611 21131
rect 16574 21128 16580 21140
rect 14599 21100 16580 21128
rect 14599 21097 14611 21100
rect 14553 21091 14611 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 17512 21100 21956 21128
rect 14918 21060 14924 21072
rect 12406 21032 14924 21060
rect 14918 21020 14924 21032
rect 14976 21020 14982 21072
rect 17218 21060 17224 21072
rect 15120 21032 17224 21060
rect 8389 20955 8447 20961
rect 9048 20964 9628 20992
rect 7466 20884 7472 20936
rect 7524 20924 7530 20936
rect 8205 20927 8263 20933
rect 8205 20924 8217 20927
rect 7524 20896 8217 20924
rect 7524 20884 7530 20896
rect 8205 20893 8217 20896
rect 8251 20893 8263 20927
rect 8205 20887 8263 20893
rect 8297 20927 8355 20933
rect 8297 20893 8309 20927
rect 8343 20924 8355 20927
rect 9048 20924 9076 20964
rect 9674 20952 9680 21004
rect 9732 20952 9738 21004
rect 10965 20995 11023 21001
rect 10965 20961 10977 20995
rect 11011 20992 11023 20995
rect 11011 20964 12434 20992
rect 11011 20961 11023 20964
rect 10965 20955 11023 20961
rect 8343 20896 9076 20924
rect 8343 20893 8355 20896
rect 8297 20887 8355 20893
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 11698 20884 11704 20936
rect 11756 20924 11762 20936
rect 11974 20924 11980 20936
rect 11756 20896 11980 20924
rect 11756 20884 11762 20896
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 12406 20924 12434 20964
rect 12618 20952 12624 21004
rect 12676 20952 12682 21004
rect 14277 20995 14335 21001
rect 14277 20961 14289 20995
rect 14323 20992 14335 20995
rect 15010 20992 15016 21004
rect 14323 20964 15016 20992
rect 14323 20961 14335 20964
rect 14277 20955 14335 20961
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 15120 21001 15148 21032
rect 17218 21020 17224 21032
rect 17276 21020 17282 21072
rect 15105 20995 15163 21001
rect 15105 20961 15117 20995
rect 15151 20961 15163 20995
rect 15105 20955 15163 20961
rect 16206 20952 16212 21004
rect 16264 20952 16270 21004
rect 16390 20952 16396 21004
rect 16448 20952 16454 21004
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 17512 20992 17540 21100
rect 17604 21032 18920 21060
rect 17604 21001 17632 21032
rect 17451 20964 17540 20992
rect 17589 20995 17647 21001
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 17589 20961 17601 20995
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 18782 20952 18788 21004
rect 18840 20952 18846 21004
rect 18892 20992 18920 21032
rect 21634 21020 21640 21072
rect 21692 21020 21698 21072
rect 21928 21060 21956 21100
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 22336 21100 23612 21128
rect 22336 21088 22342 21100
rect 23474 21060 23480 21072
rect 21928 21032 23480 21060
rect 23474 21020 23480 21032
rect 23532 21020 23538 21072
rect 23584 21060 23612 21100
rect 23750 21088 23756 21140
rect 23808 21128 23814 21140
rect 26050 21128 26056 21140
rect 23808 21100 26056 21128
rect 23808 21088 23814 21100
rect 26050 21088 26056 21100
rect 26108 21088 26114 21140
rect 26510 21088 26516 21140
rect 26568 21128 26574 21140
rect 28902 21128 28908 21140
rect 26568 21100 28908 21128
rect 26568 21088 26574 21100
rect 28902 21088 28908 21100
rect 28960 21088 28966 21140
rect 29730 21088 29736 21140
rect 29788 21128 29794 21140
rect 31846 21128 31852 21140
rect 29788 21100 31852 21128
rect 29788 21088 29794 21100
rect 31846 21088 31852 21100
rect 31904 21088 31910 21140
rect 33318 21088 33324 21140
rect 33376 21128 33382 21140
rect 34241 21131 34299 21137
rect 34241 21128 34253 21131
rect 33376 21100 34253 21128
rect 33376 21088 33382 21100
rect 34241 21097 34253 21100
rect 34287 21097 34299 21131
rect 34241 21091 34299 21097
rect 49050 21088 49056 21140
rect 49108 21128 49114 21140
rect 49421 21131 49479 21137
rect 49421 21128 49433 21131
rect 49108 21100 49433 21128
rect 49108 21088 49114 21100
rect 49421 21097 49433 21100
rect 49467 21097 49479 21131
rect 49421 21091 49479 21097
rect 23584 21032 23796 21060
rect 19702 20992 19708 21004
rect 18892 20964 19708 20992
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 22646 20992 22652 21004
rect 20128 20964 22652 20992
rect 20128 20952 20134 20964
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 23566 20992 23572 21004
rect 22787 20964 23572 20992
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 23566 20952 23572 20964
rect 23624 20952 23630 21004
rect 23768 21001 23796 21032
rect 24394 21020 24400 21072
rect 24452 21060 24458 21072
rect 25685 21063 25743 21069
rect 25685 21060 25697 21063
rect 24452 21032 25697 21060
rect 24452 21020 24458 21032
rect 25685 21029 25697 21032
rect 25731 21060 25743 21063
rect 25774 21060 25780 21072
rect 25731 21032 25780 21060
rect 25731 21029 25743 21032
rect 25685 21023 25743 21029
rect 25774 21020 25780 21032
rect 25832 21020 25838 21072
rect 27798 21060 27804 21072
rect 27356 21032 27804 21060
rect 23753 20995 23811 21001
rect 23753 20961 23765 20995
rect 23799 20961 23811 20995
rect 23753 20955 23811 20961
rect 23842 20952 23848 21004
rect 23900 20952 23906 21004
rect 25314 20952 25320 21004
rect 25372 20952 25378 21004
rect 25792 20992 25820 21020
rect 26050 20992 26056 21004
rect 25792 20964 26056 20992
rect 26050 20952 26056 20964
rect 26108 20952 26114 21004
rect 26329 20995 26387 21001
rect 26329 20961 26341 20995
rect 26375 20992 26387 20995
rect 27356 20992 27384 21032
rect 27798 21020 27804 21032
rect 27856 21020 27862 21072
rect 32493 21063 32551 21069
rect 32493 21029 32505 21063
rect 32539 21060 32551 21063
rect 35710 21060 35716 21072
rect 32539 21032 35716 21060
rect 32539 21029 32551 21032
rect 32493 21023 32551 21029
rect 35710 21020 35716 21032
rect 35768 21020 35774 21072
rect 26375 20964 27384 20992
rect 26375 20961 26387 20964
rect 26329 20955 26387 20961
rect 27706 20952 27712 21004
rect 27764 20992 27770 21004
rect 28537 20995 28595 21001
rect 28537 20992 28549 20995
rect 27764 20964 28549 20992
rect 27764 20952 27770 20964
rect 28537 20961 28549 20964
rect 28583 20961 28595 20995
rect 28537 20955 28595 20961
rect 29733 20995 29791 21001
rect 29733 20961 29745 20995
rect 29779 20992 29791 20995
rect 29914 20992 29920 21004
rect 29779 20964 29920 20992
rect 29779 20961 29791 20964
rect 29733 20955 29791 20961
rect 29914 20952 29920 20964
rect 29972 20952 29978 21004
rect 30006 20952 30012 21004
rect 30064 20952 30070 21004
rect 30098 20952 30104 21004
rect 30156 20992 30162 21004
rect 32582 20992 32588 21004
rect 30156 20964 32588 20992
rect 30156 20952 30162 20964
rect 32582 20952 32588 20964
rect 32640 20992 32646 21004
rect 33137 20995 33195 21001
rect 33137 20992 33149 20995
rect 32640 20964 33149 20992
rect 32640 20952 32646 20964
rect 33137 20961 33149 20964
rect 33183 20961 33195 20995
rect 33137 20955 33195 20961
rect 33505 20995 33563 21001
rect 33505 20961 33517 20995
rect 33551 20992 33563 20995
rect 33597 20995 33655 21001
rect 33597 20992 33609 20995
rect 33551 20964 33609 20992
rect 33551 20961 33563 20964
rect 33505 20955 33563 20961
rect 33597 20961 33609 20964
rect 33643 20992 33655 20995
rect 34146 20992 34152 21004
rect 33643 20964 34152 20992
rect 33643 20961 33655 20964
rect 33597 20955 33655 20961
rect 34146 20952 34152 20964
rect 34204 20952 34210 21004
rect 15194 20924 15200 20936
rect 12406 20896 15200 20924
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20924 16175 20927
rect 17494 20924 17500 20936
rect 16163 20896 17500 20924
rect 16163 20893 16175 20896
rect 16117 20887 16175 20893
rect 17494 20884 17500 20896
rect 17552 20884 17558 20936
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 18874 20924 18880 20936
rect 18555 20896 18880 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20924 22615 20927
rect 23290 20924 23296 20936
rect 22603 20896 23296 20924
rect 22603 20893 22615 20896
rect 22557 20887 22615 20893
rect 23290 20884 23296 20896
rect 23348 20884 23354 20936
rect 28261 20927 28319 20933
rect 28261 20893 28273 20927
rect 28307 20924 28319 20927
rect 28442 20924 28448 20936
rect 28307 20896 28448 20924
rect 28307 20893 28319 20896
rect 28261 20887 28319 20893
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 29822 20884 29828 20936
rect 29880 20924 29886 20936
rect 31113 20927 31171 20933
rect 31113 20924 31125 20927
rect 29880 20896 31125 20924
rect 29880 20884 29886 20896
rect 31113 20893 31125 20896
rect 31159 20893 31171 20927
rect 31113 20887 31171 20893
rect 32122 20884 32128 20936
rect 32180 20924 32186 20936
rect 32677 20927 32735 20933
rect 32677 20924 32689 20927
rect 32180 20896 32689 20924
rect 32180 20884 32186 20896
rect 32677 20893 32689 20896
rect 32723 20924 32735 20927
rect 32953 20927 33011 20933
rect 32953 20924 32965 20927
rect 32723 20896 32965 20924
rect 32723 20893 32735 20896
rect 32677 20887 32735 20893
rect 32953 20893 32965 20896
rect 32999 20893 33011 20927
rect 32953 20887 33011 20893
rect 10318 20856 10324 20868
rect 7392 20828 10324 20856
rect 10318 20816 10324 20828
rect 10376 20816 10382 20868
rect 11330 20816 11336 20868
rect 11388 20816 11394 20868
rect 15013 20859 15071 20865
rect 15013 20825 15025 20859
rect 15059 20856 15071 20859
rect 17862 20856 17868 20868
rect 15059 20828 17868 20856
rect 15059 20825 15071 20828
rect 15013 20819 15071 20825
rect 17862 20816 17868 20828
rect 17920 20816 17926 20868
rect 19978 20856 19984 20868
rect 18064 20828 19984 20856
rect 5902 20748 5908 20800
rect 5960 20788 5966 20800
rect 7193 20791 7251 20797
rect 7193 20788 7205 20791
rect 5960 20760 7205 20788
rect 5960 20748 5966 20760
rect 7193 20757 7205 20760
rect 7239 20757 7251 20791
rect 7193 20751 7251 20757
rect 7558 20748 7564 20800
rect 7616 20748 7622 20800
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 8846 20788 8852 20800
rect 7883 20760 8852 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 8846 20748 8852 20760
rect 8904 20748 8910 20800
rect 11422 20748 11428 20800
rect 11480 20748 11486 20800
rect 13906 20748 13912 20800
rect 13964 20748 13970 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 14921 20791 14979 20797
rect 14921 20788 14933 20791
rect 14792 20760 14933 20788
rect 14792 20748 14798 20760
rect 14921 20757 14933 20760
rect 14967 20757 14979 20791
rect 14921 20751 14979 20757
rect 15746 20748 15752 20800
rect 15804 20748 15810 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17034 20748 17040 20800
rect 17092 20788 17098 20800
rect 17313 20791 17371 20797
rect 17313 20788 17325 20791
rect 17092 20760 17325 20788
rect 17092 20748 17098 20760
rect 17313 20757 17325 20760
rect 17359 20788 17371 20791
rect 18064 20788 18092 20828
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 20990 20856 20996 20868
rect 20930 20828 20996 20856
rect 20990 20816 20996 20828
rect 21048 20856 21054 20868
rect 21634 20856 21640 20868
rect 21048 20828 21640 20856
rect 21048 20816 21054 20828
rect 21634 20816 21640 20828
rect 21692 20816 21698 20868
rect 21821 20859 21879 20865
rect 21821 20825 21833 20859
rect 21867 20856 21879 20859
rect 22370 20856 22376 20868
rect 21867 20828 22376 20856
rect 21867 20825 21879 20828
rect 21821 20819 21879 20825
rect 22370 20816 22376 20828
rect 22428 20816 22434 20868
rect 22465 20859 22523 20865
rect 22465 20825 22477 20859
rect 22511 20856 22523 20859
rect 23382 20856 23388 20868
rect 22511 20828 23388 20856
rect 22511 20825 22523 20828
rect 22465 20819 22523 20825
rect 23382 20816 23388 20828
rect 23440 20816 23446 20868
rect 25041 20859 25099 20865
rect 25041 20825 25053 20859
rect 25087 20856 25099 20859
rect 26234 20856 26240 20868
rect 25087 20828 26240 20856
rect 25087 20825 25099 20828
rect 25041 20819 25099 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 26418 20816 26424 20868
rect 26476 20856 26482 20868
rect 30650 20856 30656 20868
rect 26476 20828 26818 20856
rect 27724 20828 30656 20856
rect 26476 20816 26482 20828
rect 17359 20760 18092 20788
rect 18141 20791 18199 20797
rect 17359 20757 17371 20760
rect 17313 20751 17371 20757
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 18322 20788 18328 20800
rect 18187 20760 18328 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18322 20748 18328 20760
rect 18380 20748 18386 20800
rect 20530 20748 20536 20800
rect 20588 20788 20594 20800
rect 21177 20791 21235 20797
rect 21177 20788 21189 20791
rect 20588 20760 21189 20788
rect 20588 20748 20594 20760
rect 21177 20757 21189 20760
rect 21223 20757 21235 20791
rect 21177 20751 21235 20757
rect 22097 20791 22155 20797
rect 22097 20757 22109 20791
rect 22143 20788 22155 20791
rect 22278 20788 22284 20800
rect 22143 20760 22284 20788
rect 22143 20757 22155 20760
rect 22097 20751 22155 20757
rect 22278 20748 22284 20760
rect 22336 20748 22342 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 22704 20760 23305 20788
rect 22704 20748 22710 20760
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 23293 20751 23351 20757
rect 23658 20748 23664 20800
rect 23716 20748 23722 20800
rect 23750 20748 23756 20800
rect 23808 20788 23814 20800
rect 24673 20791 24731 20797
rect 24673 20788 24685 20791
rect 23808 20760 24685 20788
rect 23808 20748 23814 20760
rect 24673 20757 24685 20760
rect 24719 20757 24731 20791
rect 24673 20751 24731 20757
rect 25133 20791 25191 20797
rect 25133 20757 25145 20791
rect 25179 20788 25191 20791
rect 27724 20788 27752 20828
rect 30650 20816 30656 20828
rect 30708 20816 30714 20868
rect 31849 20859 31907 20865
rect 31849 20856 31861 20859
rect 30760 20828 31861 20856
rect 25179 20760 27752 20788
rect 27801 20791 27859 20797
rect 25179 20757 25191 20760
rect 25133 20751 25191 20757
rect 27801 20757 27813 20791
rect 27847 20788 27859 20791
rect 27890 20788 27896 20800
rect 27847 20760 27896 20788
rect 27847 20757 27859 20760
rect 27801 20751 27859 20757
rect 27890 20748 27896 20760
rect 27948 20748 27954 20800
rect 28994 20748 29000 20800
rect 29052 20788 29058 20800
rect 30760 20788 30788 20828
rect 31849 20825 31861 20828
rect 31895 20825 31907 20859
rect 31849 20819 31907 20825
rect 32030 20816 32036 20868
rect 32088 20816 32094 20868
rect 29052 20760 30788 20788
rect 29052 20748 29058 20760
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 34054 20748 34060 20800
rect 34112 20748 34118 20800
rect 46198 20748 46204 20800
rect 46256 20788 46262 20800
rect 47486 20788 47492 20800
rect 46256 20760 47492 20788
rect 46256 20748 46262 20760
rect 47486 20748 47492 20760
rect 47544 20748 47550 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5629 20587 5687 20593
rect 5629 20553 5641 20587
rect 5675 20584 5687 20587
rect 6914 20584 6920 20596
rect 5675 20556 6920 20584
rect 5675 20553 5687 20556
rect 5629 20547 5687 20553
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 9490 20584 9496 20596
rect 8772 20556 9496 20584
rect 4614 20476 4620 20528
rect 4672 20516 4678 20528
rect 8772 20525 8800 20556
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 9600 20556 12909 20584
rect 8757 20519 8815 20525
rect 4672 20488 7052 20516
rect 4672 20476 4678 20488
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 3421 20451 3479 20457
rect 3421 20448 3433 20451
rect 1872 20420 3433 20448
rect 934 20340 940 20392
rect 992 20380 998 20392
rect 1872 20380 1900 20420
rect 3421 20417 3433 20420
rect 3467 20417 3479 20451
rect 3421 20411 3479 20417
rect 5721 20451 5779 20457
rect 5721 20417 5733 20451
rect 5767 20448 5779 20451
rect 5994 20448 6000 20460
rect 5767 20420 6000 20448
rect 5767 20417 5779 20420
rect 5721 20411 5779 20417
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6144 20420 6561 20448
rect 6144 20408 6150 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 992 20352 1900 20380
rect 992 20340 998 20352
rect 2038 20340 2044 20392
rect 2096 20340 2102 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 7024 20389 7052 20488
rect 8757 20485 8769 20519
rect 8803 20485 8815 20519
rect 9600 20516 9628 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13035 20556 15792 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 8757 20479 8815 20485
rect 9416 20488 9628 20516
rect 7558 20408 7564 20460
rect 7616 20448 7622 20460
rect 9416 20448 9444 20488
rect 10134 20476 10140 20528
rect 10192 20476 10198 20528
rect 11790 20476 11796 20528
rect 11848 20476 11854 20528
rect 12434 20476 12440 20528
rect 12492 20516 12498 20528
rect 13538 20516 13544 20528
rect 12492 20488 13544 20516
rect 12492 20476 12498 20488
rect 13538 20476 13544 20488
rect 13596 20516 13602 20528
rect 13596 20488 13768 20516
rect 13596 20476 13602 20488
rect 13740 20457 13768 20488
rect 13998 20476 14004 20528
rect 14056 20476 14062 20528
rect 14458 20476 14464 20528
rect 14516 20476 14522 20528
rect 15764 20516 15792 20556
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17000 20556 17509 20584
rect 17000 20544 17006 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 17497 20547 17555 20553
rect 18509 20587 18567 20593
rect 18509 20553 18521 20587
rect 18555 20553 18567 20587
rect 18509 20547 18567 20553
rect 18524 20516 18552 20547
rect 18874 20544 18880 20596
rect 18932 20544 18938 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19484 20556 22784 20584
rect 19484 20544 19490 20556
rect 15764 20488 18552 20516
rect 18800 20488 19104 20516
rect 7616 20420 9444 20448
rect 13725 20451 13783 20457
rect 7616 20408 7622 20420
rect 13725 20417 13737 20451
rect 13771 20417 13783 20451
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 13725 20411 13783 20417
rect 15212 20420 16037 20448
rect 15212 20392 15240 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16666 20448 16672 20460
rect 16025 20411 16083 20417
rect 16408 20420 16672 20448
rect 5905 20383 5963 20389
rect 5905 20349 5917 20383
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 5920 20312 5948 20343
rect 7282 20340 7288 20392
rect 7340 20380 7346 20392
rect 7340 20352 7604 20380
rect 7340 20340 7346 20352
rect 6086 20312 6092 20324
rect 5920 20284 6092 20312
rect 6086 20272 6092 20284
rect 6144 20272 6150 20324
rect 6178 20272 6184 20324
rect 6236 20312 6242 20324
rect 7466 20312 7472 20324
rect 6236 20284 7472 20312
rect 6236 20272 6242 20284
rect 7466 20272 7472 20284
rect 7524 20272 7530 20324
rect 7576 20312 7604 20352
rect 8938 20340 8944 20392
rect 8996 20380 9002 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 8996 20352 9413 20380
rect 8996 20340 9002 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 10962 20380 10968 20392
rect 9723 20352 10968 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 9122 20312 9128 20324
rect 7576 20284 9128 20312
rect 9122 20272 9128 20284
rect 9180 20272 9186 20324
rect 3878 20204 3884 20256
rect 3936 20244 3942 20256
rect 4062 20244 4068 20256
rect 3936 20216 4068 20244
rect 3936 20204 3942 20216
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 7282 20244 7288 20256
rect 5307 20216 7288 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 8202 20204 8208 20256
rect 8260 20244 8266 20256
rect 8297 20247 8355 20253
rect 8297 20244 8309 20247
rect 8260 20216 8309 20244
rect 8260 20204 8266 20216
rect 8297 20213 8309 20216
rect 8343 20213 8355 20247
rect 8297 20207 8355 20213
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 8849 20247 8907 20253
rect 8849 20244 8861 20247
rect 8444 20216 8861 20244
rect 8444 20204 8450 20216
rect 8849 20213 8861 20216
rect 8895 20213 8907 20247
rect 9416 20244 9444 20343
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13219 20352 15148 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 15120 20312 15148 20352
rect 15194 20340 15200 20392
rect 15252 20340 15258 20392
rect 16408 20380 16436 20420
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 16853 20383 16911 20389
rect 16853 20380 16865 20383
rect 15304 20352 16436 20380
rect 16592 20352 16865 20380
rect 15304 20312 15332 20352
rect 15120 20284 15332 20312
rect 15470 20272 15476 20324
rect 15528 20272 15534 20324
rect 9674 20244 9680 20256
rect 9416 20216 9680 20244
rect 8849 20207 8907 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 11146 20204 11152 20256
rect 11204 20204 11210 20256
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 11388 20216 11897 20244
rect 11388 20204 11394 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11885 20207 11943 20213
rect 12526 20204 12532 20256
rect 12584 20204 12590 20256
rect 13446 20204 13452 20256
rect 13504 20204 13510 20256
rect 13630 20204 13636 20256
rect 13688 20204 13694 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 16592 20244 16620 20352
rect 16853 20349 16865 20352
rect 16899 20380 16911 20383
rect 17420 20380 17448 20411
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 18800 20448 18828 20488
rect 17644 20420 18828 20448
rect 17644 20408 17650 20420
rect 16899 20352 17448 20380
rect 17681 20383 17739 20389
rect 16899 20349 16911 20352
rect 16853 20343 16911 20349
rect 17681 20349 17693 20383
rect 17727 20349 17739 20383
rect 17681 20343 17739 20349
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17037 20315 17095 20321
rect 17037 20312 17049 20315
rect 17000 20284 17049 20312
rect 17000 20272 17006 20284
rect 17037 20281 17049 20284
rect 17083 20281 17095 20315
rect 17696 20312 17724 20343
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 19076 20389 19104 20488
rect 19720 20457 19748 20556
rect 20990 20476 20996 20528
rect 21048 20476 21054 20528
rect 21910 20476 21916 20528
rect 21968 20516 21974 20528
rect 22756 20525 22784 20556
rect 23382 20544 23388 20596
rect 23440 20544 23446 20596
rect 24029 20587 24087 20593
rect 24029 20553 24041 20587
rect 24075 20584 24087 20587
rect 24946 20584 24952 20596
rect 24075 20556 24952 20584
rect 24075 20553 24087 20556
rect 24029 20547 24087 20553
rect 24946 20544 24952 20556
rect 25004 20584 25010 20596
rect 25498 20584 25504 20596
rect 25004 20556 25504 20584
rect 25004 20544 25010 20556
rect 25498 20544 25504 20556
rect 25556 20544 25562 20596
rect 26050 20544 26056 20596
rect 26108 20584 26114 20596
rect 26513 20587 26571 20593
rect 26513 20584 26525 20587
rect 26108 20556 26525 20584
rect 26108 20544 26114 20556
rect 26513 20553 26525 20556
rect 26559 20553 26571 20587
rect 26513 20547 26571 20553
rect 27062 20544 27068 20596
rect 27120 20584 27126 20596
rect 27157 20587 27215 20593
rect 27157 20584 27169 20587
rect 27120 20556 27169 20584
rect 27120 20544 27126 20556
rect 27157 20553 27169 20556
rect 27203 20553 27215 20587
rect 27157 20547 27215 20553
rect 27617 20587 27675 20593
rect 27617 20553 27629 20587
rect 27663 20584 27675 20587
rect 30834 20584 30840 20596
rect 27663 20556 30840 20584
rect 27663 20553 27675 20556
rect 27617 20547 27675 20553
rect 30834 20544 30840 20556
rect 30892 20544 30898 20596
rect 30929 20587 30987 20593
rect 30929 20553 30941 20587
rect 30975 20584 30987 20587
rect 31662 20584 31668 20596
rect 30975 20556 31668 20584
rect 30975 20553 30987 20556
rect 30929 20547 30987 20553
rect 31662 20544 31668 20556
rect 31720 20544 31726 20596
rect 31754 20544 31760 20596
rect 31812 20584 31818 20596
rect 32122 20584 32128 20596
rect 31812 20556 32128 20584
rect 31812 20544 31818 20556
rect 32122 20544 32128 20556
rect 32180 20544 32186 20596
rect 32214 20544 32220 20596
rect 32272 20584 32278 20596
rect 32861 20587 32919 20593
rect 32861 20584 32873 20587
rect 32272 20556 32873 20584
rect 32272 20544 32278 20556
rect 32861 20553 32873 20556
rect 32907 20553 32919 20587
rect 32861 20547 32919 20553
rect 22005 20519 22063 20525
rect 22005 20516 22017 20519
rect 21968 20488 22017 20516
rect 21968 20476 21974 20488
rect 22005 20485 22017 20488
rect 22051 20485 22063 20519
rect 22005 20479 22063 20485
rect 22741 20519 22799 20525
rect 22741 20485 22753 20519
rect 22787 20485 22799 20519
rect 26418 20516 26424 20528
rect 25806 20488 26424 20516
rect 22741 20479 22799 20485
rect 26418 20476 26424 20488
rect 26476 20476 26482 20528
rect 29086 20476 29092 20528
rect 29144 20476 29150 20528
rect 31021 20519 31079 20525
rect 31021 20485 31033 20519
rect 31067 20516 31079 20519
rect 37458 20516 37464 20528
rect 31067 20488 37464 20516
rect 31067 20485 31079 20488
rect 31021 20479 31079 20485
rect 37458 20476 37464 20488
rect 37516 20476 37522 20528
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 23198 20408 23204 20460
rect 23256 20448 23262 20460
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 23256 20420 24317 20448
rect 23256 20408 23262 20420
rect 24305 20417 24317 20420
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 26326 20408 26332 20460
rect 26384 20448 26390 20460
rect 26697 20451 26755 20457
rect 26697 20448 26709 20451
rect 26384 20420 26709 20448
rect 26384 20408 26390 20420
rect 26697 20417 26709 20420
rect 26743 20448 26755 20451
rect 27338 20448 27344 20460
rect 26743 20420 27344 20448
rect 26743 20417 26755 20420
rect 26697 20411 26755 20417
rect 27338 20408 27344 20420
rect 27396 20448 27402 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 27396 20420 27537 20448
rect 27396 20408 27402 20420
rect 27525 20417 27537 20420
rect 27571 20417 27583 20451
rect 27525 20411 27583 20417
rect 31938 20408 31944 20460
rect 31996 20448 32002 20460
rect 32677 20451 32735 20457
rect 32677 20448 32689 20451
rect 31996 20420 32689 20448
rect 31996 20408 32002 20420
rect 32677 20417 32689 20420
rect 32723 20417 32735 20451
rect 32677 20411 32735 20417
rect 18969 20383 19027 20389
rect 18969 20380 18981 20383
rect 18012 20352 18981 20380
rect 18012 20340 18018 20352
rect 18969 20349 18981 20352
rect 19015 20349 19027 20383
rect 18969 20343 19027 20349
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20380 19119 20383
rect 19981 20383 20039 20389
rect 19107 20352 19748 20380
rect 19107 20349 19119 20352
rect 19061 20343 19119 20349
rect 19610 20312 19616 20324
rect 17696 20284 19616 20312
rect 17037 20275 17095 20281
rect 19610 20272 19616 20284
rect 19668 20272 19674 20324
rect 13780 20216 16620 20244
rect 13780 20204 13786 20216
rect 16666 20204 16672 20256
rect 16724 20244 16730 20256
rect 18141 20247 18199 20253
rect 18141 20244 18153 20247
rect 16724 20216 18153 20244
rect 16724 20204 16730 20216
rect 18141 20213 18153 20216
rect 18187 20213 18199 20247
rect 19720 20244 19748 20352
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20622 20380 20628 20392
rect 20027 20352 20628 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 24581 20383 24639 20389
rect 24581 20349 24593 20383
rect 24627 20380 24639 20383
rect 24670 20380 24676 20392
rect 24627 20352 24676 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 24670 20340 24676 20352
rect 24728 20340 24734 20392
rect 26053 20383 26111 20389
rect 26053 20380 26065 20383
rect 25700 20352 26065 20380
rect 25700 20324 25728 20352
rect 26053 20349 26065 20352
rect 26099 20380 26111 20383
rect 27709 20383 27767 20389
rect 26099 20352 27292 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 25682 20272 25688 20324
rect 25740 20272 25746 20324
rect 27264 20312 27292 20352
rect 27709 20349 27721 20383
rect 27755 20349 27767 20383
rect 28350 20380 28356 20392
rect 27709 20343 27767 20349
rect 27816 20352 28356 20380
rect 27724 20312 27752 20343
rect 27264 20284 27752 20312
rect 21453 20247 21511 20253
rect 21453 20244 21465 20247
rect 19720 20216 21465 20244
rect 18141 20207 18199 20213
rect 21453 20213 21465 20216
rect 21499 20213 21511 20247
rect 21453 20207 21511 20213
rect 22738 20204 22744 20256
rect 22796 20244 22802 20256
rect 26510 20244 26516 20256
rect 22796 20216 26516 20244
rect 22796 20204 22802 20216
rect 26510 20204 26516 20216
rect 26568 20204 26574 20256
rect 27706 20204 27712 20256
rect 27764 20244 27770 20256
rect 27816 20244 27844 20352
rect 28350 20340 28356 20352
rect 28408 20340 28414 20392
rect 28629 20383 28687 20389
rect 28629 20349 28641 20383
rect 28675 20380 28687 20383
rect 30190 20380 30196 20392
rect 28675 20352 30196 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 30190 20340 30196 20352
rect 30248 20340 30254 20392
rect 30282 20340 30288 20392
rect 30340 20380 30346 20392
rect 31113 20383 31171 20389
rect 31113 20380 31125 20383
rect 30340 20352 31125 20380
rect 30340 20340 30346 20352
rect 31113 20349 31125 20352
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 31018 20272 31024 20324
rect 31076 20312 31082 20324
rect 31938 20312 31944 20324
rect 31076 20284 31944 20312
rect 31076 20272 31082 20284
rect 31938 20272 31944 20284
rect 31996 20312 32002 20324
rect 32309 20315 32367 20321
rect 32309 20312 32321 20315
rect 31996 20284 32321 20312
rect 31996 20272 32002 20284
rect 32309 20281 32321 20284
rect 32355 20281 32367 20315
rect 32309 20275 32367 20281
rect 27764 20216 27844 20244
rect 27764 20204 27770 20216
rect 28350 20204 28356 20256
rect 28408 20244 28414 20256
rect 30101 20247 30159 20253
rect 30101 20244 30113 20247
rect 28408 20216 30113 20244
rect 28408 20204 28414 20216
rect 30101 20213 30113 20216
rect 30147 20213 30159 20247
rect 30101 20207 30159 20213
rect 30558 20204 30564 20256
rect 30616 20204 30622 20256
rect 30926 20204 30932 20256
rect 30984 20244 30990 20256
rect 31570 20244 31576 20256
rect 30984 20216 31576 20244
rect 30984 20204 30990 20216
rect 31570 20204 31576 20216
rect 31628 20204 31634 20256
rect 31754 20204 31760 20256
rect 31812 20204 31818 20256
rect 32122 20204 32128 20256
rect 32180 20204 32186 20256
rect 32490 20204 32496 20256
rect 32548 20204 32554 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 3418 20000 3424 20052
rect 3476 20040 3482 20052
rect 3513 20043 3571 20049
rect 3513 20040 3525 20043
rect 3476 20012 3525 20040
rect 3476 20000 3482 20012
rect 3513 20009 3525 20012
rect 3559 20040 3571 20043
rect 3973 20043 4031 20049
rect 3973 20040 3985 20043
rect 3559 20012 3985 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 3973 20009 3985 20012
rect 4019 20040 4031 20043
rect 4157 20043 4215 20049
rect 4157 20040 4169 20043
rect 4019 20012 4169 20040
rect 4019 20009 4031 20012
rect 3973 20003 4031 20009
rect 4157 20009 4169 20012
rect 4203 20040 4215 20043
rect 5258 20040 5264 20052
rect 4203 20012 5264 20040
rect 4203 20009 4215 20012
rect 4157 20003 4215 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 6270 20000 6276 20052
rect 6328 20000 6334 20052
rect 7742 20000 7748 20052
rect 7800 20040 7806 20052
rect 8294 20040 8300 20052
rect 7800 20012 8300 20040
rect 7800 20000 7806 20012
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 10042 20040 10048 20052
rect 9048 20012 10048 20040
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 5442 19904 5448 19916
rect 4571 19876 5448 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 5442 19864 5448 19876
rect 5500 19904 5506 19916
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 5500 19876 6745 19904
rect 5500 19864 5506 19876
rect 6733 19873 6745 19876
rect 6779 19904 6791 19907
rect 8938 19904 8944 19916
rect 6779 19876 8944 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 4246 19836 4252 19848
rect 1811 19808 4252 19836
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 9048 19836 9076 20012
rect 10042 20000 10048 20012
rect 10100 20040 10106 20052
rect 10873 20043 10931 20049
rect 10873 20040 10885 20043
rect 10100 20012 10885 20040
rect 10100 20000 10106 20012
rect 10873 20009 10885 20012
rect 10919 20009 10931 20043
rect 10873 20003 10931 20009
rect 11790 20000 11796 20052
rect 11848 20040 11854 20052
rect 12989 20043 13047 20049
rect 11848 20012 12940 20040
rect 11848 20000 11854 20012
rect 12434 19972 12440 19984
rect 10796 19944 12440 19972
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 10796 19904 10824 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 11333 19907 11391 19913
rect 11333 19904 11345 19907
rect 9171 19876 10824 19904
rect 10888 19876 11345 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 8404 19808 9076 19836
rect 2777 19771 2835 19777
rect 2777 19737 2789 19771
rect 2823 19768 2835 19771
rect 2866 19768 2872 19780
rect 2823 19740 2872 19768
rect 2823 19737 2835 19740
rect 2777 19731 2835 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 3510 19728 3516 19780
rect 3568 19768 3574 19780
rect 4801 19771 4859 19777
rect 3568 19740 4016 19768
rect 3568 19728 3574 19740
rect 3418 19660 3424 19712
rect 3476 19660 3482 19712
rect 3878 19660 3884 19712
rect 3936 19660 3942 19712
rect 3988 19700 4016 19740
rect 4801 19737 4813 19771
rect 4847 19768 4859 19771
rect 5074 19768 5080 19780
rect 4847 19740 5080 19768
rect 4847 19737 4859 19740
rect 4801 19731 4859 19737
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 5258 19728 5264 19780
rect 5316 19728 5322 19780
rect 7009 19771 7067 19777
rect 7009 19737 7021 19771
rect 7055 19737 7067 19771
rect 7009 19731 7067 19737
rect 6638 19700 6644 19712
rect 3988 19672 6644 19700
rect 6638 19660 6644 19672
rect 6696 19660 6702 19712
rect 7024 19700 7052 19731
rect 7466 19728 7472 19780
rect 7524 19728 7530 19780
rect 8404 19700 8432 19808
rect 10410 19796 10416 19848
rect 10468 19836 10474 19848
rect 10888 19836 10916 19876
rect 11333 19873 11345 19876
rect 11379 19904 11391 19907
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 11379 19876 11437 19904
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 11425 19873 11437 19876
rect 11471 19904 11483 19907
rect 12066 19904 12072 19916
rect 11471 19876 12072 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 12345 19907 12403 19913
rect 12345 19873 12357 19907
rect 12391 19904 12403 19907
rect 12710 19904 12716 19916
rect 12391 19876 12716 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 10468 19808 10916 19836
rect 10468 19796 10474 19808
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11296 19808 12173 19836
rect 11296 19796 11302 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12912 19836 12940 20012
rect 12989 20009 13001 20043
rect 13035 20040 13047 20043
rect 13354 20040 13360 20052
rect 13035 20012 13360 20040
rect 13035 20009 13047 20012
rect 12989 20003 13047 20009
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 17954 20040 17960 20052
rect 13464 20012 17960 20040
rect 13464 19913 13492 20012
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19886 20040 19892 20052
rect 18739 20012 19892 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19886 20000 19892 20012
rect 19944 20000 19950 20052
rect 20714 20000 20720 20052
rect 20772 20040 20778 20052
rect 27617 20043 27675 20049
rect 20772 20012 27200 20040
rect 20772 20000 20778 20012
rect 14274 19932 14280 19984
rect 14332 19932 14338 19984
rect 14458 19932 14464 19984
rect 14516 19932 14522 19984
rect 16761 19975 16819 19981
rect 16761 19941 16773 19975
rect 16807 19972 16819 19975
rect 17034 19972 17040 19984
rect 16807 19944 17040 19972
rect 16807 19941 16819 19944
rect 16761 19935 16819 19941
rect 17034 19932 17040 19944
rect 17092 19932 17098 19984
rect 17218 19932 17224 19984
rect 17276 19932 17282 19984
rect 19334 19972 19340 19984
rect 17328 19944 19340 19972
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19873 13507 19907
rect 13449 19867 13507 19873
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 13679 19876 14841 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14829 19873 14841 19876
rect 14875 19904 14887 19907
rect 15470 19904 15476 19916
rect 14875 19876 15476 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 17328 19904 17356 19944
rect 19334 19932 19340 19944
rect 19392 19932 19398 19984
rect 27172 19972 27200 20012
rect 27617 20009 27629 20043
rect 27663 20040 27675 20043
rect 27798 20040 27804 20052
rect 27663 20012 27804 20040
rect 27663 20009 27675 20012
rect 27617 20003 27675 20009
rect 27798 20000 27804 20012
rect 27856 20000 27862 20052
rect 29730 20000 29736 20052
rect 29788 20000 29794 20052
rect 29914 20000 29920 20052
rect 29972 20040 29978 20052
rect 30193 20043 30251 20049
rect 30193 20040 30205 20043
rect 29972 20012 30205 20040
rect 29972 20000 29978 20012
rect 30193 20009 30205 20012
rect 30239 20009 30251 20043
rect 30193 20003 30251 20009
rect 31018 20000 31024 20052
rect 31076 20040 31082 20052
rect 31849 20043 31907 20049
rect 31849 20040 31861 20043
rect 31076 20012 31861 20040
rect 31076 20000 31082 20012
rect 31849 20009 31861 20012
rect 31895 20040 31907 20043
rect 35158 20040 35164 20052
rect 31895 20012 35164 20040
rect 31895 20009 31907 20012
rect 31849 20003 31907 20009
rect 35158 20000 35164 20012
rect 35216 20000 35222 20052
rect 49234 20040 49240 20052
rect 35866 20012 49240 20040
rect 35866 19972 35894 20012
rect 49234 20000 49240 20012
rect 49292 20000 49298 20052
rect 27172 19944 35894 19972
rect 16080 19876 17356 19904
rect 17865 19907 17923 19913
rect 16080 19864 16086 19876
rect 17865 19873 17877 19907
rect 17911 19904 17923 19907
rect 18966 19904 18972 19916
rect 17911 19876 18972 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 18966 19864 18972 19876
rect 19024 19904 19030 19916
rect 19426 19904 19432 19916
rect 19024 19876 19432 19904
rect 19024 19864 19030 19876
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 20530 19904 20536 19916
rect 19668 19876 20536 19904
rect 19668 19864 19674 19876
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 21542 19864 21548 19916
rect 21600 19904 21606 19916
rect 22005 19907 22063 19913
rect 22005 19904 22017 19907
rect 21600 19876 22017 19904
rect 21600 19864 21606 19876
rect 22005 19873 22017 19876
rect 22051 19904 22063 19907
rect 23842 19904 23848 19916
rect 22051 19876 23848 19904
rect 22051 19873 22063 19876
rect 22005 19867 22063 19873
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 25317 19907 25375 19913
rect 25317 19873 25329 19907
rect 25363 19904 25375 19907
rect 26142 19904 26148 19916
rect 25363 19876 26148 19904
rect 25363 19873 25375 19876
rect 25317 19867 25375 19873
rect 26142 19864 26148 19876
rect 26200 19864 26206 19916
rect 26510 19864 26516 19916
rect 26568 19904 26574 19916
rect 26568 19876 27384 19904
rect 26568 19864 26574 19876
rect 12912 19808 13492 19836
rect 12161 19799 12219 19805
rect 9401 19771 9459 19777
rect 9401 19737 9413 19771
rect 9447 19737 9459 19771
rect 9401 19731 9459 19737
rect 7024 19672 8432 19700
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8570 19700 8576 19712
rect 8527 19672 8576 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 9416 19700 9444 19731
rect 10134 19728 10140 19780
rect 10192 19728 10198 19780
rect 12710 19728 12716 19780
rect 12768 19768 12774 19780
rect 13357 19771 13415 19777
rect 13357 19768 13369 19771
rect 12768 19740 13369 19768
rect 12768 19728 12774 19740
rect 13357 19737 13369 19740
rect 13403 19737 13415 19771
rect 13464 19768 13492 19808
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 18322 19836 18328 19848
rect 17727 19808 18328 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19058 19836 19064 19848
rect 18923 19808 19064 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19702 19796 19708 19848
rect 19760 19836 19766 19848
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 19760 19808 20269 19836
rect 19760 19796 19766 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 22370 19796 22376 19848
rect 22428 19836 22434 19848
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22428 19808 22569 19836
rect 22428 19796 22434 19808
rect 22557 19805 22569 19808
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 23753 19839 23811 19845
rect 23753 19805 23765 19839
rect 23799 19836 23811 19839
rect 24946 19836 24952 19848
rect 23799 19808 24952 19836
rect 23799 19805 23811 19808
rect 23753 19799 23811 19805
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25832 19808 25881 19836
rect 25832 19796 25838 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 27356 19836 27384 19876
rect 27614 19864 27620 19916
rect 27672 19904 27678 19916
rect 28629 19907 28687 19913
rect 28629 19904 28641 19907
rect 27672 19876 28641 19904
rect 27672 19864 27678 19876
rect 28629 19873 28641 19876
rect 28675 19873 28687 19907
rect 31297 19907 31355 19913
rect 31297 19904 31309 19907
rect 28629 19867 28687 19873
rect 29012 19876 31309 19904
rect 29012 19848 29040 19876
rect 31297 19873 31309 19876
rect 31343 19873 31355 19907
rect 31297 19867 31355 19873
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 27356 19808 28365 19836
rect 25869 19799 25927 19805
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 28994 19796 29000 19848
rect 29052 19796 29058 19848
rect 29914 19796 29920 19848
rect 29972 19796 29978 19848
rect 31205 19839 31263 19845
rect 31205 19805 31217 19839
rect 31251 19836 31263 19839
rect 41322 19836 41328 19848
rect 31251 19808 41328 19836
rect 31251 19805 31263 19808
rect 31205 19799 31263 19805
rect 41322 19796 41328 19808
rect 41380 19796 41386 19848
rect 14826 19768 14832 19780
rect 13464 19740 14832 19768
rect 13357 19731 13415 19737
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 16666 19768 16672 19780
rect 15212 19740 15318 19768
rect 16224 19740 16672 19768
rect 11146 19700 11152 19712
rect 9416 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11790 19660 11796 19712
rect 11848 19660 11854 19712
rect 12253 19703 12311 19709
rect 12253 19669 12265 19703
rect 12299 19700 12311 19703
rect 13262 19700 13268 19712
rect 12299 19672 13268 19700
rect 12299 19669 12311 19672
rect 12253 19663 12311 19669
rect 13262 19660 13268 19672
rect 13320 19660 13326 19712
rect 13814 19660 13820 19712
rect 13872 19660 13878 19712
rect 14458 19660 14464 19712
rect 14516 19700 14522 19712
rect 15212 19700 15240 19740
rect 16224 19700 16252 19740
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19768 17003 19771
rect 19613 19771 19671 19777
rect 19613 19768 19625 19771
rect 16991 19740 19625 19768
rect 16991 19737 17003 19740
rect 16945 19731 17003 19737
rect 19613 19737 19625 19740
rect 19659 19768 19671 19771
rect 19978 19768 19984 19780
rect 19659 19740 19984 19768
rect 19659 19737 19671 19740
rect 19613 19731 19671 19737
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 20990 19728 20996 19780
rect 21048 19728 21054 19780
rect 23566 19728 23572 19780
rect 23624 19768 23630 19780
rect 25498 19768 25504 19780
rect 23624 19740 25504 19768
rect 23624 19728 23630 19740
rect 25498 19728 25504 19740
rect 25556 19768 25562 19780
rect 26145 19771 26203 19777
rect 26145 19768 26157 19771
rect 25556 19740 26157 19768
rect 25556 19728 25562 19740
rect 26145 19737 26157 19740
rect 26191 19737 26203 19771
rect 26145 19731 26203 19737
rect 26418 19728 26424 19780
rect 26476 19768 26482 19780
rect 26602 19768 26608 19780
rect 26476 19740 26608 19768
rect 26476 19728 26482 19740
rect 26602 19728 26608 19740
rect 26660 19728 26666 19780
rect 29822 19768 29828 19780
rect 27724 19740 29828 19768
rect 14516 19672 16252 19700
rect 16301 19703 16359 19709
rect 14516 19660 14522 19672
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 16390 19700 16396 19712
rect 16347 19672 16396 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 17586 19660 17592 19712
rect 17644 19660 17650 19712
rect 18414 19660 18420 19712
rect 18472 19660 18478 19712
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19886 19700 19892 19712
rect 19751 19672 19892 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 20070 19660 20076 19712
rect 20128 19700 20134 19712
rect 20714 19700 20720 19712
rect 20128 19672 20720 19700
rect 20128 19660 20134 19672
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 22428 19672 22661 19700
rect 22428 19660 22434 19672
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 22649 19663 22707 19669
rect 23290 19660 23296 19712
rect 23348 19660 23354 19712
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 23842 19660 23848 19712
rect 23900 19700 23906 19712
rect 24673 19703 24731 19709
rect 24673 19700 24685 19703
rect 23900 19672 24685 19700
rect 23900 19660 23906 19672
rect 24673 19669 24685 19672
rect 24719 19669 24731 19703
rect 24673 19663 24731 19669
rect 25038 19660 25044 19712
rect 25096 19660 25102 19712
rect 25133 19703 25191 19709
rect 25133 19669 25145 19703
rect 25179 19700 25191 19703
rect 27724 19700 27752 19740
rect 29822 19728 29828 19740
rect 29880 19728 29886 19780
rect 25179 19672 27752 19700
rect 25179 19669 25191 19672
rect 25133 19663 25191 19669
rect 27798 19660 27804 19712
rect 27856 19700 27862 19712
rect 27893 19703 27951 19709
rect 27893 19700 27905 19703
rect 27856 19672 27905 19700
rect 27856 19660 27862 19672
rect 27893 19669 27905 19672
rect 27939 19700 27951 19703
rect 29086 19700 29092 19712
rect 27939 19672 29092 19700
rect 27939 19669 27951 19672
rect 27893 19663 27951 19669
rect 29086 19660 29092 19672
rect 29144 19660 29150 19712
rect 30190 19660 30196 19712
rect 30248 19700 30254 19712
rect 30377 19703 30435 19709
rect 30377 19700 30389 19703
rect 30248 19672 30389 19700
rect 30248 19660 30254 19672
rect 30377 19669 30389 19672
rect 30423 19669 30435 19703
rect 30377 19663 30435 19669
rect 30742 19660 30748 19712
rect 30800 19660 30806 19712
rect 31018 19660 31024 19712
rect 31076 19700 31082 19712
rect 31113 19703 31171 19709
rect 31113 19700 31125 19703
rect 31076 19672 31125 19700
rect 31076 19660 31082 19672
rect 31113 19669 31125 19672
rect 31159 19669 31171 19703
rect 31113 19663 31171 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 5261 19499 5319 19505
rect 2608 19468 4476 19496
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19360 1823 19363
rect 2608 19360 2636 19468
rect 4338 19388 4344 19440
rect 4396 19388 4402 19440
rect 4448 19428 4476 19468
rect 5261 19465 5273 19499
rect 5307 19496 5319 19499
rect 5442 19496 5448 19508
rect 5307 19468 5448 19496
rect 5307 19465 5319 19468
rect 5261 19459 5319 19465
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 5718 19456 5724 19508
rect 5776 19456 5782 19508
rect 5828 19468 6408 19496
rect 4448 19400 5580 19428
rect 1811 19332 2636 19360
rect 1811 19329 1823 19332
rect 1765 19323 1823 19329
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 4890 19360 4896 19372
rect 3651 19332 4896 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 4890 19320 4896 19332
rect 4948 19320 4954 19372
rect 5552 19292 5580 19400
rect 5629 19363 5687 19369
rect 5629 19329 5641 19363
rect 5675 19360 5687 19363
rect 5718 19360 5724 19372
rect 5675 19332 5724 19360
rect 5675 19329 5687 19332
rect 5629 19323 5687 19329
rect 5718 19320 5724 19332
rect 5776 19320 5782 19372
rect 5828 19292 5856 19468
rect 6380 19428 6408 19468
rect 6454 19456 6460 19508
rect 6512 19496 6518 19508
rect 10318 19496 10324 19508
rect 6512 19468 10324 19496
rect 6512 19456 6518 19468
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 10413 19499 10471 19505
rect 10413 19465 10425 19499
rect 10459 19496 10471 19499
rect 11882 19496 11888 19508
rect 10459 19468 11888 19496
rect 10459 19465 10471 19468
rect 10413 19459 10471 19465
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 14550 19496 14556 19508
rect 11992 19468 14556 19496
rect 11992 19440 12020 19468
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14826 19456 14832 19508
rect 14884 19456 14890 19508
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 16942 19496 16948 19508
rect 16632 19468 16948 19496
rect 16632 19456 16638 19468
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 17034 19456 17040 19508
rect 17092 19496 17098 19508
rect 17221 19499 17279 19505
rect 17221 19496 17233 19499
rect 17092 19468 17233 19496
rect 17092 19456 17098 19468
rect 17221 19465 17233 19468
rect 17267 19465 17279 19499
rect 17221 19459 17279 19465
rect 17865 19499 17923 19505
rect 17865 19465 17877 19499
rect 17911 19465 17923 19499
rect 17865 19459 17923 19465
rect 7098 19428 7104 19440
rect 6380 19400 7104 19428
rect 7098 19388 7104 19400
rect 7156 19388 7162 19440
rect 8478 19388 8484 19440
rect 8536 19428 8542 19440
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 8536 19400 9321 19428
rect 8536 19388 8542 19400
rect 9309 19397 9321 19400
rect 9355 19397 9367 19431
rect 11974 19428 11980 19440
rect 9309 19391 9367 19397
rect 11716 19400 11980 19428
rect 6549 19363 6607 19369
rect 6549 19360 6561 19363
rect 6288 19332 6561 19360
rect 5552 19264 5856 19292
rect 5902 19252 5908 19304
rect 5960 19252 5966 19304
rect 2682 19184 2688 19236
rect 2740 19224 2746 19236
rect 6288 19224 6316 19332
rect 6549 19329 6561 19332
rect 6595 19329 6607 19363
rect 6549 19323 6607 19329
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 7469 19363 7527 19369
rect 7469 19360 7481 19363
rect 6696 19332 7481 19360
rect 6696 19320 6702 19332
rect 7469 19329 7481 19332
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 8754 19360 8760 19372
rect 8619 19332 8760 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 8754 19320 8760 19332
rect 8812 19320 8818 19372
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10778 19360 10784 19372
rect 10367 19332 10784 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 11606 19360 11612 19372
rect 10919 19332 11612 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 11716 19369 11744 19400
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 12066 19388 12072 19440
rect 12124 19428 12130 19440
rect 12124 19400 12466 19428
rect 12124 19388 12130 19400
rect 13262 19388 13268 19440
rect 13320 19428 13326 19440
rect 17880 19428 17908 19459
rect 19058 19456 19064 19508
rect 19116 19456 19122 19508
rect 19426 19456 19432 19508
rect 19484 19496 19490 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 19484 19468 21465 19496
rect 19484 19456 19490 19468
rect 21453 19465 21465 19468
rect 21499 19465 21511 19499
rect 21453 19459 21511 19465
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 23290 19496 23296 19508
rect 22419 19468 23296 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 26421 19499 26479 19505
rect 26421 19496 26433 19499
rect 26292 19468 26433 19496
rect 26292 19456 26298 19468
rect 26421 19465 26433 19468
rect 26467 19465 26479 19499
rect 26421 19459 26479 19465
rect 27706 19456 27712 19508
rect 27764 19456 27770 19508
rect 30374 19496 30380 19508
rect 28276 19468 30380 19496
rect 13320 19400 17908 19428
rect 18325 19431 18383 19437
rect 13320 19388 13326 19400
rect 18325 19397 18337 19431
rect 18371 19428 18383 19431
rect 19334 19428 19340 19440
rect 18371 19400 19340 19428
rect 18371 19397 18383 19400
rect 18325 19391 18383 19397
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 20070 19428 20076 19440
rect 19720 19400 20076 19428
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 13906 19320 13912 19372
rect 13964 19360 13970 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 13964 19332 14749 19360
rect 13964 19320 13970 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 14844 19332 15056 19360
rect 10962 19252 10968 19304
rect 11020 19252 11026 19304
rect 11977 19295 12035 19301
rect 11977 19261 11989 19295
rect 12023 19292 12035 19295
rect 13630 19292 13636 19304
rect 12023 19264 13636 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13998 19252 14004 19304
rect 14056 19292 14062 19304
rect 14844 19292 14872 19332
rect 14056 19264 14872 19292
rect 14056 19252 14062 19264
rect 14918 19252 14924 19304
rect 14976 19252 14982 19304
rect 15028 19292 15056 19332
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 15896 19332 16988 19360
rect 15896 19320 15902 19332
rect 15028 19264 15976 19292
rect 8294 19224 8300 19236
rect 2740 19196 6316 19224
rect 6840 19196 8300 19224
rect 2740 19184 2746 19196
rect 5718 19116 5724 19168
rect 5776 19156 5782 19168
rect 6840 19156 6868 19196
rect 8294 19184 8300 19196
rect 8352 19224 8358 19236
rect 9490 19224 9496 19236
rect 8352 19196 9496 19224
rect 8352 19184 8358 19196
rect 9490 19184 9496 19196
rect 9548 19184 9554 19236
rect 10137 19227 10195 19233
rect 10137 19193 10149 19227
rect 10183 19224 10195 19227
rect 11698 19224 11704 19236
rect 10183 19196 11704 19224
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 11698 19184 11704 19196
rect 11756 19184 11762 19236
rect 13354 19184 13360 19236
rect 13412 19224 13418 19236
rect 13725 19227 13783 19233
rect 13725 19224 13737 19227
rect 13412 19196 13737 19224
rect 13412 19184 13418 19196
rect 13725 19193 13737 19196
rect 13771 19224 13783 19227
rect 13814 19224 13820 19236
rect 13771 19196 13820 19224
rect 13771 19193 13783 19196
rect 13725 19187 13783 19193
rect 13814 19184 13820 19196
rect 13872 19224 13878 19236
rect 13872 19196 14044 19224
rect 13872 19184 13878 19196
rect 5776 19128 6868 19156
rect 5776 19116 5782 19128
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 10870 19156 10876 19168
rect 6972 19128 10876 19156
rect 6972 19116 6978 19128
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 14016 19165 14044 19196
rect 14366 19184 14372 19236
rect 14424 19184 14430 19236
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 15841 19227 15899 19233
rect 15841 19224 15853 19227
rect 15160 19196 15853 19224
rect 15160 19184 15166 19196
rect 15841 19193 15853 19196
rect 15887 19193 15899 19227
rect 15948 19224 15976 19264
rect 16298 19252 16304 19304
rect 16356 19292 16362 19304
rect 16850 19292 16856 19304
rect 16356 19264 16856 19292
rect 16356 19252 16362 19264
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 16960 19292 16988 19332
rect 17402 19320 17408 19372
rect 17460 19320 17466 19372
rect 17862 19320 17868 19372
rect 17920 19360 17926 19372
rect 18233 19363 18291 19369
rect 18233 19360 18245 19363
rect 17920 19332 18245 19360
rect 17920 19320 17926 19332
rect 18233 19329 18245 19332
rect 18279 19360 18291 19363
rect 18279 19332 19012 19360
rect 18279 19329 18291 19332
rect 18233 19323 18291 19329
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 16960 19264 18429 19292
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18984 19292 19012 19332
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 19116 19332 19257 19360
rect 19116 19320 19122 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19720 19360 19748 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 21726 19428 21732 19440
rect 21468 19400 21732 19428
rect 19245 19323 19303 19329
rect 19352 19332 19748 19360
rect 19352 19292 19380 19332
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21468 19360 21496 19400
rect 21726 19388 21732 19400
rect 21784 19388 21790 19440
rect 22465 19431 22523 19437
rect 22465 19397 22477 19431
rect 22511 19428 22523 19431
rect 22646 19428 22652 19440
rect 22511 19400 22652 19428
rect 22511 19397 22523 19400
rect 22465 19391 22523 19397
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 23474 19388 23480 19440
rect 23532 19428 23538 19440
rect 24029 19431 24087 19437
rect 24029 19428 24041 19431
rect 23532 19400 24041 19428
rect 23532 19388 23538 19400
rect 24029 19397 24041 19400
rect 24075 19397 24087 19431
rect 24029 19391 24087 19397
rect 25314 19388 25320 19440
rect 25372 19428 25378 19440
rect 28166 19428 28172 19440
rect 25372 19400 28172 19428
rect 25372 19388 25378 19400
rect 28166 19388 28172 19400
rect 28224 19388 28230 19440
rect 21140 19332 21496 19360
rect 21140 19320 21146 19332
rect 21542 19320 21548 19372
rect 21600 19360 21606 19372
rect 23750 19360 23756 19372
rect 21600 19332 23756 19360
rect 21600 19320 21606 19332
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 24118 19320 24124 19372
rect 24176 19320 24182 19372
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19329 25007 19363
rect 24949 19323 25007 19329
rect 18984 19264 19380 19292
rect 18417 19255 18475 19261
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 22646 19292 22652 19304
rect 20680 19264 22652 19292
rect 20680 19252 20686 19264
rect 22646 19252 22652 19264
rect 22704 19252 22710 19304
rect 23842 19292 23848 19304
rect 22848 19264 23848 19292
rect 16758 19224 16764 19236
rect 15948 19196 16764 19224
rect 15841 19187 15899 19193
rect 16758 19184 16764 19196
rect 16816 19184 16822 19236
rect 16868 19224 16896 19252
rect 19720 19224 19748 19252
rect 16868 19196 19748 19224
rect 20990 19184 20996 19236
rect 21048 19224 21054 19236
rect 22848 19224 22876 19264
rect 23842 19252 23848 19264
rect 23900 19252 23906 19304
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24854 19292 24860 19304
rect 24351 19264 24860 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 23293 19227 23351 19233
rect 23293 19224 23305 19227
rect 21048 19196 22876 19224
rect 23032 19196 23305 19224
rect 21048 19184 21054 19196
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 11020 19128 13461 19156
rect 11020 19116 11026 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 14001 19159 14059 19165
rect 14001 19125 14013 19159
rect 14047 19156 14059 19159
rect 14185 19159 14243 19165
rect 14185 19156 14197 19159
rect 14047 19128 14197 19156
rect 14047 19125 14059 19128
rect 14001 19119 14059 19125
rect 14185 19125 14197 19128
rect 14231 19156 14243 19159
rect 15010 19156 15016 19168
rect 14231 19128 15016 19156
rect 14231 19125 14243 19128
rect 14185 19119 14243 19125
rect 15010 19116 15016 19128
rect 15068 19156 15074 19168
rect 15197 19159 15255 19165
rect 15197 19156 15209 19159
rect 15068 19128 15209 19156
rect 15068 19116 15074 19128
rect 15197 19125 15209 19128
rect 15243 19156 15255 19159
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 15243 19128 15393 19156
rect 15243 19125 15255 19128
rect 15197 19119 15255 19125
rect 15381 19125 15393 19128
rect 15427 19156 15439 19159
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15427 19128 16037 19156
rect 15427 19125 15439 19128
rect 15381 19119 15439 19125
rect 16025 19125 16037 19128
rect 16071 19156 16083 19159
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 16071 19128 16221 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 16209 19125 16221 19128
rect 16255 19156 16267 19159
rect 16393 19159 16451 19165
rect 16393 19156 16405 19159
rect 16255 19128 16405 19156
rect 16255 19125 16267 19128
rect 16209 19119 16267 19125
rect 16393 19125 16405 19128
rect 16439 19156 16451 19159
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16439 19128 16681 19156
rect 16439 19125 16451 19128
rect 16393 19119 16451 19125
rect 16669 19125 16681 19128
rect 16715 19156 16727 19159
rect 16853 19159 16911 19165
rect 16853 19156 16865 19159
rect 16715 19128 16865 19156
rect 16715 19125 16727 19128
rect 16669 19119 16727 19125
rect 16853 19125 16865 19128
rect 16899 19156 16911 19159
rect 17037 19159 17095 19165
rect 17037 19156 17049 19159
rect 16899 19128 17049 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 17037 19125 17049 19128
rect 17083 19156 17095 19159
rect 17497 19159 17555 19165
rect 17497 19156 17509 19159
rect 17083 19128 17509 19156
rect 17083 19125 17095 19128
rect 17037 19119 17095 19125
rect 17497 19125 17509 19128
rect 17543 19156 17555 19159
rect 17681 19159 17739 19165
rect 17681 19156 17693 19159
rect 17543 19128 17693 19156
rect 17543 19125 17555 19128
rect 17497 19119 17555 19125
rect 17681 19125 17693 19128
rect 17727 19156 17739 19159
rect 17862 19156 17868 19168
rect 17727 19128 17868 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18782 19116 18788 19168
rect 18840 19156 18846 19168
rect 19968 19159 20026 19165
rect 19968 19156 19980 19159
rect 18840 19128 19980 19156
rect 18840 19116 18846 19128
rect 19968 19125 19980 19128
rect 20014 19156 20026 19159
rect 21174 19156 21180 19168
rect 20014 19128 21180 19156
rect 20014 19125 20026 19128
rect 19968 19119 20026 19125
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 22002 19116 22008 19168
rect 22060 19116 22066 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 23032 19156 23060 19196
rect 23293 19193 23305 19196
rect 23339 19224 23351 19227
rect 24964 19224 24992 19323
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 28276 19360 28304 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 30469 19499 30527 19505
rect 30469 19465 30481 19499
rect 30515 19496 30527 19499
rect 34698 19496 34704 19508
rect 30515 19468 34704 19496
rect 30515 19465 30527 19468
rect 30469 19459 30527 19465
rect 34698 19456 34704 19468
rect 34756 19456 34762 19508
rect 29086 19388 29092 19440
rect 29144 19388 29150 19440
rect 30392 19428 30420 19456
rect 31018 19428 31024 19440
rect 30392 19400 31024 19428
rect 31018 19388 31024 19400
rect 31076 19388 31082 19440
rect 27396 19332 28304 19360
rect 27396 19320 27402 19332
rect 25774 19252 25780 19304
rect 25832 19252 25838 19304
rect 26970 19252 26976 19304
rect 27028 19252 27034 19304
rect 27154 19252 27160 19304
rect 27212 19292 27218 19304
rect 27908 19301 27936 19332
rect 30650 19320 30656 19372
rect 30708 19360 30714 19372
rect 31113 19363 31171 19369
rect 31113 19360 31125 19363
rect 30708 19332 31125 19360
rect 30708 19320 30714 19332
rect 31113 19329 31125 19332
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 27433 19295 27491 19301
rect 27433 19292 27445 19295
rect 27212 19264 27445 19292
rect 27212 19252 27218 19264
rect 27433 19261 27445 19264
rect 27479 19261 27491 19295
rect 27433 19255 27491 19261
rect 27893 19295 27951 19301
rect 27893 19261 27905 19295
rect 27939 19261 27951 19295
rect 27893 19255 27951 19261
rect 27982 19252 27988 19304
rect 28040 19292 28046 19304
rect 28261 19295 28319 19301
rect 28261 19292 28273 19295
rect 28040 19264 28273 19292
rect 28040 19252 28046 19264
rect 28261 19261 28273 19264
rect 28307 19261 28319 19295
rect 30466 19292 30472 19304
rect 28261 19255 28319 19261
rect 28368 19264 30472 19292
rect 25314 19224 25320 19236
rect 23339 19196 25320 19224
rect 23339 19193 23351 19196
rect 23293 19187 23351 19193
rect 25314 19184 25320 19196
rect 25372 19184 25378 19236
rect 25406 19184 25412 19236
rect 25464 19224 25470 19236
rect 28368 19224 28396 19264
rect 30466 19252 30472 19264
rect 30524 19252 30530 19304
rect 25464 19196 28396 19224
rect 25464 19184 25470 19196
rect 22152 19128 23060 19156
rect 23109 19159 23167 19165
rect 22152 19116 22158 19128
rect 23109 19125 23121 19159
rect 23155 19156 23167 19159
rect 23382 19156 23388 19168
rect 23155 19128 23388 19156
rect 23155 19125 23167 19128
rect 23109 19119 23167 19125
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 23566 19116 23572 19168
rect 23624 19156 23630 19168
rect 23661 19159 23719 19165
rect 23661 19156 23673 19159
rect 23624 19128 23673 19156
rect 23624 19116 23630 19128
rect 23661 19125 23673 19128
rect 23707 19125 23719 19159
rect 23661 19119 23719 19125
rect 26786 19116 26792 19168
rect 26844 19156 26850 19168
rect 27249 19159 27307 19165
rect 27249 19156 27261 19159
rect 26844 19128 27261 19156
rect 26844 19116 26850 19128
rect 27249 19125 27261 19128
rect 27295 19156 27307 19159
rect 27522 19156 27528 19168
rect 27295 19128 27528 19156
rect 27295 19125 27307 19128
rect 27249 19119 27307 19125
rect 27522 19116 27528 19128
rect 27580 19116 27586 19168
rect 28166 19116 28172 19168
rect 28224 19156 28230 19168
rect 28518 19159 28576 19165
rect 28518 19156 28530 19159
rect 28224 19128 28530 19156
rect 28224 19116 28230 19128
rect 28518 19125 28530 19128
rect 28564 19125 28576 19159
rect 28518 19119 28576 19125
rect 28626 19116 28632 19168
rect 28684 19156 28690 19168
rect 30009 19159 30067 19165
rect 30009 19156 30021 19159
rect 28684 19128 30021 19156
rect 28684 19116 28690 19128
rect 30009 19125 30021 19128
rect 30055 19156 30067 19159
rect 30282 19156 30288 19168
rect 30055 19128 30288 19156
rect 30055 19125 30067 19128
rect 30009 19119 30067 19125
rect 30282 19116 30288 19128
rect 30340 19116 30346 19168
rect 30926 19116 30932 19168
rect 30984 19116 30990 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 9766 18952 9772 18964
rect 3927 18924 9772 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 3988 18825 4016 18924
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 11112 18924 11621 18952
rect 11112 18912 11118 18924
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 11609 18915 11667 18921
rect 12268 18924 14657 18952
rect 8573 18887 8631 18893
rect 8573 18853 8585 18887
rect 8619 18884 8631 18887
rect 9122 18884 9128 18896
rect 8619 18856 9128 18884
rect 8619 18853 8631 18856
rect 8573 18847 8631 18853
rect 9122 18844 9128 18856
rect 9180 18884 9186 18896
rect 10134 18884 10140 18896
rect 9180 18856 10140 18884
rect 9180 18844 9186 18856
rect 10134 18844 10140 18856
rect 10192 18844 10198 18896
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1452 18788 2053 18816
rect 1452 18776 1458 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 3973 18819 4031 18825
rect 3973 18785 3985 18819
rect 4019 18785 4031 18819
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 3973 18779 4031 18785
rect 4632 18788 6837 18816
rect 4632 18760 4660 18788
rect 6825 18785 6837 18788
rect 6871 18816 6883 18819
rect 8478 18816 8484 18828
rect 6871 18788 8484 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10226 18816 10232 18828
rect 10091 18788 10232 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 11112 18788 11161 18816
rect 11112 18776 11118 18788
rect 11149 18785 11161 18788
rect 11195 18785 11207 18819
rect 11149 18779 11207 18785
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11296 18788 12173 18816
rect 11296 18776 11302 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 4246 18748 4252 18760
rect 1811 18720 4252 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9824 18720 9873 18748
rect 9824 18708 9830 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 10965 18751 11023 18757
rect 10965 18748 10977 18751
rect 10928 18720 10977 18748
rect 10928 18708 10934 18720
rect 10965 18717 10977 18720
rect 11011 18748 11023 18751
rect 12268 18748 12296 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 14645 18915 14703 18921
rect 14921 18955 14979 18961
rect 14921 18921 14933 18955
rect 14967 18952 14979 18955
rect 15010 18952 15016 18964
rect 14967 18924 15016 18952
rect 14967 18921 14979 18924
rect 14921 18915 14979 18921
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 22002 18952 22008 18964
rect 15120 18924 22008 18952
rect 13722 18844 13728 18896
rect 13780 18884 13786 18896
rect 14185 18887 14243 18893
rect 14185 18884 14197 18887
rect 13780 18856 14197 18884
rect 13780 18844 13786 18856
rect 14185 18853 14197 18856
rect 14231 18884 14243 18887
rect 14458 18884 14464 18896
rect 14231 18856 14464 18884
rect 14231 18853 14243 18856
rect 14185 18847 14243 18853
rect 14458 18844 14464 18856
rect 14516 18844 14522 18896
rect 13538 18776 13544 18828
rect 13596 18776 13602 18828
rect 13909 18819 13967 18825
rect 13909 18785 13921 18819
rect 13955 18816 13967 18819
rect 14826 18816 14832 18828
rect 13955 18788 14832 18816
rect 13955 18785 13967 18788
rect 13909 18779 13967 18785
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 14553 18751 14611 18757
rect 11011 18720 12296 18748
rect 12360 18720 12940 18748
rect 11011 18717 11023 18720
rect 10965 18711 11023 18717
rect 4893 18683 4951 18689
rect 4893 18649 4905 18683
rect 4939 18680 4951 18683
rect 4982 18680 4988 18692
rect 4939 18652 4988 18680
rect 4939 18649 4951 18652
rect 4893 18643 4951 18649
rect 4982 18640 4988 18652
rect 5040 18640 5046 18692
rect 6178 18680 6184 18692
rect 6118 18652 6184 18680
rect 6178 18640 6184 18652
rect 6236 18640 6242 18692
rect 6454 18640 6460 18692
rect 6512 18680 6518 18692
rect 7098 18680 7104 18692
rect 6512 18652 7104 18680
rect 6512 18640 6518 18652
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 7558 18640 7564 18692
rect 7616 18640 7622 18692
rect 8846 18680 8852 18692
rect 8404 18652 8852 18680
rect 2498 18572 2504 18624
rect 2556 18612 2562 18624
rect 3329 18615 3387 18621
rect 3329 18612 3341 18615
rect 2556 18584 3341 18612
rect 2556 18572 2562 18584
rect 3329 18581 3341 18584
rect 3375 18581 3387 18615
rect 3329 18575 3387 18581
rect 3602 18572 3608 18624
rect 3660 18572 3666 18624
rect 5074 18572 5080 18624
rect 5132 18612 5138 18624
rect 6365 18615 6423 18621
rect 6365 18612 6377 18615
rect 5132 18584 6377 18612
rect 5132 18572 5138 18584
rect 6365 18581 6377 18584
rect 6411 18612 6423 18615
rect 8404 18612 8432 18652
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 9125 18683 9183 18689
rect 9125 18649 9137 18683
rect 9171 18680 9183 18683
rect 10042 18680 10048 18692
rect 9171 18652 10048 18680
rect 9171 18649 9183 18652
rect 9125 18643 9183 18649
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 12360 18680 12388 18720
rect 10520 18652 12388 18680
rect 10520 18624 10548 18652
rect 12802 18640 12808 18692
rect 12860 18640 12866 18692
rect 12912 18680 12940 18720
rect 14553 18717 14565 18751
rect 14599 18748 14611 18751
rect 15120 18748 15148 18924
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22646 18912 22652 18964
rect 22704 18952 22710 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22704 18924 22937 18952
rect 22704 18912 22710 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 22925 18915 22983 18921
rect 23290 18912 23296 18964
rect 23348 18952 23354 18964
rect 25406 18952 25412 18964
rect 23348 18924 25412 18952
rect 23348 18912 23354 18924
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 25498 18912 25504 18964
rect 25556 18952 25562 18964
rect 27157 18955 27215 18961
rect 27157 18952 27169 18955
rect 25556 18924 27169 18952
rect 25556 18912 25562 18924
rect 27157 18921 27169 18924
rect 27203 18921 27215 18955
rect 46934 18952 46940 18964
rect 27157 18915 27215 18921
rect 31726 18924 46940 18952
rect 17586 18844 17592 18896
rect 17644 18884 17650 18896
rect 21082 18884 21088 18896
rect 17644 18856 21088 18884
rect 17644 18844 17650 18856
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 22462 18844 22468 18896
rect 22520 18884 22526 18896
rect 23385 18887 23443 18893
rect 23385 18884 23397 18887
rect 22520 18856 23397 18884
rect 22520 18844 22526 18856
rect 23385 18853 23397 18856
rect 23431 18853 23443 18887
rect 23385 18847 23443 18853
rect 26694 18844 26700 18896
rect 26752 18884 26758 18896
rect 31726 18884 31754 18924
rect 46934 18912 46940 18924
rect 46992 18912 46998 18964
rect 26752 18856 31754 18884
rect 26752 18844 26758 18856
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 16206 18816 16212 18828
rect 15243 18788 16212 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 16206 18776 16212 18788
rect 16264 18776 16270 18828
rect 16666 18816 16672 18828
rect 16592 18788 16672 18816
rect 14599 18720 15148 18748
rect 16592 18734 16620 18788
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 17494 18776 17500 18828
rect 17552 18776 17558 18828
rect 18598 18776 18604 18828
rect 18656 18776 18662 18828
rect 18693 18819 18751 18825
rect 18693 18785 18705 18819
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 18708 18748 18736 18779
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 19760 18788 20361 18816
rect 19760 18776 19766 18788
rect 20349 18785 20361 18788
rect 20395 18816 20407 18819
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 20395 18788 21189 18816
rect 20395 18785 20407 18788
rect 20349 18779 20407 18785
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 21876 18788 23520 18816
rect 21876 18776 21882 18788
rect 16816 18720 18736 18748
rect 19613 18751 19671 18757
rect 16816 18708 16822 18720
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19659 18720 20944 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 15010 18680 15016 18692
rect 12912 18652 15016 18680
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 15470 18640 15476 18692
rect 15528 18680 15534 18692
rect 20070 18680 20076 18692
rect 15528 18652 15884 18680
rect 15528 18640 15534 18652
rect 6411 18584 8432 18612
rect 6411 18581 6423 18584
rect 6365 18575 6423 18581
rect 9398 18572 9404 18624
rect 9456 18572 9462 18624
rect 9769 18615 9827 18621
rect 9769 18581 9781 18615
rect 9815 18612 9827 18615
rect 10502 18612 10508 18624
rect 9815 18584 10508 18612
rect 9815 18581 9827 18584
rect 9769 18575 9827 18581
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 10597 18615 10655 18621
rect 10597 18581 10609 18615
rect 10643 18612 10655 18615
rect 11698 18612 11704 18624
rect 10643 18584 11704 18612
rect 10643 18581 10655 18584
rect 10597 18575 10655 18581
rect 11698 18572 11704 18584
rect 11756 18612 11762 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11756 18584 11989 18612
rect 11756 18572 11762 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 14826 18612 14832 18624
rect 12124 18584 14832 18612
rect 12124 18572 12130 18584
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 15105 18615 15163 18621
rect 15105 18581 15117 18615
rect 15151 18612 15163 18615
rect 15286 18612 15292 18624
rect 15151 18584 15292 18612
rect 15151 18581 15163 18584
rect 15105 18575 15163 18581
rect 15286 18572 15292 18584
rect 15344 18572 15350 18624
rect 15856 18612 15884 18652
rect 16776 18652 20076 18680
rect 16390 18612 16396 18624
rect 15856 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18612 16454 18624
rect 16776 18612 16804 18652
rect 20070 18640 20076 18652
rect 20128 18640 20134 18692
rect 16448 18584 16804 18612
rect 16448 18572 16454 18584
rect 16942 18572 16948 18624
rect 17000 18572 17006 18624
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 18141 18615 18199 18621
rect 18141 18612 18153 18615
rect 18012 18584 18153 18612
rect 18012 18572 18018 18584
rect 18141 18581 18153 18584
rect 18187 18581 18199 18615
rect 18141 18575 18199 18581
rect 18509 18615 18567 18621
rect 18509 18581 18521 18615
rect 18555 18612 18567 18615
rect 18690 18612 18696 18624
rect 18555 18584 18696 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 19334 18572 19340 18624
rect 19392 18572 19398 18624
rect 20806 18572 20812 18624
rect 20864 18572 20870 18624
rect 20916 18612 20944 18720
rect 21726 18640 21732 18692
rect 21784 18680 21790 18692
rect 23492 18680 23520 18788
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 23716 18788 24593 18816
rect 23716 18776 23722 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25774 18816 25780 18828
rect 25455 18788 25780 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 29822 18776 29828 18828
rect 29880 18816 29886 18828
rect 30285 18819 30343 18825
rect 30285 18816 30297 18819
rect 29880 18788 30297 18816
rect 29880 18776 29886 18788
rect 30285 18785 30297 18788
rect 30331 18785 30343 18819
rect 30285 18779 30343 18785
rect 23566 18708 23572 18760
rect 23624 18708 23630 18760
rect 23842 18708 23848 18760
rect 23900 18748 23906 18760
rect 25041 18751 25099 18757
rect 25041 18748 25053 18751
rect 23900 18720 25053 18748
rect 23900 18708 23906 18720
rect 25041 18717 25053 18720
rect 25087 18717 25099 18751
rect 25041 18711 25099 18717
rect 26786 18708 26792 18760
rect 26844 18708 26850 18760
rect 27614 18708 27620 18760
rect 27672 18708 27678 18760
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 27893 18751 27951 18757
rect 27893 18748 27905 18751
rect 27764 18720 27905 18748
rect 27764 18708 27770 18720
rect 27893 18717 27905 18720
rect 27939 18717 27951 18751
rect 27893 18711 27951 18717
rect 30193 18751 30251 18757
rect 30193 18717 30205 18751
rect 30239 18748 30251 18751
rect 30558 18748 30564 18760
rect 30239 18720 30564 18748
rect 30239 18717 30251 18720
rect 30193 18711 30251 18717
rect 30558 18708 30564 18720
rect 30616 18708 30622 18760
rect 21784 18652 21942 18680
rect 23492 18652 25636 18680
rect 21784 18640 21790 18652
rect 22094 18612 22100 18624
rect 20916 18584 22100 18612
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 23937 18615 23995 18621
rect 23937 18612 23949 18615
rect 23900 18584 23949 18612
rect 23900 18572 23906 18584
rect 23937 18581 23949 18584
rect 23983 18581 23995 18615
rect 23937 18575 23995 18581
rect 24026 18572 24032 18624
rect 24084 18612 24090 18624
rect 24121 18615 24179 18621
rect 24121 18612 24133 18615
rect 24084 18584 24133 18612
rect 24084 18572 24090 18584
rect 24121 18581 24133 18584
rect 24167 18581 24179 18615
rect 25608 18612 25636 18652
rect 25682 18640 25688 18692
rect 25740 18640 25746 18692
rect 29086 18640 29092 18692
rect 29144 18680 29150 18692
rect 30745 18683 30803 18689
rect 30745 18680 30757 18683
rect 29144 18652 30757 18680
rect 29144 18640 29150 18652
rect 30745 18649 30757 18652
rect 30791 18680 30803 18683
rect 30926 18680 30932 18692
rect 30791 18652 30932 18680
rect 30791 18649 30803 18652
rect 30745 18643 30803 18649
rect 30926 18640 30932 18652
rect 30984 18640 30990 18692
rect 29638 18612 29644 18624
rect 25608 18584 29644 18612
rect 24121 18575 24179 18581
rect 29638 18572 29644 18584
rect 29696 18572 29702 18624
rect 29730 18572 29736 18624
rect 29788 18572 29794 18624
rect 30098 18572 30104 18624
rect 30156 18572 30162 18624
rect 43438 18572 43444 18624
rect 43496 18612 43502 18624
rect 48498 18612 48504 18624
rect 43496 18584 48504 18612
rect 43496 18572 43502 18584
rect 48498 18572 48504 18584
rect 48556 18572 48562 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 2240 18380 6500 18408
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2240 18272 2268 18380
rect 5902 18340 5908 18352
rect 3620 18312 5908 18340
rect 3620 18281 3648 18312
rect 5902 18300 5908 18312
rect 5960 18300 5966 18352
rect 1811 18244 2268 18272
rect 3605 18275 3663 18281
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 5626 18232 5632 18284
rect 5684 18232 5690 18284
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 3694 18164 3700 18216
rect 3752 18204 3758 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3752 18176 3893 18204
rect 3752 18164 3758 18176
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 5350 18204 5356 18216
rect 3881 18167 3939 18173
rect 4908 18176 5356 18204
rect 3418 18096 3424 18148
rect 3476 18136 3482 18148
rect 4908 18136 4936 18176
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 5718 18164 5724 18216
rect 5776 18164 5782 18216
rect 5902 18164 5908 18216
rect 5960 18204 5966 18216
rect 6362 18204 6368 18216
rect 5960 18176 6368 18204
rect 5960 18164 5966 18176
rect 6362 18164 6368 18176
rect 6420 18164 6426 18216
rect 6472 18204 6500 18380
rect 6748 18380 13584 18408
rect 6748 18281 6776 18380
rect 7742 18300 7748 18352
rect 7800 18300 7806 18352
rect 12802 18340 12808 18352
rect 9876 18312 12808 18340
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 8444 18244 8493 18272
rect 8444 18232 8450 18244
rect 8481 18241 8493 18244
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8294 18204 8300 18216
rect 6472 18176 8300 18204
rect 8294 18164 8300 18176
rect 8352 18164 8358 18216
rect 8496 18204 8524 18235
rect 8570 18232 8576 18284
rect 8628 18272 8634 18284
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 8628 18244 9229 18272
rect 8628 18232 8634 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9876 18213 9904 18312
rect 12802 18300 12808 18312
rect 12860 18340 12866 18352
rect 13556 18340 13584 18380
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 13780 18380 15393 18408
rect 13780 18368 13786 18380
rect 15381 18377 15393 18380
rect 15427 18377 15439 18411
rect 15381 18371 15439 18377
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 16666 18408 16672 18420
rect 16347 18380 16672 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 17313 18411 17371 18417
rect 17313 18377 17325 18411
rect 17359 18408 17371 18411
rect 20717 18411 20775 18417
rect 20717 18408 20729 18411
rect 17359 18380 20729 18408
rect 17359 18377 17371 18380
rect 17313 18371 17371 18377
rect 20717 18377 20729 18380
rect 20763 18377 20775 18411
rect 20717 18371 20775 18377
rect 21082 18368 21088 18420
rect 21140 18368 21146 18420
rect 21174 18368 21180 18420
rect 21232 18408 21238 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 21232 18380 24869 18408
rect 21232 18368 21238 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 26694 18408 26700 18420
rect 24857 18371 24915 18377
rect 24964 18380 26700 18408
rect 14461 18343 14519 18349
rect 12860 18312 13216 18340
rect 13556 18312 13768 18340
rect 12860 18300 12866 18312
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10008 18244 10793 18272
rect 10008 18232 10014 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18272 11759 18275
rect 12066 18272 12072 18284
rect 11747 18244 12072 18272
rect 11747 18241 11759 18244
rect 11701 18235 11759 18241
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12618 18272 12624 18284
rect 12345 18235 12403 18241
rect 12452 18244 12624 18272
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 8496 18176 9873 18204
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 9861 18167 9919 18173
rect 9968 18176 10885 18204
rect 3476 18108 4936 18136
rect 3476 18096 3482 18108
rect 4982 18096 4988 18148
rect 5040 18136 5046 18148
rect 6638 18136 6644 18148
rect 5040 18108 6644 18136
rect 5040 18096 5046 18108
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 7558 18096 7564 18148
rect 7616 18136 7622 18148
rect 9122 18136 9128 18148
rect 7616 18108 9128 18136
rect 7616 18096 7622 18108
rect 9122 18096 9128 18108
rect 9180 18136 9186 18148
rect 9180 18108 9444 18136
rect 9180 18096 9186 18108
rect 5261 18071 5319 18077
rect 5261 18037 5273 18071
rect 5307 18068 5319 18071
rect 6730 18068 6736 18080
rect 5307 18040 6736 18068
rect 5307 18037 5319 18040
rect 5261 18031 5319 18037
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 8202 18068 8208 18080
rect 7340 18040 8208 18068
rect 7340 18028 7346 18040
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 9306 18068 9312 18080
rect 8352 18040 9312 18068
rect 8352 18028 8358 18040
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 9416 18068 9444 18108
rect 9490 18096 9496 18148
rect 9548 18136 9554 18148
rect 9968 18136 9996 18176
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 11057 18207 11115 18213
rect 11057 18173 11069 18207
rect 11103 18204 11115 18207
rect 11422 18204 11428 18216
rect 11103 18176 11428 18204
rect 11103 18173 11115 18176
rect 11057 18167 11115 18173
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 11790 18164 11796 18216
rect 11848 18204 11854 18216
rect 12360 18204 12388 18235
rect 12452 18213 12480 18244
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 13188 18281 13216 18312
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13633 18275 13691 18281
rect 13633 18272 13645 18275
rect 13173 18235 13231 18241
rect 13556 18244 13645 18272
rect 11848 18176 12388 18204
rect 12437 18207 12495 18213
rect 11848 18164 11854 18176
rect 12437 18173 12449 18207
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12529 18207 12587 18213
rect 12529 18173 12541 18207
rect 12575 18173 12587 18207
rect 13188 18204 13216 18235
rect 13556 18204 13584 18244
rect 13633 18241 13645 18244
rect 13679 18241 13691 18275
rect 13740 18272 13768 18312
rect 14461 18309 14473 18343
rect 14507 18340 14519 18343
rect 14550 18340 14556 18352
rect 14507 18312 14556 18340
rect 14507 18309 14519 18312
rect 14461 18303 14519 18309
rect 14550 18300 14556 18312
rect 14608 18300 14614 18352
rect 15010 18300 15016 18352
rect 15068 18340 15074 18352
rect 18141 18343 18199 18349
rect 15068 18312 17356 18340
rect 15068 18300 15074 18312
rect 16022 18272 16028 18284
rect 13740 18244 16028 18272
rect 13633 18235 13691 18241
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16482 18232 16488 18284
rect 16540 18232 16546 18284
rect 16666 18232 16672 18284
rect 16724 18272 16730 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16724 18244 17233 18272
rect 16724 18232 16730 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17328 18272 17356 18312
rect 18141 18309 18153 18343
rect 18187 18340 18199 18343
rect 20990 18340 20996 18352
rect 18187 18312 20996 18340
rect 18187 18309 18199 18312
rect 18141 18303 18199 18309
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 21100 18340 21128 18368
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21100 18312 22017 18340
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22005 18303 22063 18309
rect 22557 18343 22615 18349
rect 22557 18309 22569 18343
rect 22603 18340 22615 18343
rect 22830 18340 22836 18352
rect 22603 18312 22836 18340
rect 22603 18309 22615 18312
rect 22557 18303 22615 18309
rect 22830 18300 22836 18312
rect 22888 18300 22894 18352
rect 23382 18340 23388 18352
rect 23124 18312 23388 18340
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 17328 18244 18337 18272
rect 17221 18235 17279 18241
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 19334 18232 19340 18284
rect 19392 18272 19398 18284
rect 19889 18275 19947 18281
rect 19889 18272 19901 18275
rect 19392 18244 19901 18272
rect 19392 18232 19398 18244
rect 19889 18241 19901 18244
rect 19935 18241 19947 18275
rect 19889 18235 19947 18241
rect 15102 18204 15108 18216
rect 13188 18176 15108 18204
rect 12529 18167 12587 18173
rect 9548 18108 9996 18136
rect 10413 18139 10471 18145
rect 9548 18096 9554 18108
rect 10413 18105 10425 18139
rect 10459 18136 10471 18139
rect 10459 18108 12112 18136
rect 10459 18105 10471 18108
rect 10413 18099 10471 18105
rect 9677 18071 9735 18077
rect 9677 18068 9689 18071
rect 9416 18040 9689 18068
rect 9677 18037 9689 18040
rect 9723 18037 9735 18071
rect 9677 18031 9735 18037
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9916 18040 10057 18068
rect 9916 18028 9922 18040
rect 10045 18037 10057 18040
rect 10091 18068 10103 18071
rect 10594 18068 10600 18080
rect 10091 18040 10600 18068
rect 10091 18037 10103 18040
rect 10045 18031 10103 18037
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 11977 18071 12035 18077
rect 11977 18068 11989 18071
rect 11940 18040 11989 18068
rect 11940 18028 11946 18040
rect 11977 18037 11989 18040
rect 12023 18037 12035 18071
rect 12084 18068 12112 18108
rect 12250 18096 12256 18148
rect 12308 18136 12314 18148
rect 12544 18136 12572 18167
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16942 18204 16948 18216
rect 15703 18176 16948 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 12308 18108 12572 18136
rect 12308 18096 12314 18108
rect 15010 18096 15016 18148
rect 15068 18096 15074 18148
rect 15488 18136 15516 18167
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17494 18164 17500 18216
rect 17552 18164 17558 18216
rect 18874 18164 18880 18216
rect 18932 18164 18938 18216
rect 19521 18139 19579 18145
rect 19521 18136 19533 18139
rect 15488 18108 19533 18136
rect 19521 18105 19533 18108
rect 19567 18105 19579 18139
rect 19904 18136 19932 18235
rect 19978 18232 19984 18284
rect 20036 18232 20042 18284
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18272 21143 18275
rect 21131 18244 21588 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 20070 18164 20076 18216
rect 20128 18164 20134 18216
rect 20990 18164 20996 18216
rect 21048 18204 21054 18216
rect 21177 18207 21235 18213
rect 21177 18204 21189 18207
rect 21048 18176 21189 18204
rect 21048 18164 21054 18176
rect 21177 18173 21189 18176
rect 21223 18173 21235 18207
rect 21177 18167 21235 18173
rect 21361 18207 21419 18213
rect 21361 18173 21373 18207
rect 21407 18173 21419 18207
rect 21560 18204 21588 18244
rect 21726 18232 21732 18284
rect 21784 18272 21790 18284
rect 23124 18272 23152 18312
rect 23382 18300 23388 18312
rect 23440 18340 23446 18352
rect 23842 18340 23848 18352
rect 23440 18312 23848 18340
rect 23440 18300 23446 18312
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 24762 18300 24768 18352
rect 24820 18340 24826 18352
rect 24964 18340 24992 18380
rect 26694 18368 26700 18380
rect 26752 18368 26758 18420
rect 27157 18411 27215 18417
rect 27157 18377 27169 18411
rect 27203 18408 27215 18411
rect 30098 18408 30104 18420
rect 27203 18380 30104 18408
rect 27203 18377 27215 18380
rect 27157 18371 27215 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 30466 18368 30472 18420
rect 30524 18408 30530 18420
rect 30653 18411 30711 18417
rect 30653 18408 30665 18411
rect 30524 18380 30665 18408
rect 30524 18368 30530 18380
rect 30653 18377 30665 18380
rect 30699 18408 30711 18411
rect 31297 18411 31355 18417
rect 31297 18408 31309 18411
rect 30699 18380 31309 18408
rect 30699 18377 30711 18380
rect 30653 18371 30711 18377
rect 31297 18377 31309 18380
rect 31343 18408 31355 18411
rect 31343 18380 31754 18408
rect 31343 18377 31355 18380
rect 31297 18371 31355 18377
rect 24820 18312 24992 18340
rect 24820 18300 24826 18312
rect 25314 18300 25320 18352
rect 25372 18300 25378 18352
rect 26050 18300 26056 18352
rect 26108 18300 26114 18352
rect 28353 18343 28411 18349
rect 28353 18309 28365 18343
rect 28399 18340 28411 18343
rect 28626 18340 28632 18352
rect 28399 18312 28632 18340
rect 28399 18309 28411 18312
rect 28353 18303 28411 18309
rect 28626 18300 28632 18312
rect 28684 18300 28690 18352
rect 29086 18300 29092 18352
rect 29144 18300 29150 18352
rect 31726 18340 31754 18380
rect 43346 18340 43352 18352
rect 31726 18312 43352 18340
rect 43346 18300 43352 18312
rect 43404 18300 43410 18352
rect 21784 18244 23152 18272
rect 25332 18272 25360 18300
rect 26513 18275 26571 18281
rect 26513 18272 26525 18275
rect 25332 18244 26525 18272
rect 21784 18232 21790 18244
rect 26513 18241 26525 18244
rect 26559 18241 26571 18275
rect 26513 18235 26571 18241
rect 27798 18232 27804 18284
rect 27856 18272 27862 18284
rect 28077 18275 28135 18281
rect 28077 18272 28089 18275
rect 27856 18244 28089 18272
rect 27856 18232 27862 18244
rect 28077 18241 28089 18244
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 29638 18232 29644 18284
rect 29696 18272 29702 18284
rect 30745 18275 30803 18281
rect 30745 18272 30757 18275
rect 29696 18244 30757 18272
rect 29696 18232 29702 18244
rect 30745 18241 30757 18244
rect 30791 18272 30803 18275
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 30791 18244 31493 18272
rect 30791 18241 30803 18244
rect 30745 18235 30803 18241
rect 31481 18241 31493 18244
rect 31527 18272 31539 18275
rect 31527 18244 35894 18272
rect 31527 18241 31539 18244
rect 31481 18235 31539 18241
rect 22830 18204 22836 18216
rect 21560 18176 22836 18204
rect 21361 18167 21419 18173
rect 19978 18136 19984 18148
rect 19904 18108 19984 18136
rect 19521 18099 19579 18105
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 12710 18068 12716 18080
rect 12084 18040 12716 18068
rect 11977 18031 12035 18037
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 13354 18028 13360 18080
rect 13412 18028 13418 18080
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 15654 18068 15660 18080
rect 14608 18040 15660 18068
rect 14608 18028 14614 18040
rect 15654 18028 15660 18040
rect 15712 18068 15718 18080
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15712 18040 16037 18068
rect 15712 18028 15718 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 16853 18071 16911 18077
rect 16853 18037 16865 18071
rect 16899 18068 16911 18071
rect 17862 18068 17868 18080
rect 16899 18040 17868 18068
rect 16899 18037 16911 18040
rect 16853 18031 16911 18037
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 21376 18068 21404 18167
rect 22830 18164 22836 18176
rect 22888 18164 22894 18216
rect 23109 18207 23167 18213
rect 23109 18173 23121 18207
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 26234 18204 26240 18216
rect 23431 18176 26240 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 18380 18040 21404 18068
rect 23124 18068 23152 18167
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 27062 18164 27068 18216
rect 27120 18204 27126 18216
rect 30837 18207 30895 18213
rect 27120 18176 30328 18204
rect 27120 18164 27126 18176
rect 30300 18145 30328 18176
rect 30837 18173 30849 18207
rect 30883 18173 30895 18207
rect 35866 18204 35894 18244
rect 45002 18204 45008 18216
rect 35866 18176 45008 18204
rect 30837 18167 30895 18173
rect 30285 18139 30343 18145
rect 30285 18105 30297 18139
rect 30331 18105 30343 18139
rect 30285 18099 30343 18105
rect 30374 18096 30380 18148
rect 30432 18136 30438 18148
rect 30852 18136 30880 18167
rect 45002 18164 45008 18176
rect 45060 18164 45066 18216
rect 39574 18136 39580 18148
rect 30432 18108 39580 18136
rect 30432 18096 30438 18108
rect 39574 18096 39580 18108
rect 39632 18096 39638 18148
rect 24670 18068 24676 18080
rect 23124 18040 24676 18068
rect 18380 18028 18386 18040
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 26694 18028 26700 18080
rect 26752 18028 26758 18080
rect 27338 18028 27344 18080
rect 27396 18068 27402 18080
rect 29822 18068 29828 18080
rect 27396 18040 29828 18068
rect 27396 18028 27402 18040
rect 29822 18028 29828 18040
rect 29880 18028 29886 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 3605 17867 3663 17873
rect 3605 17833 3617 17867
rect 3651 17864 3663 17867
rect 8386 17864 8392 17876
rect 3651 17836 8392 17864
rect 3651 17833 3663 17836
rect 3605 17827 3663 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 8570 17824 8576 17876
rect 8628 17864 8634 17876
rect 9398 17864 9404 17876
rect 8628 17836 9404 17864
rect 8628 17824 8634 17836
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 10376 17836 10609 17864
rect 10376 17824 10382 17836
rect 10597 17833 10609 17836
rect 10643 17833 10655 17867
rect 16114 17864 16120 17876
rect 10597 17827 10655 17833
rect 10704 17836 16120 17864
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 4433 17799 4491 17805
rect 4433 17796 4445 17799
rect 1912 17768 4445 17796
rect 1912 17756 1918 17768
rect 4433 17765 4445 17768
rect 4479 17765 4491 17799
rect 4433 17759 4491 17765
rect 6638 17756 6644 17808
rect 6696 17756 6702 17808
rect 7098 17756 7104 17808
rect 7156 17796 7162 17808
rect 7156 17768 7788 17796
rect 7156 17756 7162 17768
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 1780 17700 7389 17728
rect 1780 17669 1808 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7760 17728 7788 17768
rect 7834 17756 7840 17808
rect 7892 17756 7898 17808
rect 8404 17796 8432 17824
rect 10704 17796 10732 17836
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 16758 17864 16764 17876
rect 16408 17836 16764 17864
rect 8404 17768 9168 17796
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7760 17700 8401 17728
rect 7377 17691 7435 17697
rect 8389 17697 8401 17700
rect 8435 17728 8447 17731
rect 9030 17728 9036 17740
rect 8435 17700 9036 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 9140 17672 9168 17768
rect 9232 17768 10732 17796
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17629 1823 17663
rect 1765 17623 1823 17629
rect 3602 17620 3608 17672
rect 3660 17660 3666 17672
rect 3878 17660 3884 17672
rect 3660 17632 3884 17660
rect 3660 17620 3666 17632
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4614 17660 4620 17672
rect 4212 17632 4620 17660
rect 4212 17620 4218 17632
rect 4614 17620 4620 17632
rect 4672 17660 4678 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4672 17632 4905 17660
rect 4672 17620 4678 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 8202 17620 8208 17672
rect 8260 17620 8266 17672
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 1210 17552 1216 17604
rect 1268 17592 1274 17604
rect 2501 17595 2559 17601
rect 2501 17592 2513 17595
rect 1268 17564 2513 17592
rect 1268 17552 1274 17564
rect 2501 17561 2513 17564
rect 2547 17561 2559 17595
rect 2501 17555 2559 17561
rect 4246 17552 4252 17604
rect 4304 17552 4310 17604
rect 5169 17595 5227 17601
rect 5169 17561 5181 17595
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 3418 17484 3424 17536
rect 3476 17484 3482 17536
rect 3786 17484 3792 17536
rect 3844 17484 3850 17536
rect 5184 17524 5212 17555
rect 6178 17552 6184 17604
rect 6236 17552 6242 17604
rect 7193 17595 7251 17601
rect 7193 17561 7205 17595
rect 7239 17592 7251 17595
rect 7282 17592 7288 17604
rect 7239 17564 7288 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 7282 17552 7288 17564
rect 7340 17552 7346 17604
rect 8297 17595 8355 17601
rect 8297 17561 8309 17595
rect 8343 17592 8355 17595
rect 8570 17592 8576 17604
rect 8343 17564 8576 17592
rect 8343 17561 8355 17564
rect 8297 17555 8355 17561
rect 8570 17552 8576 17564
rect 8628 17552 8634 17604
rect 7466 17524 7472 17536
rect 5184 17496 7472 17524
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 9232 17524 9260 17768
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 11882 17796 11888 17808
rect 10928 17768 11888 17796
rect 10928 17756 10934 17768
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 13630 17756 13636 17808
rect 13688 17796 13694 17808
rect 13725 17799 13783 17805
rect 13725 17796 13737 17799
rect 13688 17768 13737 17796
rect 13688 17756 13694 17768
rect 13725 17765 13737 17768
rect 13771 17765 13783 17799
rect 13725 17759 13783 17765
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 16025 17799 16083 17805
rect 16025 17796 16037 17799
rect 15344 17768 16037 17796
rect 15344 17756 15350 17768
rect 16025 17765 16037 17768
rect 16071 17796 16083 17799
rect 16408 17796 16436 17836
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17184 17836 23612 17864
rect 17184 17824 17190 17836
rect 16071 17768 16436 17796
rect 16071 17765 16083 17768
rect 16025 17759 16083 17765
rect 17678 17756 17684 17808
rect 17736 17796 17742 17808
rect 17736 17768 19748 17796
rect 17736 17756 17742 17768
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9732 17700 9873 17728
rect 9732 17688 9738 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10134 17688 10140 17740
rect 10192 17728 10198 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10192 17700 11161 17728
rect 10192 17688 10198 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 14366 17728 14372 17740
rect 11149 17691 11207 17697
rect 11716 17700 14372 17728
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11716 17660 11744 17700
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 16298 17688 16304 17740
rect 16356 17688 16362 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16942 17728 16948 17740
rect 16623 17700 16948 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 17034 17688 17040 17740
rect 17092 17728 17098 17740
rect 19720 17737 19748 17768
rect 20070 17756 20076 17808
rect 20128 17796 20134 17808
rect 21818 17796 21824 17808
rect 20128 17768 21824 17796
rect 20128 17756 20134 17768
rect 21818 17756 21824 17768
rect 21876 17756 21882 17808
rect 23584 17796 23612 17836
rect 26234 17824 26240 17876
rect 26292 17864 26298 17876
rect 27338 17873 27344 17876
rect 26605 17867 26663 17873
rect 26605 17864 26617 17867
rect 26292 17836 26617 17864
rect 26292 17824 26298 17836
rect 26605 17833 26617 17836
rect 26651 17833 26663 17867
rect 26605 17827 26663 17833
rect 27322 17867 27344 17873
rect 27322 17833 27334 17867
rect 27322 17827 27344 17833
rect 27338 17824 27344 17827
rect 27396 17824 27402 17876
rect 27430 17824 27436 17876
rect 27488 17864 27494 17876
rect 28994 17864 29000 17876
rect 27488 17836 29000 17864
rect 27488 17824 27494 17836
rect 28994 17824 29000 17836
rect 29052 17824 29058 17876
rect 29086 17824 29092 17876
rect 29144 17824 29150 17876
rect 31938 17824 31944 17876
rect 31996 17824 32002 17876
rect 24302 17796 24308 17808
rect 23584 17768 24308 17796
rect 24302 17756 24308 17768
rect 24360 17756 24366 17808
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 29733 17799 29791 17805
rect 29733 17796 29745 17799
rect 28500 17768 29745 17796
rect 28500 17756 28506 17768
rect 29733 17765 29745 17768
rect 29779 17765 29791 17799
rect 30374 17796 30380 17808
rect 29733 17759 29791 17765
rect 30300 17768 30380 17796
rect 19429 17731 19487 17737
rect 19429 17728 19441 17731
rect 17092 17700 19441 17728
rect 17092 17688 17098 17700
rect 19429 17697 19441 17700
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 20438 17688 20444 17740
rect 20496 17728 20502 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 20496 17700 21281 17728
rect 20496 17688 20502 17700
rect 21269 17697 21281 17700
rect 21315 17728 21327 17731
rect 24486 17728 24492 17740
rect 21315 17700 24492 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 24486 17688 24492 17700
rect 24544 17688 24550 17740
rect 24670 17688 24676 17740
rect 24728 17728 24734 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24728 17700 24869 17728
rect 24728 17688 24734 17700
rect 24857 17697 24869 17700
rect 24903 17728 24915 17731
rect 25774 17728 25780 17740
rect 24903 17700 25780 17728
rect 24903 17697 24915 17700
rect 24857 17691 24915 17697
rect 25774 17688 25780 17700
rect 25832 17728 25838 17740
rect 27065 17731 27123 17737
rect 27065 17728 27077 17731
rect 25832 17700 27077 17728
rect 25832 17688 25838 17700
rect 27065 17697 27077 17700
rect 27111 17728 27123 17731
rect 27798 17728 27804 17740
rect 27111 17700 27804 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 27798 17688 27804 17700
rect 27856 17688 27862 17740
rect 30190 17688 30196 17740
rect 30248 17688 30254 17740
rect 30300 17737 30328 17768
rect 30374 17756 30380 17768
rect 30432 17756 30438 17808
rect 30285 17731 30343 17737
rect 30285 17697 30297 17731
rect 30331 17697 30343 17731
rect 31481 17731 31539 17737
rect 31481 17728 31493 17731
rect 30285 17691 30343 17697
rect 30852 17700 31493 17728
rect 11011 17632 11744 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 13354 17620 13360 17672
rect 13412 17620 13418 17672
rect 14918 17660 14924 17672
rect 13648 17632 14924 17660
rect 9398 17552 9404 17604
rect 9456 17592 9462 17604
rect 11057 17595 11115 17601
rect 11057 17592 11069 17595
rect 9456 17564 11069 17592
rect 9456 17552 9462 17564
rect 11057 17561 11069 17564
rect 11103 17561 11115 17595
rect 12158 17592 12164 17604
rect 11057 17555 11115 17561
rect 11256 17564 12164 17592
rect 7616 17496 9260 17524
rect 7616 17484 7622 17496
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 11256 17524 11284 17564
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 12250 17552 12256 17604
rect 12308 17552 12314 17604
rect 10376 17496 11284 17524
rect 10376 17484 10382 17496
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 11609 17527 11667 17533
rect 11609 17524 11621 17527
rect 11388 17496 11621 17524
rect 11388 17484 11394 17496
rect 11609 17493 11621 17496
rect 11655 17493 11667 17527
rect 11609 17487 11667 17493
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 13648 17524 13676 17632
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 15378 17620 15384 17672
rect 15436 17620 15442 17672
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 17736 17632 18337 17660
rect 17736 17620 17742 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21726 17660 21732 17672
rect 20956 17632 21732 17660
rect 20956 17620 20962 17632
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 22002 17620 22008 17672
rect 22060 17660 22066 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22060 17632 22293 17660
rect 22060 17620 22066 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 22281 17623 22339 17629
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17592 14427 17595
rect 15396 17592 15424 17620
rect 16298 17592 16304 17604
rect 14415 17564 14964 17592
rect 15396 17564 16304 17592
rect 14415 17561 14427 17564
rect 14369 17555 14427 17561
rect 14936 17536 14964 17564
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 17880 17564 18828 17592
rect 11940 17496 13676 17524
rect 11940 17484 11946 17496
rect 14458 17484 14464 17536
rect 14516 17484 14522 17536
rect 14918 17484 14924 17536
rect 14976 17484 14982 17536
rect 15102 17484 15108 17536
rect 15160 17484 15166 17536
rect 15378 17484 15384 17536
rect 15436 17484 15442 17536
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 17880 17524 17908 17564
rect 16448 17496 17908 17524
rect 18049 17527 18107 17533
rect 16448 17484 16454 17496
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18322 17524 18328 17536
rect 18095 17496 18328 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 18690 17484 18696 17536
rect 18748 17484 18754 17536
rect 18800 17524 18828 17564
rect 18874 17552 18880 17604
rect 18932 17592 18938 17604
rect 21085 17595 21143 17601
rect 21085 17592 21097 17595
rect 18932 17564 21097 17592
rect 18932 17552 18938 17564
rect 21085 17561 21097 17564
rect 21131 17561 21143 17595
rect 21085 17555 21143 17561
rect 21266 17552 21272 17604
rect 21324 17592 21330 17604
rect 22557 17595 22615 17601
rect 22557 17592 22569 17595
rect 21324 17564 22569 17592
rect 21324 17552 21330 17564
rect 22557 17561 22569 17564
rect 22603 17561 22615 17595
rect 22557 17555 22615 17561
rect 23198 17552 23204 17604
rect 23256 17552 23262 17604
rect 25133 17595 25191 17601
rect 25133 17592 25145 17595
rect 24044 17564 25145 17592
rect 20717 17527 20775 17533
rect 20717 17524 20729 17527
rect 18800 17496 20729 17524
rect 20717 17493 20729 17496
rect 20763 17493 20775 17527
rect 20717 17487 20775 17493
rect 21174 17484 21180 17536
rect 21232 17484 21238 17536
rect 21634 17484 21640 17536
rect 21692 17524 21698 17536
rect 24044 17533 24072 17564
rect 25133 17561 25145 17564
rect 25179 17592 25191 17595
rect 25406 17592 25412 17604
rect 25179 17564 25412 17592
rect 25179 17561 25191 17564
rect 25133 17555 25191 17561
rect 25406 17552 25412 17564
rect 25464 17552 25470 17604
rect 26694 17592 26700 17604
rect 26358 17564 26700 17592
rect 26694 17552 26700 17564
rect 26752 17592 26758 17604
rect 30101 17595 30159 17601
rect 30101 17592 30113 17595
rect 26752 17564 27830 17592
rect 28644 17564 30113 17592
rect 26752 17552 26758 17564
rect 21913 17527 21971 17533
rect 21913 17524 21925 17527
rect 21692 17496 21925 17524
rect 21692 17484 21698 17496
rect 21913 17493 21925 17496
rect 21959 17493 21971 17527
rect 21913 17487 21971 17493
rect 24029 17527 24087 17533
rect 24029 17493 24041 17527
rect 24075 17493 24087 17527
rect 24029 17487 24087 17493
rect 24394 17484 24400 17536
rect 24452 17524 24458 17536
rect 28644 17524 28672 17564
rect 30101 17561 30113 17564
rect 30147 17592 30159 17595
rect 30742 17592 30748 17604
rect 30147 17564 30748 17592
rect 30147 17561 30159 17564
rect 30101 17555 30159 17561
rect 30742 17552 30748 17564
rect 30800 17552 30806 17604
rect 24452 17496 28672 17524
rect 24452 17484 24458 17496
rect 28810 17484 28816 17536
rect 28868 17524 28874 17536
rect 30852 17524 30880 17700
rect 31481 17697 31493 17700
rect 31527 17697 31539 17731
rect 31481 17691 31539 17697
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17660 31355 17663
rect 31938 17660 31944 17672
rect 31343 17632 31944 17660
rect 31343 17629 31355 17632
rect 31297 17623 31355 17629
rect 31938 17620 31944 17632
rect 31996 17620 32002 17672
rect 31389 17595 31447 17601
rect 31389 17561 31401 17595
rect 31435 17592 31447 17595
rect 37550 17592 37556 17604
rect 31435 17564 37556 17592
rect 31435 17561 31447 17564
rect 31389 17555 31447 17561
rect 37550 17552 37556 17564
rect 37608 17552 37614 17604
rect 28868 17496 30880 17524
rect 28868 17484 28874 17496
rect 30926 17484 30932 17536
rect 30984 17484 30990 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 5261 17323 5319 17329
rect 2746 17292 4568 17320
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2746 17184 2774 17292
rect 4430 17212 4436 17264
rect 4488 17212 4494 17264
rect 4540 17252 4568 17292
rect 5261 17289 5273 17323
rect 5307 17320 5319 17323
rect 7285 17323 7343 17329
rect 7285 17320 7297 17323
rect 5307 17292 7297 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 7285 17289 7297 17292
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7432 17292 8033 17320
rect 7432 17280 7438 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 8481 17323 8539 17329
rect 8481 17289 8493 17323
rect 8527 17320 8539 17323
rect 8570 17320 8576 17332
rect 8527 17292 8576 17320
rect 8527 17289 8539 17292
rect 8481 17283 8539 17289
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 9582 17320 9588 17332
rect 9539 17292 9588 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 9953 17323 10011 17329
rect 9953 17289 9965 17323
rect 9999 17320 10011 17323
rect 10410 17320 10416 17332
rect 9999 17292 10416 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 11664 17292 12541 17320
rect 11664 17280 11670 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 12897 17323 12955 17329
rect 12897 17320 12909 17323
rect 12529 17283 12587 17289
rect 12636 17292 12909 17320
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 4540 17224 10977 17252
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 1811 17156 2774 17184
rect 3605 17187 3663 17193
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 3651 17156 5304 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 5276 16980 5304 17156
rect 5350 17144 5356 17196
rect 5408 17184 5414 17196
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5408 17156 5641 17184
rect 5408 17144 5414 17156
rect 5629 17153 5641 17156
rect 5675 17153 5687 17187
rect 6086 17184 6092 17196
rect 5629 17147 5687 17153
rect 5828 17156 6092 17184
rect 5828 17125 5856 17156
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6454 17144 6460 17196
rect 6512 17144 6518 17196
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17184 7251 17187
rect 7834 17184 7840 17196
rect 7239 17156 7840 17184
rect 7239 17153 7251 17156
rect 7193 17147 7251 17153
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 8386 17144 8392 17196
rect 8444 17144 8450 17196
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 8496 17156 9137 17184
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 6472 17116 6500 17144
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 6472 17088 7389 17116
rect 5813 17079 5871 17085
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 5736 17048 5764 17079
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 8496 17116 8524 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 7984 17088 8524 17116
rect 8665 17119 8723 17125
rect 7984 17076 7990 17088
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 8846 17116 8852 17128
rect 8711 17088 8852 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 9140 17116 9168 17147
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 10318 17184 10324 17196
rect 9968 17156 10324 17184
rect 9766 17116 9772 17128
rect 9140 17088 9772 17116
rect 9766 17076 9772 17088
rect 9824 17116 9830 17128
rect 9968 17116 9996 17156
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 10778 17144 10784 17196
rect 10836 17144 10842 17196
rect 11330 17144 11336 17196
rect 11388 17184 11394 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11388 17156 11805 17184
rect 11388 17144 11394 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12636 17184 12664 17292
rect 12897 17289 12909 17292
rect 12943 17289 12955 17323
rect 12897 17283 12955 17289
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 13630 17320 13636 17332
rect 13136 17292 13636 17320
rect 13136 17280 13142 17292
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 13722 17280 13728 17332
rect 13780 17280 13786 17332
rect 15013 17323 15071 17329
rect 15013 17289 15025 17323
rect 15059 17320 15071 17323
rect 15059 17292 21404 17320
rect 15059 17289 15071 17292
rect 15013 17283 15071 17289
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 15028 17252 15056 17283
rect 13035 17224 15056 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 18322 17212 18328 17264
rect 18380 17252 18386 17264
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 18380 17224 18429 17252
rect 18380 17212 18386 17224
rect 18417 17221 18429 17224
rect 18463 17221 18475 17255
rect 18417 17215 18475 17221
rect 20070 17212 20076 17264
rect 20128 17252 20134 17264
rect 20349 17255 20407 17261
rect 20349 17252 20361 17255
rect 20128 17224 20361 17252
rect 20128 17212 20134 17224
rect 20349 17221 20361 17224
rect 20395 17252 20407 17255
rect 20395 17224 21036 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 12584 17156 12664 17184
rect 12584 17144 12590 17156
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13504 17156 14105 17184
rect 13504 17144 13510 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17184 15255 17187
rect 15286 17184 15292 17196
rect 15243 17156 15292 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 17126 17184 17132 17196
rect 16347 17156 17132 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 17218 17144 17224 17196
rect 17276 17144 17282 17196
rect 20162 17184 20168 17196
rect 19550 17156 20168 17184
rect 20162 17144 20168 17156
rect 20220 17184 20226 17196
rect 20898 17184 20904 17196
rect 20220 17156 20904 17184
rect 20220 17144 20226 17156
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 9824 17088 9996 17116
rect 9824 17076 9830 17088
rect 10042 17076 10048 17128
rect 10100 17076 10106 17128
rect 13078 17076 13084 17128
rect 13136 17076 13142 17128
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 14185 17119 14243 17125
rect 14185 17116 14197 17119
rect 13872 17088 14197 17116
rect 13872 17076 13878 17088
rect 14185 17085 14197 17088
rect 14231 17085 14243 17119
rect 14185 17079 14243 17085
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 15470 17116 15476 17128
rect 14415 17088 15476 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 5408 17020 5764 17048
rect 5408 17008 5414 17020
rect 6454 17008 6460 17060
rect 6512 17008 6518 17060
rect 6822 17008 6828 17060
rect 6880 17008 6886 17060
rect 11977 17051 12035 17057
rect 11977 17048 11989 17051
rect 7484 17020 11989 17048
rect 7484 16980 7512 17020
rect 11977 17017 11989 17020
rect 12023 17017 12035 17051
rect 14200 17048 14228 17079
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 15838 17076 15844 17128
rect 15896 17116 15902 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 15896 17088 17325 17116
rect 15896 17076 15902 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 14737 17051 14795 17057
rect 14737 17048 14749 17051
rect 14200 17020 14749 17048
rect 11977 17011 12035 17017
rect 14737 17017 14749 17020
rect 14783 17017 14795 17051
rect 14737 17011 14795 17017
rect 15028 17020 16068 17048
rect 5276 16952 7512 16980
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 10226 16980 10232 16992
rect 9088 16952 10232 16980
rect 9088 16940 9094 16952
rect 10226 16940 10232 16952
rect 10284 16980 10290 16992
rect 10870 16980 10876 16992
rect 10284 16952 10876 16980
rect 10284 16940 10290 16952
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 11333 16983 11391 16989
rect 11333 16949 11345 16983
rect 11379 16980 11391 16983
rect 11698 16980 11704 16992
rect 11379 16952 11704 16980
rect 11379 16949 11391 16952
rect 11333 16943 11391 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 15028 16980 15056 17020
rect 12860 16952 15056 16980
rect 15473 16983 15531 16989
rect 12860 16940 12866 16952
rect 15473 16949 15485 16983
rect 15519 16980 15531 16983
rect 15746 16980 15752 16992
rect 15519 16952 15752 16980
rect 15519 16949 15531 16952
rect 15473 16943 15531 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 16040 16980 16068 17020
rect 16114 17008 16120 17060
rect 16172 17008 16178 17060
rect 17034 17008 17040 17060
rect 17092 17048 17098 17060
rect 18156 17048 18184 17079
rect 19702 17076 19708 17128
rect 19760 17116 19766 17128
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 19760 17088 20269 17116
rect 19760 17076 19766 17088
rect 20257 17085 20269 17088
rect 20303 17116 20315 17119
rect 20622 17116 20628 17128
rect 20303 17088 20628 17116
rect 20303 17085 20315 17088
rect 20257 17079 20315 17085
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 21008 17116 21036 17224
rect 21082 17144 21088 17196
rect 21140 17144 21146 17196
rect 21376 17184 21404 17292
rect 21450 17280 21456 17332
rect 21508 17320 21514 17332
rect 23661 17323 23719 17329
rect 23661 17320 23673 17323
rect 21508 17292 23673 17320
rect 21508 17280 21514 17292
rect 23661 17289 23673 17292
rect 23707 17320 23719 17323
rect 24394 17320 24400 17332
rect 23707 17292 24400 17320
rect 23707 17289 23719 17292
rect 23661 17283 23719 17289
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 24762 17280 24768 17332
rect 24820 17280 24826 17332
rect 28810 17320 28816 17332
rect 24964 17292 28816 17320
rect 21634 17212 21640 17264
rect 21692 17252 21698 17264
rect 22465 17255 22523 17261
rect 22465 17252 22477 17255
rect 21692 17224 22477 17252
rect 21692 17212 21698 17224
rect 22465 17221 22477 17224
rect 22511 17252 22523 17255
rect 23290 17252 23296 17264
rect 22511 17224 23296 17252
rect 22511 17221 22523 17224
rect 22465 17215 22523 17221
rect 23290 17212 23296 17224
rect 23348 17212 23354 17264
rect 23753 17255 23811 17261
rect 23753 17221 23765 17255
rect 23799 17252 23811 17255
rect 24026 17252 24032 17264
rect 23799 17224 24032 17252
rect 23799 17221 23811 17224
rect 23753 17215 23811 17221
rect 24026 17212 24032 17224
rect 24084 17212 24090 17264
rect 24302 17212 24308 17264
rect 24360 17252 24366 17264
rect 24780 17252 24808 17280
rect 24964 17261 24992 17292
rect 28810 17280 28816 17292
rect 28868 17280 28874 17332
rect 29086 17280 29092 17332
rect 29144 17320 29150 17332
rect 29825 17323 29883 17329
rect 29825 17320 29837 17323
rect 29144 17292 29837 17320
rect 29144 17280 29150 17292
rect 29825 17289 29837 17292
rect 29871 17289 29883 17323
rect 29825 17283 29883 17289
rect 30190 17280 30196 17332
rect 30248 17320 30254 17332
rect 30561 17323 30619 17329
rect 30561 17320 30573 17323
rect 30248 17292 30573 17320
rect 30248 17280 30254 17292
rect 30561 17289 30573 17292
rect 30607 17320 30619 17323
rect 36998 17320 37004 17332
rect 30607 17292 37004 17320
rect 30607 17289 30619 17292
rect 30561 17283 30619 17289
rect 36998 17280 37004 17292
rect 37056 17280 37062 17332
rect 24360 17224 24808 17252
rect 24949 17255 25007 17261
rect 24360 17212 24366 17224
rect 24949 17221 24961 17255
rect 24995 17221 25007 17255
rect 26694 17252 26700 17264
rect 26174 17224 26700 17252
rect 24949 17215 25007 17221
rect 26694 17212 26700 17224
rect 26752 17252 26758 17264
rect 26752 17224 28566 17252
rect 26752 17212 26758 17224
rect 30742 17212 30748 17264
rect 30800 17252 30806 17264
rect 30837 17255 30895 17261
rect 30837 17252 30849 17255
rect 30800 17224 30849 17252
rect 30800 17212 30806 17224
rect 30837 17221 30849 17224
rect 30883 17252 30895 17255
rect 30883 17224 31754 17252
rect 30883 17221 30895 17224
rect 30837 17215 30895 17221
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 21376 17156 22385 17184
rect 22373 17153 22385 17156
rect 22419 17184 22431 17187
rect 22830 17184 22836 17196
rect 22419 17156 22836 17184
rect 22419 17153 22431 17156
rect 22373 17147 22431 17153
rect 22830 17144 22836 17156
rect 22888 17144 22894 17196
rect 24670 17144 24676 17196
rect 24728 17144 24734 17196
rect 27798 17144 27804 17196
rect 27856 17144 27862 17196
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 21008 17088 21189 17116
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17085 21419 17119
rect 21361 17079 21419 17085
rect 21266 17048 21272 17060
rect 17092 17020 18184 17048
rect 19904 17020 21272 17048
rect 17092 17008 17098 17020
rect 16758 16980 16764 16992
rect 16040 16952 16764 16980
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 16850 16940 16856 16992
rect 16908 16940 16914 16992
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 19904 16989 19932 17020
rect 21266 17008 21272 17020
rect 21324 17008 21330 17060
rect 21376 17048 21404 17079
rect 21634 17076 21640 17128
rect 21692 17116 21698 17128
rect 22557 17119 22615 17125
rect 22557 17116 22569 17119
rect 21692 17088 22569 17116
rect 21692 17076 21698 17088
rect 22557 17085 22569 17088
rect 22603 17085 22615 17119
rect 22557 17079 22615 17085
rect 23845 17119 23903 17125
rect 23845 17085 23857 17119
rect 23891 17085 23903 17119
rect 23845 17079 23903 17085
rect 23860 17048 23888 17079
rect 24486 17076 24492 17128
rect 24544 17116 24550 17128
rect 26421 17119 26479 17125
rect 26421 17116 26433 17119
rect 24544 17088 26433 17116
rect 24544 17076 24550 17088
rect 26421 17085 26433 17088
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27706 17116 27712 17128
rect 27203 17088 27712 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 27706 17076 27712 17088
rect 27764 17076 27770 17128
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17116 28135 17119
rect 30374 17116 30380 17128
rect 28123 17088 30380 17116
rect 28123 17085 28135 17088
rect 28077 17079 28135 17085
rect 30374 17076 30380 17088
rect 30432 17076 30438 17128
rect 21376 17020 22232 17048
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 17552 16952 19901 16980
rect 17552 16940 17558 16952
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 20714 16940 20720 16992
rect 20772 16940 20778 16992
rect 20806 16940 20812 16992
rect 20864 16980 20870 16992
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 20864 16952 22017 16980
rect 20864 16940 20870 16952
rect 22005 16949 22017 16952
rect 22051 16949 22063 16983
rect 22204 16980 22232 17020
rect 22664 17020 23888 17048
rect 22664 16992 22692 17020
rect 22646 16980 22652 16992
rect 22204 16952 22652 16980
rect 22005 16943 22063 16949
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 23290 16940 23296 16992
rect 23348 16940 23354 16992
rect 24670 16940 24676 16992
rect 24728 16980 24734 16992
rect 25130 16980 25136 16992
rect 24728 16952 25136 16980
rect 24728 16940 24734 16952
rect 25130 16940 25136 16952
rect 25188 16940 25194 16992
rect 26694 16940 26700 16992
rect 26752 16940 26758 16992
rect 27154 16940 27160 16992
rect 27212 16980 27218 16992
rect 29549 16983 29607 16989
rect 29549 16980 29561 16983
rect 27212 16952 29561 16980
rect 27212 16940 27218 16952
rect 29549 16949 29561 16952
rect 29595 16949 29607 16983
rect 31726 16980 31754 17224
rect 42794 16980 42800 16992
rect 31726 16952 42800 16980
rect 29549 16943 29607 16949
rect 42794 16940 42800 16952
rect 42852 16940 42858 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 842 16736 848 16788
rect 900 16776 906 16788
rect 1118 16776 1124 16788
rect 900 16748 1124 16776
rect 900 16736 906 16748
rect 1118 16736 1124 16748
rect 1176 16736 1182 16788
rect 3602 16736 3608 16788
rect 3660 16736 3666 16788
rect 3970 16736 3976 16788
rect 4028 16776 4034 16788
rect 5350 16776 5356 16788
rect 4028 16748 5356 16776
rect 4028 16736 4034 16748
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 5810 16736 5816 16788
rect 5868 16776 5874 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5868 16748 6009 16776
rect 5868 16736 5874 16748
rect 5997 16745 6009 16748
rect 6043 16745 6055 16779
rect 7558 16776 7564 16788
rect 5997 16739 6055 16745
rect 6104 16748 7564 16776
rect 4246 16668 4252 16720
rect 4304 16708 4310 16720
rect 6104 16708 6132 16748
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 7760 16748 7972 16776
rect 4304 16680 6132 16708
rect 4304 16668 4310 16680
rect 566 16600 572 16652
rect 624 16640 630 16652
rect 842 16640 848 16652
rect 624 16612 848 16640
rect 624 16600 630 16612
rect 842 16600 848 16612
rect 900 16600 906 16652
rect 2222 16600 2228 16652
rect 2280 16640 2286 16652
rect 3329 16643 3387 16649
rect 3329 16640 3341 16643
rect 2280 16612 3341 16640
rect 2280 16600 2286 16612
rect 3329 16609 3341 16612
rect 3375 16640 3387 16643
rect 5902 16640 5908 16652
rect 3375 16612 5908 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 5994 16600 6000 16652
rect 6052 16640 6058 16652
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 6052 16612 7113 16640
rect 6052 16600 6058 16612
rect 7101 16609 7113 16612
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 7760 16640 7788 16748
rect 7944 16708 7972 16748
rect 8110 16736 8116 16788
rect 8168 16776 8174 16788
rect 11606 16776 11612 16788
rect 8168 16748 11612 16776
rect 8168 16736 8174 16748
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 12526 16776 12532 16788
rect 12176 16748 12532 16776
rect 7944 16680 8524 16708
rect 7331 16612 7788 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 8496 16649 8524 16680
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 9490 16708 9496 16720
rect 8628 16680 9496 16708
rect 8628 16668 8634 16680
rect 9490 16668 9496 16680
rect 9548 16708 9554 16720
rect 9766 16708 9772 16720
rect 9548 16680 9772 16708
rect 9548 16668 9554 16680
rect 9766 16668 9772 16680
rect 9824 16668 9830 16720
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 10045 16711 10103 16717
rect 10045 16708 10057 16711
rect 9916 16680 10057 16708
rect 9916 16668 9922 16680
rect 10045 16677 10057 16680
rect 10091 16677 10103 16711
rect 10045 16671 10103 16677
rect 10336 16680 10732 16708
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 8168 16612 8309 16640
rect 8168 16600 8174 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 10336 16640 10364 16680
rect 8527 16612 10364 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 10704 16649 10732 16680
rect 10870 16668 10876 16720
rect 10928 16708 10934 16720
rect 12176 16708 12204 16748
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 16117 16779 16175 16785
rect 16117 16776 16129 16779
rect 12676 16748 13492 16776
rect 12676 16736 12682 16748
rect 10928 16680 12204 16708
rect 10928 16668 10934 16680
rect 12342 16668 12348 16720
rect 12400 16668 12406 16720
rect 10689 16643 10747 16649
rect 10468 16612 10548 16640
rect 10468 16600 10474 16612
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 4065 16575 4123 16581
rect 1811 16544 4016 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 3988 16504 4016 16544
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 5074 16572 5080 16584
rect 4111 16544 5080 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 5074 16532 5080 16544
rect 5132 16532 5138 16584
rect 5166 16532 5172 16584
rect 5224 16532 5230 16584
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 5276 16544 9413 16572
rect 5276 16504 5304 16544
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9401 16535 9459 16541
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 10520 16581 10548 16612
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 11882 16640 11888 16652
rect 10735 16612 11888 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 10505 16575 10563 16581
rect 9824 16544 10180 16572
rect 9824 16532 9830 16544
rect 3988 16476 5304 16504
rect 5905 16507 5963 16513
rect 2501 16467 2559 16473
rect 5905 16473 5917 16507
rect 5951 16504 5963 16507
rect 7282 16504 7288 16516
rect 5951 16476 7288 16504
rect 5951 16473 5963 16476
rect 5905 16467 5963 16473
rect 7282 16464 7288 16476
rect 7340 16464 7346 16516
rect 9030 16504 9036 16516
rect 8128 16476 9036 16504
rect 2590 16396 2596 16448
rect 2648 16436 2654 16448
rect 6454 16436 6460 16448
rect 2648 16408 6460 16436
rect 2648 16396 2654 16408
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 6822 16436 6828 16448
rect 6687 16408 6828 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6972 16408 7021 16436
rect 6972 16396 6978 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7009 16399 7067 16405
rect 7837 16439 7895 16445
rect 7837 16405 7849 16439
rect 7883 16436 7895 16439
rect 8128 16436 8156 16476
rect 9030 16464 9036 16476
rect 9088 16464 9094 16516
rect 9217 16507 9275 16513
rect 9217 16473 9229 16507
rect 9263 16473 9275 16507
rect 9217 16467 9275 16473
rect 7883 16408 8156 16436
rect 7883 16405 7895 16408
rect 7837 16399 7895 16405
rect 8202 16396 8208 16448
rect 8260 16396 8266 16448
rect 9232 16436 9260 16467
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 9858 16504 9864 16516
rect 9364 16476 9864 16504
rect 9364 16464 9370 16476
rect 9858 16464 9864 16476
rect 9916 16464 9922 16516
rect 10152 16504 10180 16544
rect 10505 16541 10517 16575
rect 10551 16541 10563 16575
rect 10505 16535 10563 16541
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 12360 16572 12388 16668
rect 13464 16649 13492 16748
rect 13556 16748 16129 16776
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 11655 16544 12388 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 13556 16572 13584 16748
rect 16117 16745 16129 16748
rect 16163 16776 16175 16779
rect 16206 16776 16212 16788
rect 16163 16748 16212 16776
rect 16163 16745 16175 16748
rect 16117 16739 16175 16745
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16356 16748 16405 16776
rect 16356 16736 16362 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 19702 16776 19708 16788
rect 16816 16748 19708 16776
rect 16816 16736 16822 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 30926 16776 30932 16788
rect 21232 16748 30932 16776
rect 21232 16736 21238 16748
rect 30926 16736 30932 16748
rect 30984 16736 30990 16788
rect 18322 16708 18328 16720
rect 13648 16680 18328 16708
rect 13648 16649 13676 16680
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 22278 16668 22284 16720
rect 22336 16708 22342 16720
rect 25685 16711 25743 16717
rect 25685 16708 25697 16711
rect 22336 16680 22600 16708
rect 22336 16668 22342 16680
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 14516 16612 15485 16640
rect 14516 16600 14522 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 16298 16640 16304 16652
rect 15703 16612 16304 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16640 16819 16643
rect 17218 16640 17224 16652
rect 16807 16612 17224 16640
rect 16807 16609 16819 16612
rect 16761 16603 16819 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20438 16640 20444 16652
rect 19751 16612 20444 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 22572 16649 22600 16680
rect 25148 16680 25697 16708
rect 25148 16652 25176 16680
rect 25685 16677 25697 16680
rect 25731 16708 25743 16711
rect 25866 16708 25872 16720
rect 25731 16680 25872 16708
rect 25731 16677 25743 16680
rect 25685 16671 25743 16677
rect 25866 16668 25872 16680
rect 25924 16668 25930 16720
rect 25958 16668 25964 16720
rect 26016 16668 26022 16720
rect 28276 16680 28948 16708
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 20772 16612 22477 16640
rect 20772 16600 20778 16612
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16609 22615 16643
rect 22557 16603 22615 16609
rect 22830 16600 22836 16652
rect 22888 16640 22894 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 22888 16612 23765 16640
rect 22888 16600 22894 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 25130 16600 25136 16652
rect 25188 16600 25194 16652
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16640 25375 16643
rect 25774 16640 25780 16652
rect 25363 16612 25780 16640
rect 25363 16609 25375 16612
rect 25317 16603 25375 16609
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 27062 16600 27068 16652
rect 27120 16600 27126 16652
rect 27154 16600 27160 16652
rect 27212 16600 27218 16652
rect 28276 16649 28304 16680
rect 28261 16643 28319 16649
rect 28261 16609 28273 16643
rect 28307 16609 28319 16643
rect 28261 16603 28319 16609
rect 28445 16643 28503 16649
rect 28445 16609 28457 16643
rect 28491 16640 28503 16643
rect 28810 16640 28816 16652
rect 28491 16612 28816 16640
rect 28491 16609 28503 16612
rect 28445 16603 28503 16609
rect 28810 16600 28816 16612
rect 28868 16600 28874 16652
rect 28920 16649 28948 16680
rect 28905 16643 28963 16649
rect 28905 16609 28917 16643
rect 28951 16640 28963 16643
rect 31938 16640 31944 16652
rect 28951 16612 31944 16640
rect 28951 16609 28963 16612
rect 28905 16603 28963 16609
rect 31938 16600 31944 16612
rect 31996 16600 32002 16652
rect 12584 16544 13584 16572
rect 14553 16575 14611 16581
rect 12584 16532 12590 16544
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 15286 16572 15292 16584
rect 14599 16544 15292 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 15378 16532 15384 16584
rect 15436 16532 15442 16584
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16572 18291 16575
rect 18322 16572 18328 16584
rect 18279 16544 18328 16572
rect 18279 16541 18291 16544
rect 18233 16535 18291 16541
rect 10152 16476 11836 16504
rect 9582 16436 9588 16448
rect 9232 16408 9588 16436
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 9766 16396 9772 16448
rect 9824 16396 9830 16448
rect 10413 16439 10471 16445
rect 10413 16405 10425 16439
rect 10459 16436 10471 16439
rect 10502 16436 10508 16448
rect 10459 16408 10508 16436
rect 10459 16405 10471 16408
rect 10413 16399 10471 16405
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 11238 16396 11244 16448
rect 11296 16396 11302 16448
rect 11698 16396 11704 16448
rect 11756 16396 11762 16448
rect 11808 16436 11836 16476
rect 11882 16464 11888 16516
rect 11940 16504 11946 16516
rect 12342 16504 12348 16516
rect 11940 16476 12348 16504
rect 11940 16464 11946 16476
rect 12342 16464 12348 16476
rect 12400 16464 12406 16516
rect 12802 16464 12808 16516
rect 12860 16504 12866 16516
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 12860 16476 13369 16504
rect 12860 16464 12866 16476
rect 13357 16473 13369 16476
rect 13403 16473 13415 16507
rect 16666 16504 16672 16516
rect 13357 16467 13415 16473
rect 14292 16476 16672 16504
rect 12158 16436 12164 16448
rect 11808 16408 12164 16436
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 12989 16439 13047 16445
rect 12989 16405 13001 16439
rect 13035 16436 13047 16439
rect 14292 16436 14320 16476
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 17218 16504 17224 16516
rect 17000 16476 17224 16504
rect 17000 16464 17006 16476
rect 17218 16464 17224 16476
rect 17276 16504 17282 16516
rect 17604 16504 17632 16535
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16572 22431 16575
rect 23290 16572 23296 16584
rect 22419 16544 23296 16572
rect 22419 16541 22431 16544
rect 22373 16535 22431 16541
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 24302 16572 24308 16584
rect 23615 16544 24308 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 24302 16532 24308 16544
rect 24360 16532 24366 16584
rect 25038 16532 25044 16584
rect 25096 16572 25102 16584
rect 25096 16544 26740 16572
rect 25096 16532 25102 16544
rect 19334 16504 19340 16516
rect 17276 16476 17540 16504
rect 17604 16476 19340 16504
rect 17276 16464 17282 16476
rect 13035 16408 14320 16436
rect 13035 16405 13047 16408
rect 12989 16399 13047 16405
rect 14366 16396 14372 16448
rect 14424 16396 14430 16448
rect 14826 16396 14832 16448
rect 14884 16436 14890 16448
rect 15013 16439 15071 16445
rect 15013 16436 15025 16439
rect 14884 16408 15025 16436
rect 14884 16396 14890 16408
rect 15013 16405 15025 16408
rect 15059 16405 15071 16439
rect 15013 16399 15071 16405
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 16114 16436 16120 16448
rect 15252 16408 16120 16436
rect 15252 16396 15258 16408
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 16206 16396 16212 16448
rect 16264 16396 16270 16448
rect 16758 16396 16764 16448
rect 16816 16436 16822 16448
rect 17405 16439 17463 16445
rect 17405 16436 17417 16439
rect 16816 16408 17417 16436
rect 16816 16396 16822 16408
rect 17405 16405 17417 16408
rect 17451 16405 17463 16439
rect 17512 16436 17540 16476
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 20162 16464 20168 16516
rect 20220 16464 20226 16516
rect 21450 16464 21456 16516
rect 21508 16464 21514 16516
rect 23661 16507 23719 16513
rect 23661 16473 23673 16507
rect 23707 16504 23719 16507
rect 23842 16504 23848 16516
rect 23707 16476 23848 16504
rect 23707 16473 23719 16476
rect 23661 16467 23719 16473
rect 23842 16464 23848 16476
rect 23900 16464 23906 16516
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 24176 16476 26648 16504
rect 24176 16464 24182 16476
rect 17678 16436 17684 16448
rect 17512 16408 17684 16436
rect 17405 16399 17463 16405
rect 17678 16396 17684 16408
rect 17736 16396 17742 16448
rect 18049 16439 18107 16445
rect 18049 16405 18061 16439
rect 18095 16436 18107 16439
rect 18506 16436 18512 16448
rect 18095 16408 18512 16436
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 18598 16396 18604 16448
rect 18656 16436 18662 16448
rect 18693 16439 18751 16445
rect 18693 16436 18705 16439
rect 18656 16408 18705 16436
rect 18656 16396 18662 16408
rect 18693 16405 18705 16408
rect 18739 16405 18751 16439
rect 18693 16399 18751 16405
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 20772 16408 22017 16436
rect 20772 16396 20778 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 22462 16396 22468 16448
rect 22520 16436 22526 16448
rect 23201 16439 23259 16445
rect 23201 16436 23213 16439
rect 22520 16408 23213 16436
rect 22520 16396 22526 16408
rect 23201 16405 23213 16408
rect 23247 16405 23259 16439
rect 23201 16399 23259 16405
rect 23750 16396 23756 16448
rect 23808 16436 23814 16448
rect 24673 16439 24731 16445
rect 24673 16436 24685 16439
rect 23808 16408 24685 16436
rect 23808 16396 23814 16408
rect 24673 16405 24685 16408
rect 24719 16405 24731 16439
rect 24673 16399 24731 16405
rect 25038 16396 25044 16448
rect 25096 16436 25102 16448
rect 25958 16436 25964 16448
rect 25096 16408 25964 16436
rect 25096 16396 25102 16408
rect 25958 16396 25964 16408
rect 26016 16396 26022 16448
rect 26620 16445 26648 16476
rect 26605 16439 26663 16445
rect 26605 16405 26617 16439
rect 26651 16405 26663 16439
rect 26712 16436 26740 16544
rect 27706 16532 27712 16584
rect 27764 16572 27770 16584
rect 28169 16575 28227 16581
rect 28169 16572 28181 16575
rect 27764 16544 28181 16572
rect 27764 16532 27770 16544
rect 28169 16541 28181 16544
rect 28215 16541 28227 16575
rect 28169 16535 28227 16541
rect 26973 16507 27031 16513
rect 26973 16473 26985 16507
rect 27019 16504 27031 16507
rect 28442 16504 28448 16516
rect 27019 16476 28448 16504
rect 27019 16473 27031 16476
rect 26973 16467 27031 16473
rect 28442 16464 28448 16476
rect 28500 16464 28506 16516
rect 27801 16439 27859 16445
rect 27801 16436 27813 16439
rect 26712 16408 27813 16436
rect 26605 16399 26663 16405
rect 27801 16405 27813 16408
rect 27847 16405 27859 16439
rect 27801 16399 27859 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 7190 16192 7196 16244
rect 7248 16232 7254 16244
rect 7285 16235 7343 16241
rect 7285 16232 7297 16235
rect 7248 16204 7297 16232
rect 7248 16192 7254 16204
rect 7285 16201 7297 16204
rect 7331 16201 7343 16235
rect 8846 16232 8852 16244
rect 7285 16195 7343 16201
rect 7484 16204 8852 16232
rect 4338 16124 4344 16176
rect 4396 16124 4402 16176
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 1811 16068 2774 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2746 16028 2774 16068
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 5626 16056 5632 16108
rect 5684 16056 5690 16108
rect 5721 16099 5779 16105
rect 5721 16065 5733 16099
rect 5767 16096 5779 16099
rect 5994 16096 6000 16108
rect 5767 16068 6000 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 5994 16056 6000 16068
rect 6052 16096 6058 16108
rect 7484 16096 7512 16204
rect 8846 16192 8852 16204
rect 8904 16192 8910 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9732 16204 10640 16232
rect 9732 16192 9738 16204
rect 8386 16164 8392 16176
rect 6052 16068 7512 16096
rect 7576 16136 8392 16164
rect 6052 16056 6058 16068
rect 4706 16028 4712 16040
rect 2746 16000 4712 16028
rect 2041 15991 2099 15997
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 5902 15988 5908 16040
rect 5960 16028 5966 16040
rect 6546 16028 6552 16040
rect 5960 16000 6552 16028
rect 5960 15988 5966 16000
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 6638 15988 6644 16040
rect 6696 15988 6702 16040
rect 7576 16028 7604 16136
rect 8386 16124 8392 16136
rect 8444 16164 8450 16176
rect 10612 16173 10640 16204
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11606 16232 11612 16244
rect 11204 16204 11612 16232
rect 11204 16192 11210 16204
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 12250 16192 12256 16244
rect 12308 16232 12314 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 12308 16204 13737 16232
rect 12308 16192 12314 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 14734 16192 14740 16244
rect 14792 16232 14798 16244
rect 14792 16204 17080 16232
rect 14792 16192 14798 16204
rect 8757 16167 8815 16173
rect 8757 16164 8769 16167
rect 8444 16136 8769 16164
rect 8444 16124 8450 16136
rect 8757 16133 8769 16136
rect 8803 16133 8815 16167
rect 8757 16127 8815 16133
rect 10597 16167 10655 16173
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 10778 16164 10784 16176
rect 10643 16136 10784 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 10778 16124 10784 16136
rect 10836 16164 10842 16176
rect 12526 16164 12532 16176
rect 10836 16136 12532 16164
rect 10836 16124 10842 16136
rect 12526 16124 12532 16136
rect 12584 16124 12590 16176
rect 14645 16167 14703 16173
rect 14645 16133 14657 16167
rect 14691 16164 14703 16167
rect 16482 16164 16488 16176
rect 14691 16136 16488 16164
rect 14691 16133 14703 16136
rect 14645 16127 14703 16133
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 16942 16164 16948 16176
rect 16592 16136 16948 16164
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16096 7803 16099
rect 7926 16096 7932 16108
rect 7791 16068 7932 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 7926 16056 7932 16068
rect 7984 16056 7990 16108
rect 8478 16056 8484 16108
rect 8536 16056 8542 16108
rect 9858 16056 9864 16108
rect 9916 16056 9922 16108
rect 10134 16096 10140 16108
rect 9968 16068 10140 16096
rect 7392 16000 7604 16028
rect 7837 16031 7895 16037
rect 6178 15920 6184 15972
rect 6236 15960 6242 15972
rect 7392 15960 7420 16000
rect 7837 15997 7849 16031
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 6236 15932 7420 15960
rect 6236 15920 6242 15932
rect 7466 15920 7472 15972
rect 7524 15960 7530 15972
rect 7852 15960 7880 15991
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 9968 16028 9996 16068
rect 10134 16056 10140 16068
rect 10192 16096 10198 16108
rect 10686 16096 10692 16108
rect 10192 16068 10692 16096
rect 10192 16056 10198 16068
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 10928 16068 11161 16096
rect 10928 16056 10934 16068
rect 11149 16065 11161 16068
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 11974 16056 11980 16108
rect 12032 16056 12038 16108
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 14918 16096 14924 16108
rect 14783 16068 14924 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 14918 16056 14924 16068
rect 14976 16096 14982 16108
rect 16301 16099 16359 16105
rect 14976 16068 15608 16096
rect 14976 16056 14982 16068
rect 8444 16000 9996 16028
rect 8444 15988 8450 16000
rect 10226 15988 10232 16040
rect 10284 15988 10290 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 16028 12311 16031
rect 13538 16028 13544 16040
rect 12299 16000 13544 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 14829 15991 14887 15997
rect 14936 16000 15485 16028
rect 7524 15932 7880 15960
rect 7524 15920 7530 15932
rect 10962 15920 10968 15972
rect 11020 15920 11026 15972
rect 14844 15960 14872 15991
rect 13280 15932 14872 15960
rect 5258 15852 5264 15904
rect 5316 15852 5322 15904
rect 5810 15852 5816 15904
rect 5868 15892 5874 15904
rect 7926 15892 7932 15904
rect 5868 15864 7932 15892
rect 5868 15852 5874 15864
rect 7926 15852 7932 15864
rect 7984 15892 7990 15904
rect 11422 15892 11428 15904
rect 7984 15864 11428 15892
rect 7984 15852 7990 15864
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 13280 15892 13308 15932
rect 12676 15864 13308 15892
rect 12676 15852 12682 15864
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13688 15864 14289 15892
rect 13688 15852 13694 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 14734 15852 14740 15904
rect 14792 15892 14798 15904
rect 14936 15892 14964 16000
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 15580 16028 15608 16068
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16390 16096 16396 16108
rect 16347 16068 16396 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16592 16028 16620 16136
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 17052 16164 17080 16204
rect 17126 16192 17132 16244
rect 17184 16192 17190 16244
rect 18598 16232 18604 16244
rect 17788 16204 18604 16232
rect 17788 16164 17816 16204
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 20441 16235 20499 16241
rect 20441 16232 20453 16235
rect 18748 16204 20453 16232
rect 18748 16192 18754 16204
rect 20441 16201 20453 16204
rect 20487 16201 20499 16235
rect 20806 16232 20812 16244
rect 20441 16195 20499 16201
rect 20548 16204 20812 16232
rect 17052 16136 17816 16164
rect 17865 16167 17923 16173
rect 17865 16133 17877 16167
rect 17911 16164 17923 16167
rect 20548 16164 20576 16204
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 21266 16192 21272 16244
rect 21324 16192 21330 16244
rect 21468 16204 24900 16232
rect 17911 16136 20576 16164
rect 17911 16133 17923 16136
rect 17865 16127 17923 16133
rect 16666 16056 16672 16108
rect 16724 16096 16730 16108
rect 17773 16099 17831 16105
rect 17773 16096 17785 16099
rect 16724 16068 17785 16096
rect 16724 16056 16730 16068
rect 17773 16065 17785 16068
rect 17819 16065 17831 16099
rect 18601 16099 18659 16105
rect 17773 16059 17831 16065
rect 17880 16068 18092 16096
rect 15580 16000 16620 16028
rect 16761 16031 16819 16037
rect 15473 15991 15531 15997
rect 16761 15997 16773 16031
rect 16807 16028 16819 16031
rect 17218 16028 17224 16040
rect 16807 16000 17224 16028
rect 16807 15997 16819 16000
rect 16761 15991 16819 15997
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 17880 16028 17908 16068
rect 17368 16000 17908 16028
rect 17957 16031 18015 16037
rect 17368 15988 17374 16000
rect 17957 15997 17969 16031
rect 18003 15997 18015 16031
rect 18064 16028 18092 16068
rect 18601 16065 18613 16099
rect 18647 16096 18659 16099
rect 19150 16096 19156 16108
rect 18647 16068 19156 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 19702 16056 19708 16108
rect 19760 16096 19766 16108
rect 21468 16105 21496 16204
rect 24872 16164 24900 16204
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 26605 16235 26663 16241
rect 26605 16232 26617 16235
rect 25004 16204 26617 16232
rect 25004 16192 25010 16204
rect 26605 16201 26617 16204
rect 26651 16201 26663 16235
rect 26605 16195 26663 16201
rect 25222 16164 25228 16176
rect 24872 16136 25228 16164
rect 25222 16124 25228 16136
rect 25280 16124 25286 16176
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 19760 16068 20545 16096
rect 19760 16056 19766 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16065 21511 16099
rect 21453 16059 21511 16065
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16096 22339 16099
rect 22554 16096 22560 16108
rect 22327 16068 22560 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16096 23719 16099
rect 24302 16096 24308 16108
rect 23707 16068 24308 16096
rect 23707 16065 23719 16068
rect 23661 16059 23719 16065
rect 24302 16056 24308 16068
rect 24360 16056 24366 16108
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 24670 16096 24676 16108
rect 24627 16068 24676 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 24670 16056 24676 16068
rect 24728 16056 24734 16108
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 26234 16056 26240 16108
rect 26292 16096 26298 16108
rect 26694 16096 26700 16108
rect 26292 16068 26700 16096
rect 26292 16056 26298 16068
rect 26694 16056 26700 16068
rect 26752 16096 26758 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26752 16068 26985 16096
rect 26752 16056 26758 16068
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18064 16000 18889 16028
rect 17957 15991 18015 15997
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 16028 20775 16031
rect 21266 16028 21272 16040
rect 20763 16000 21272 16028
rect 20763 15997 20775 16000
rect 20717 15991 20775 15997
rect 17405 15963 17463 15969
rect 17405 15960 17417 15963
rect 16500 15932 17417 15960
rect 14792 15864 14964 15892
rect 14792 15852 14798 15864
rect 15194 15852 15200 15904
rect 15252 15892 15258 15904
rect 16117 15895 16175 15901
rect 16117 15892 16129 15895
rect 15252 15864 16129 15892
rect 15252 15852 15258 15864
rect 16117 15861 16129 15864
rect 16163 15861 16175 15895
rect 16117 15855 16175 15861
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 16500 15892 16528 15932
rect 17405 15929 17417 15932
rect 17451 15929 17463 15963
rect 17405 15923 17463 15929
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 17972 15960 18000 15991
rect 21266 15988 21272 16000
rect 21324 15988 21330 16040
rect 21358 15988 21364 16040
rect 21416 16028 21422 16040
rect 21910 16028 21916 16040
rect 21416 16000 21916 16028
rect 21416 15988 21422 16000
rect 21910 15988 21916 16000
rect 21968 16028 21974 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 21968 16000 22017 16028
rect 21968 15988 21974 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 23474 16028 23480 16040
rect 22005 15991 22063 15997
rect 22112 16000 23480 16028
rect 17552 15932 18000 15960
rect 17552 15920 17558 15932
rect 16264 15864 16528 15892
rect 20073 15895 20131 15901
rect 16264 15852 16270 15864
rect 20073 15861 20085 15895
rect 20119 15892 20131 15895
rect 22112 15892 22140 16000
rect 23474 15988 23480 16000
rect 23532 15988 23538 16040
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 23842 16028 23848 16040
rect 23799 16000 23848 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 23937 16031 23995 16037
rect 23937 15997 23949 16031
rect 23983 16028 23995 16031
rect 24026 16028 24032 16040
rect 23983 16000 24032 16028
rect 23983 15997 23995 16000
rect 23937 15991 23995 15997
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24762 15988 24768 16040
rect 24820 16028 24826 16040
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24820 16000 25145 16028
rect 24820 15988 24826 16000
rect 25133 15997 25145 16000
rect 25179 16028 25191 16031
rect 27154 16028 27160 16040
rect 25179 16000 27160 16028
rect 25179 15997 25191 16000
rect 25133 15991 25191 15997
rect 27154 15988 27160 16000
rect 27212 15988 27218 16040
rect 26142 15920 26148 15972
rect 26200 15960 26206 15972
rect 29730 15960 29736 15972
rect 26200 15932 29736 15960
rect 26200 15920 26206 15932
rect 29730 15920 29736 15932
rect 29788 15920 29794 15972
rect 20119 15864 22140 15892
rect 20119 15861 20131 15864
rect 20073 15855 20131 15861
rect 22646 15852 22652 15904
rect 22704 15892 22710 15904
rect 23293 15895 23351 15901
rect 23293 15892 23305 15895
rect 22704 15864 23305 15892
rect 22704 15852 22710 15864
rect 23293 15861 23305 15864
rect 23339 15861 23351 15895
rect 23293 15855 23351 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 2924 15660 3433 15688
rect 2924 15648 2930 15660
rect 3421 15657 3433 15660
rect 3467 15688 3479 15691
rect 3467 15660 8340 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 3605 15623 3663 15629
rect 3605 15589 3617 15623
rect 3651 15620 3663 15623
rect 3970 15620 3976 15632
rect 3651 15592 3976 15620
rect 3651 15589 3663 15592
rect 3605 15583 3663 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 5350 15620 5356 15632
rect 4356 15592 5356 15620
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 3694 15512 3700 15564
rect 3752 15552 3758 15564
rect 4356 15552 4384 15592
rect 5350 15580 5356 15592
rect 5408 15580 5414 15632
rect 7834 15580 7840 15632
rect 7892 15580 7898 15632
rect 3752 15524 4384 15552
rect 3752 15512 3758 15524
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 3418 15484 3424 15496
rect 1811 15456 3424 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 4632 15484 4660 15515
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5592 15524 5641 15552
rect 5592 15512 5598 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 5810 15512 5816 15564
rect 5868 15512 5874 15564
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6788 15524 6837 15552
rect 6788 15512 6794 15524
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 6914 15512 6920 15564
rect 6972 15512 6978 15564
rect 8312 15561 8340 15660
rect 8754 15648 8760 15700
rect 8812 15688 8818 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8812 15660 9321 15688
rect 8812 15648 8818 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 12802 15688 12808 15700
rect 9309 15651 9367 15657
rect 10244 15660 12808 15688
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 8386 15512 8392 15564
rect 8444 15512 8450 15564
rect 10244 15561 10272 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 12912 15660 14320 15688
rect 10318 15580 10324 15632
rect 10376 15620 10382 15632
rect 10873 15623 10931 15629
rect 10873 15620 10885 15623
rect 10376 15592 10885 15620
rect 10376 15580 10382 15592
rect 10873 15589 10885 15592
rect 10919 15589 10931 15623
rect 10873 15583 10931 15589
rect 12066 15580 12072 15632
rect 12124 15580 12130 15632
rect 12158 15580 12164 15632
rect 12216 15620 12222 15632
rect 12912 15620 12940 15660
rect 12216 15592 12940 15620
rect 14292 15620 14320 15660
rect 15838 15648 15844 15700
rect 15896 15648 15902 15700
rect 19429 15691 19487 15697
rect 19429 15688 19441 15691
rect 15948 15660 19441 15688
rect 15948 15620 15976 15660
rect 19429 15657 19441 15660
rect 19475 15657 19487 15691
rect 19429 15651 19487 15657
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 19889 15691 19947 15697
rect 19889 15688 19901 15691
rect 19668 15660 19901 15688
rect 19668 15648 19674 15660
rect 19889 15657 19901 15660
rect 19935 15657 19947 15691
rect 19889 15651 19947 15657
rect 21910 15648 21916 15700
rect 21968 15688 21974 15700
rect 22557 15691 22615 15697
rect 22557 15688 22569 15691
rect 21968 15660 22569 15688
rect 21968 15648 21974 15660
rect 22557 15657 22569 15660
rect 22603 15657 22615 15691
rect 22557 15651 22615 15657
rect 23842 15648 23848 15700
rect 23900 15688 23906 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 23900 15660 24501 15688
rect 23900 15648 23906 15660
rect 24489 15657 24501 15660
rect 24535 15688 24547 15691
rect 24670 15688 24676 15700
rect 24535 15660 24676 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 24670 15648 24676 15660
rect 24728 15648 24734 15700
rect 26326 15620 26332 15632
rect 14292 15592 15976 15620
rect 25700 15592 26332 15620
rect 12216 15580 12222 15592
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15521 10287 15555
rect 10229 15515 10287 15521
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 10744 15524 11437 15552
rect 10744 15512 10750 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11425 15515 11483 15521
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12894 15552 12900 15564
rect 12759 15524 12900 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 14090 15552 14096 15564
rect 13412 15524 14096 15552
rect 13412 15512 13418 15524
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 15010 15512 15016 15564
rect 15068 15512 15074 15564
rect 16114 15512 16120 15564
rect 16172 15552 16178 15564
rect 16485 15555 16543 15561
rect 16172 15524 16344 15552
rect 16172 15512 16178 15524
rect 5902 15484 5908 15496
rect 4632 15456 5908 15484
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 12437 15487 12495 15493
rect 12437 15484 12449 15487
rect 6696 15456 12449 15484
rect 6696 15444 6702 15456
rect 12437 15453 12449 15456
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13722 15484 13728 15496
rect 13311 15456 13728 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 14829 15487 14887 15493
rect 14829 15484 14841 15487
rect 14792 15456 14841 15484
rect 14792 15444 14798 15456
rect 14829 15453 14841 15456
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 16206 15444 16212 15496
rect 16264 15444 16270 15496
rect 5537 15419 5595 15425
rect 5537 15416 5549 15419
rect 3988 15388 5549 15416
rect 3988 15357 4016 15388
rect 5537 15385 5549 15388
rect 5583 15385 5595 15419
rect 5537 15379 5595 15385
rect 6733 15419 6791 15425
rect 6733 15385 6745 15419
rect 6779 15416 6791 15419
rect 6779 15388 8340 15416
rect 6779 15385 6791 15388
rect 6733 15379 6791 15385
rect 3973 15351 4031 15357
rect 3973 15317 3985 15351
rect 4019 15317 4031 15351
rect 3973 15311 4031 15317
rect 4338 15308 4344 15360
rect 4396 15308 4402 15360
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5350 15348 5356 15360
rect 5215 15320 5356 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 5994 15348 6000 15360
rect 5868 15320 6000 15348
rect 5868 15308 5874 15320
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 6362 15308 6368 15360
rect 6420 15308 6426 15360
rect 6454 15308 6460 15360
rect 6512 15348 6518 15360
rect 7466 15348 7472 15360
rect 6512 15320 7472 15348
rect 6512 15308 6518 15320
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 7616 15320 8217 15348
rect 7616 15308 7622 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8312 15348 8340 15388
rect 8478 15376 8484 15428
rect 8536 15416 8542 15428
rect 9217 15419 9275 15425
rect 9217 15416 9229 15419
rect 8536 15388 9229 15416
rect 8536 15376 8542 15388
rect 9217 15385 9229 15388
rect 9263 15385 9275 15419
rect 9217 15379 9275 15385
rect 11146 15376 11152 15428
rect 11204 15416 11210 15428
rect 11241 15419 11299 15425
rect 11241 15416 11253 15419
rect 11204 15388 11253 15416
rect 11204 15376 11210 15388
rect 11241 15385 11253 15388
rect 11287 15385 11299 15419
rect 11241 15379 11299 15385
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 14921 15419 14979 15425
rect 14921 15416 14933 15419
rect 12308 15388 13584 15416
rect 12308 15376 12314 15388
rect 9490 15348 9496 15360
rect 8312 15320 9496 15348
rect 8205 15311 8263 15317
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 9769 15351 9827 15357
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 9858 15348 9864 15360
rect 9815 15320 9864 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 11333 15351 11391 15357
rect 11333 15348 11345 15351
rect 10008 15320 11345 15348
rect 10008 15308 10014 15320
rect 11333 15317 11345 15320
rect 11379 15348 11391 15351
rect 11606 15348 11612 15360
rect 11379 15320 11612 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 13556 15357 13584 15388
rect 13740 15388 14933 15416
rect 13740 15360 13768 15388
rect 14921 15385 14933 15388
rect 14967 15385 14979 15419
rect 16224 15416 16252 15444
rect 14921 15379 14979 15385
rect 15396 15388 16252 15416
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15317 13599 15351
rect 13541 15311 13599 15317
rect 13722 15308 13728 15360
rect 13780 15308 13786 15360
rect 14182 15308 14188 15360
rect 14240 15348 14246 15360
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 14240 15320 14473 15348
rect 14240 15308 14246 15320
rect 14461 15317 14473 15320
rect 14507 15317 14519 15351
rect 14461 15311 14519 15317
rect 14642 15308 14648 15360
rect 14700 15348 14706 15360
rect 15396 15348 15424 15388
rect 14700 15320 15424 15348
rect 14700 15308 14706 15320
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 16316 15357 16344 15524
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 16500 15416 16528 15515
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19484 15524 20269 15552
rect 19484 15512 19490 15524
rect 20257 15521 20269 15524
rect 20303 15552 20315 15555
rect 20622 15552 20628 15564
rect 20303 15524 20628 15552
rect 20303 15521 20315 15524
rect 20257 15515 20315 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 20990 15512 20996 15564
rect 21048 15552 21054 15564
rect 25700 15561 25728 15592
rect 26326 15580 26332 15592
rect 26384 15620 26390 15632
rect 26421 15623 26479 15629
rect 26421 15620 26433 15623
rect 26384 15592 26433 15620
rect 26384 15580 26390 15592
rect 26421 15589 26433 15592
rect 26467 15589 26479 15623
rect 26421 15583 26479 15589
rect 25685 15555 25743 15561
rect 25685 15552 25697 15555
rect 21048 15524 22048 15552
rect 21048 15512 21054 15524
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 20162 15484 20168 15496
rect 19659 15456 20168 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 22020 15480 22048 15524
rect 22204 15524 25697 15552
rect 22204 15480 22232 15524
rect 25685 15521 25697 15524
rect 25731 15521 25743 15555
rect 25685 15515 25743 15521
rect 25774 15512 25780 15564
rect 25832 15512 25838 15564
rect 22020 15452 22232 15480
rect 22833 15487 22891 15493
rect 22833 15453 22845 15487
rect 22879 15484 22891 15487
rect 22922 15484 22928 15496
rect 22879 15456 22928 15484
rect 22879 15453 22891 15456
rect 22833 15447 22891 15453
rect 22922 15444 22928 15456
rect 22980 15484 22986 15496
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 22980 15456 23121 15484
rect 22980 15444 22986 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 25590 15444 25596 15496
rect 25648 15484 25654 15496
rect 26329 15487 26387 15493
rect 26329 15484 26341 15487
rect 25648 15456 26341 15484
rect 25648 15444 25654 15456
rect 26329 15453 26341 15456
rect 26375 15484 26387 15487
rect 26970 15484 26976 15496
rect 26375 15456 26976 15484
rect 26375 15453 26387 15456
rect 26329 15447 26387 15453
rect 26970 15444 26976 15456
rect 27028 15484 27034 15496
rect 27028 15456 35894 15484
rect 27028 15444 27034 15456
rect 17310 15416 17316 15428
rect 16500 15388 17316 15416
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17770 15376 17776 15428
rect 17828 15376 17834 15428
rect 19978 15376 19984 15428
rect 20036 15416 20042 15428
rect 20533 15419 20591 15425
rect 20533 15416 20545 15419
rect 20036 15388 20545 15416
rect 20036 15376 20042 15388
rect 20533 15385 20545 15388
rect 20579 15385 20591 15419
rect 21758 15388 22232 15416
rect 20533 15379 20591 15385
rect 16209 15351 16267 15357
rect 16209 15348 16221 15351
rect 15528 15320 16221 15348
rect 15528 15308 15534 15320
rect 16209 15317 16221 15320
rect 16255 15317 16267 15351
rect 16209 15311 16267 15317
rect 16301 15351 16359 15357
rect 16301 15317 16313 15351
rect 16347 15348 16359 15351
rect 16390 15348 16396 15360
rect 16347 15320 16396 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 17460 15320 18797 15348
rect 17460 15308 17466 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 19150 15308 19156 15360
rect 19208 15348 19214 15360
rect 21450 15348 21456 15360
rect 19208 15320 21456 15348
rect 19208 15308 19214 15320
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21968 15320 22017 15348
rect 21968 15308 21974 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22204 15348 22232 15388
rect 23934 15376 23940 15428
rect 23992 15376 23998 15428
rect 35866 15416 35894 15456
rect 43438 15416 43444 15428
rect 35866 15388 43444 15416
rect 43438 15376 43444 15388
rect 43496 15376 43502 15428
rect 22373 15351 22431 15357
rect 22373 15348 22385 15351
rect 22204 15320 22385 15348
rect 22005 15311 22063 15317
rect 22373 15317 22385 15320
rect 22419 15348 22431 15351
rect 23382 15348 23388 15360
rect 22419 15320 23388 15348
rect 22419 15317 22431 15320
rect 22373 15311 22431 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 25222 15308 25228 15360
rect 25280 15308 25286 15360
rect 26326 15308 26332 15360
rect 26384 15348 26390 15360
rect 46198 15348 46204 15360
rect 26384 15320 46204 15348
rect 26384 15308 26390 15320
rect 46198 15308 46204 15320
rect 46256 15308 46262 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 566 15104 572 15156
rect 624 15144 630 15156
rect 1118 15144 1124 15156
rect 624 15116 1124 15144
rect 624 15104 630 15116
rect 1118 15104 1124 15116
rect 1176 15104 1182 15156
rect 3510 15104 3516 15156
rect 3568 15104 3574 15156
rect 4706 15104 4712 15156
rect 4764 15144 4770 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 4764 15116 6745 15144
rect 4764 15104 4770 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 6733 15107 6791 15113
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 8478 15144 8484 15156
rect 7524 15116 8484 15144
rect 7524 15104 7530 15116
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 8665 15147 8723 15153
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 9214 15144 9220 15156
rect 8711 15116 9220 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 9585 15147 9643 15153
rect 9585 15113 9597 15147
rect 9631 15144 9643 15147
rect 11238 15144 11244 15156
rect 9631 15116 11244 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12768 15116 13001 15144
rect 12768 15104 12774 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 15470 15144 15476 15156
rect 13320 15116 15476 15144
rect 13320 15104 13326 15116
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 22094 15144 22100 15156
rect 18472 15116 22100 15144
rect 18472 15104 18478 15116
rect 22094 15104 22100 15116
rect 22152 15144 22158 15156
rect 22922 15144 22928 15156
rect 22152 15116 22928 15144
rect 22152 15104 22158 15116
rect 22922 15104 22928 15116
rect 22980 15144 22986 15156
rect 23290 15144 23296 15156
rect 22980 15116 23296 15144
rect 22980 15104 22986 15116
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 5994 15076 6000 15088
rect 5658 15048 6000 15076
rect 5994 15036 6000 15048
rect 6052 15076 6058 15088
rect 6270 15076 6276 15088
rect 6052 15048 6276 15076
rect 6052 15036 6058 15048
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 6641 15079 6699 15085
rect 6641 15045 6653 15079
rect 6687 15076 6699 15079
rect 8386 15076 8392 15088
rect 6687 15048 8392 15076
rect 6687 15045 6699 15048
rect 6641 15039 6699 15045
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 1811 14980 2774 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 1118 14900 1124 14952
rect 1176 14940 1182 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1176 14912 2053 14940
rect 1176 14900 1182 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2746 14940 2774 14980
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3568 14980 3709 15008
rect 3568 14968 3574 14980
rect 3697 14977 3709 14980
rect 3743 15008 3755 15011
rect 3878 15008 3884 15020
rect 3743 14980 3884 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4154 14968 4160 15020
rect 4212 14968 4218 15020
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 6656 15008 6684 15039
rect 8386 15036 8392 15048
rect 8444 15036 8450 15088
rect 9030 15036 9036 15088
rect 9088 15076 9094 15088
rect 9677 15079 9735 15085
rect 9677 15076 9689 15079
rect 9088 15048 9689 15076
rect 9088 15036 9094 15048
rect 9677 15045 9689 15048
rect 9723 15045 9735 15079
rect 9677 15039 9735 15045
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 10226 15076 10232 15088
rect 9824 15048 10232 15076
rect 9824 15036 9830 15048
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 10778 15036 10784 15088
rect 10836 15036 10842 15088
rect 10962 15036 10968 15088
rect 11020 15076 11026 15088
rect 14185 15079 14243 15085
rect 14185 15076 14197 15079
rect 11020 15048 14197 15076
rect 11020 15036 11026 15048
rect 14185 15045 14197 15048
rect 14231 15076 14243 15079
rect 14734 15076 14740 15088
rect 14231 15048 14740 15076
rect 14231 15045 14243 15048
rect 14185 15039 14243 15045
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 14829 15079 14887 15085
rect 14829 15045 14841 15079
rect 14875 15076 14887 15079
rect 14918 15076 14924 15088
rect 14875 15048 14924 15076
rect 14875 15045 14887 15048
rect 14829 15039 14887 15045
rect 14918 15036 14924 15048
rect 14976 15036 14982 15088
rect 17770 15076 17776 15088
rect 16054 15048 17776 15076
rect 17770 15036 17776 15048
rect 17828 15076 17834 15088
rect 18138 15076 18144 15088
rect 17828 15048 18144 15076
rect 17828 15036 17834 15048
rect 18138 15036 18144 15048
rect 18196 15076 18202 15088
rect 19153 15079 19211 15085
rect 19153 15076 19165 15079
rect 18196 15048 19165 15076
rect 18196 15036 18202 15048
rect 19153 15045 19165 15048
rect 19199 15045 19211 15079
rect 19153 15039 19211 15045
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 20714 15076 20720 15088
rect 20211 15048 20720 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 22281 15079 22339 15085
rect 22281 15045 22293 15079
rect 22327 15076 22339 15079
rect 22554 15076 22560 15088
rect 22327 15048 22560 15076
rect 22327 15045 22339 15048
rect 22281 15039 22339 15045
rect 22554 15036 22560 15048
rect 22612 15036 22618 15088
rect 24964 15076 24992 15104
rect 25133 15079 25191 15085
rect 25133 15076 25145 15079
rect 24964 15048 25145 15076
rect 25133 15045 25145 15048
rect 25179 15045 25191 15079
rect 25133 15039 25191 15045
rect 6236 14980 6684 15008
rect 6236 14968 6242 14980
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 7653 15011 7711 15017
rect 7653 15008 7665 15011
rect 7340 14980 7665 15008
rect 7340 14968 7346 14980
rect 7653 14977 7665 14980
rect 7699 15008 7711 15011
rect 7699 14980 8064 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 2746 14912 5488 14940
rect 2041 14903 2099 14909
rect 5460 14872 5488 14912
rect 6270 14900 6276 14952
rect 6328 14940 6334 14952
rect 7745 14943 7803 14949
rect 7745 14940 7757 14943
rect 6328 14912 7757 14940
rect 6328 14900 6334 14912
rect 7745 14909 7757 14912
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 7190 14872 7196 14884
rect 5460 14844 7196 14872
rect 7190 14832 7196 14844
rect 7248 14832 7254 14884
rect 7760 14872 7788 14903
rect 7926 14900 7932 14952
rect 7984 14900 7990 14952
rect 8036 14940 8064 14980
rect 8570 14968 8576 15020
rect 8628 14968 8634 15020
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 8904 14980 10885 15008
rect 8904 14968 8910 14980
rect 10873 14977 10885 14980
rect 10919 15008 10931 15011
rect 10919 14980 11928 15008
rect 10919 14977 10931 14980
rect 10873 14971 10931 14977
rect 9861 14943 9919 14949
rect 8036 14912 9352 14940
rect 8386 14872 8392 14884
rect 7760 14844 8392 14872
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 8478 14832 8484 14884
rect 8536 14872 8542 14884
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 8536 14844 9229 14872
rect 8536 14832 8542 14844
rect 9217 14841 9229 14844
rect 9263 14841 9275 14875
rect 9217 14835 9275 14841
rect 4420 14807 4478 14813
rect 4420 14773 4432 14807
rect 4466 14804 4478 14807
rect 4890 14804 4896 14816
rect 4466 14776 4896 14804
rect 4466 14773 4478 14776
rect 4420 14767 4478 14773
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 5905 14807 5963 14813
rect 5905 14804 5917 14807
rect 5132 14776 5917 14804
rect 5132 14764 5138 14776
rect 5905 14773 5917 14776
rect 5951 14804 5963 14807
rect 6914 14804 6920 14816
rect 5951 14776 6920 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 9324 14804 9352 14912
rect 9861 14909 9873 14943
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14909 11759 14943
rect 11900 14940 11928 14980
rect 11974 14968 11980 15020
rect 12032 14968 12038 15020
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 12894 15008 12900 15020
rect 12676 14980 12900 15008
rect 12676 14968 12682 14980
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13495 14980 14013 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 14001 14977 14013 14980
rect 14047 15008 14059 15011
rect 14366 15008 14372 15020
rect 14047 14980 14372 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 19518 14968 19524 15020
rect 19576 15008 19582 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19576 14980 20085 15008
rect 19576 14968 19582 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20180 14980 20484 15008
rect 13262 14940 13268 14952
rect 11900 14912 13268 14940
rect 11701 14903 11759 14909
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 9876 14872 9904 14903
rect 10778 14872 10784 14884
rect 9732 14844 10784 14872
rect 9732 14832 9738 14844
rect 10778 14832 10784 14844
rect 10836 14832 10842 14884
rect 10980 14872 11008 14903
rect 10888 14844 11008 14872
rect 11716 14872 11744 14903
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13538 14900 13544 14952
rect 13596 14900 13602 14952
rect 13648 14912 14228 14940
rect 11716 14844 12940 14872
rect 10226 14804 10232 14816
rect 9324 14776 10232 14804
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 10410 14764 10416 14816
rect 10468 14764 10474 14816
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 10888 14804 10916 14844
rect 10560 14776 10916 14804
rect 10560 14764 10566 14776
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 12710 14804 12716 14816
rect 11112 14776 12716 14804
rect 11112 14764 11118 14776
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 12912 14804 12940 14844
rect 13648 14804 13676 14912
rect 14200 14872 14228 14912
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 14332 14912 14565 14940
rect 14332 14900 14338 14912
rect 14553 14909 14565 14912
rect 14599 14909 14611 14943
rect 16850 14940 16856 14952
rect 14553 14903 14611 14909
rect 14660 14912 16856 14940
rect 14660 14872 14688 14912
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 18966 14900 18972 14952
rect 19024 14940 19030 14952
rect 20180 14940 20208 14980
rect 19024 14912 20208 14940
rect 20349 14943 20407 14949
rect 19024 14900 19030 14912
rect 20349 14909 20361 14943
rect 20395 14909 20407 14943
rect 20456 14940 20484 14980
rect 20622 14968 20628 15020
rect 20680 15008 20686 15020
rect 22002 15008 22008 15020
rect 20680 14980 22008 15008
rect 20680 14968 20686 14980
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 23382 14968 23388 15020
rect 23440 15008 23446 15020
rect 23440 14980 23612 15008
rect 23440 14968 23446 14980
rect 23584 14952 23612 14980
rect 23934 14968 23940 15020
rect 23992 15008 23998 15020
rect 24857 15011 24915 15017
rect 24857 15008 24869 15011
rect 23992 14980 24869 15008
rect 23992 14968 23998 14980
rect 24857 14977 24869 14980
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 26234 14968 26240 15020
rect 26292 14968 26298 15020
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20456 14912 20913 14940
rect 20349 14903 20407 14909
rect 20901 14909 20913 14912
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 16758 14872 16764 14884
rect 14200 14844 14688 14872
rect 15856 14844 16764 14872
rect 12912 14776 13676 14804
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 15856 14804 15884 14844
rect 16758 14832 16764 14844
rect 16816 14832 16822 14884
rect 19705 14875 19763 14881
rect 17512 14844 19472 14872
rect 13872 14776 15884 14804
rect 13872 14764 13878 14776
rect 16298 14764 16304 14816
rect 16356 14764 16362 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16669 14807 16727 14813
rect 16669 14804 16681 14807
rect 16448 14776 16681 14804
rect 16448 14764 16454 14776
rect 16669 14773 16681 14776
rect 16715 14804 16727 14807
rect 17512 14804 17540 14844
rect 16715 14776 17540 14804
rect 16715 14773 16727 14776
rect 16669 14767 16727 14773
rect 17586 14764 17592 14816
rect 17644 14804 17650 14816
rect 18966 14804 18972 14816
rect 17644 14776 18972 14804
rect 17644 14764 17650 14776
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 19334 14764 19340 14816
rect 19392 14764 19398 14816
rect 19444 14804 19472 14844
rect 19705 14841 19717 14875
rect 19751 14872 19763 14875
rect 19794 14872 19800 14884
rect 19751 14844 19800 14872
rect 19751 14841 19763 14844
rect 19705 14835 19763 14841
rect 19794 14832 19800 14844
rect 19852 14832 19858 14884
rect 20364 14872 20392 14903
rect 23566 14900 23572 14952
rect 23624 14940 23630 14952
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 23624 14912 24041 14940
rect 23624 14900 23630 14912
rect 24029 14909 24041 14912
rect 24075 14940 24087 14943
rect 24213 14943 24271 14949
rect 24213 14940 24225 14943
rect 24075 14912 24225 14940
rect 24075 14909 24087 14912
rect 24029 14903 24087 14909
rect 24213 14909 24225 14912
rect 24259 14940 24271 14943
rect 26252 14940 26280 14968
rect 26973 14943 27031 14949
rect 26973 14940 26985 14943
rect 24259 14912 26985 14940
rect 24259 14909 24271 14912
rect 24213 14903 24271 14909
rect 26973 14909 26985 14912
rect 27019 14909 27031 14943
rect 26973 14903 27031 14909
rect 21910 14872 21916 14884
rect 20364 14844 21916 14872
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 23658 14832 23664 14884
rect 23716 14872 23722 14884
rect 23753 14875 23811 14881
rect 23753 14872 23765 14875
rect 23716 14844 23765 14872
rect 23716 14832 23722 14844
rect 23753 14841 23765 14844
rect 23799 14841 23811 14875
rect 24854 14872 24860 14884
rect 23753 14835 23811 14841
rect 23952 14844 24860 14872
rect 23952 14804 23980 14844
rect 24854 14832 24860 14844
rect 24912 14832 24918 14884
rect 19444 14776 23980 14804
rect 26602 14764 26608 14816
rect 26660 14764 26666 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 6454 14600 6460 14612
rect 3936 14572 6460 14600
rect 3936 14560 3942 14572
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 10962 14600 10968 14612
rect 6788 14572 10968 14600
rect 6788 14560 6794 14572
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 13354 14600 13360 14612
rect 11624 14572 13360 14600
rect 3973 14535 4031 14541
rect 3973 14501 3985 14535
rect 4019 14532 4031 14535
rect 4019 14504 5580 14532
rect 4019 14501 4031 14504
rect 3973 14495 4031 14501
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14464 4951 14467
rect 5074 14464 5080 14476
rect 4939 14436 5080 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5552 14464 5580 14504
rect 6822 14492 6828 14544
rect 6880 14532 6886 14544
rect 6880 14504 8248 14532
rect 6880 14492 6886 14504
rect 6178 14464 6184 14476
rect 5552 14436 6184 14464
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 7193 14467 7251 14473
rect 7193 14433 7205 14467
rect 7239 14464 7251 14467
rect 7558 14464 7564 14476
rect 7239 14436 7564 14464
rect 7239 14433 7251 14436
rect 7193 14427 7251 14433
rect 7558 14424 7564 14436
rect 7616 14464 7622 14476
rect 7834 14464 7840 14476
rect 7616 14436 7840 14464
rect 7616 14424 7622 14436
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 1762 14356 1768 14408
rect 1820 14356 1826 14408
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14396 4675 14399
rect 5166 14396 5172 14408
rect 4663 14368 5172 14396
rect 4663 14365 4675 14368
rect 4617 14359 4675 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5442 14356 5448 14408
rect 5500 14356 5506 14408
rect 8220 14405 8248 14504
rect 8386 14492 8392 14544
rect 8444 14532 8450 14544
rect 11624 14541 11652 14572
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13725 14603 13783 14609
rect 13725 14600 13737 14603
rect 13596 14572 13737 14600
rect 13596 14560 13602 14572
rect 13725 14569 13737 14572
rect 13771 14569 13783 14603
rect 13725 14563 13783 14569
rect 14090 14560 14096 14612
rect 14148 14560 14154 14612
rect 14366 14560 14372 14612
rect 14424 14560 14430 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 14976 14572 18613 14600
rect 14976 14560 14982 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 18601 14563 18659 14569
rect 18690 14560 18696 14612
rect 18748 14600 18754 14612
rect 22370 14600 22376 14612
rect 18748 14572 22376 14600
rect 18748 14560 18754 14572
rect 22370 14560 22376 14572
rect 22428 14560 22434 14612
rect 26970 14560 26976 14612
rect 27028 14560 27034 14612
rect 11609 14535 11667 14541
rect 11609 14532 11621 14535
rect 8444 14504 11621 14532
rect 8444 14492 8450 14504
rect 11609 14501 11621 14504
rect 11655 14501 11667 14535
rect 11609 14495 11667 14501
rect 18138 14492 18144 14544
rect 18196 14532 18202 14544
rect 18877 14535 18935 14541
rect 18877 14532 18889 14535
rect 18196 14504 18889 14532
rect 18196 14492 18202 14504
rect 18877 14501 18889 14504
rect 18923 14501 18935 14535
rect 18877 14495 18935 14501
rect 21726 14492 21732 14544
rect 21784 14492 21790 14544
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 24029 14535 24087 14541
rect 24029 14532 24041 14535
rect 23716 14504 24041 14532
rect 23716 14492 23722 14504
rect 24029 14501 24041 14504
rect 24075 14532 24087 14535
rect 25774 14532 25780 14544
rect 24075 14504 25780 14532
rect 24075 14501 24087 14504
rect 24029 14495 24087 14501
rect 25774 14492 25780 14504
rect 25832 14492 25838 14544
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 9674 14464 9680 14476
rect 8527 14436 9680 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 9953 14467 10011 14473
rect 9953 14464 9965 14467
rect 9824 14436 9965 14464
rect 9824 14424 9830 14436
rect 9953 14433 9965 14436
rect 9999 14433 10011 14467
rect 9953 14427 10011 14433
rect 10042 14424 10048 14476
rect 10100 14464 10106 14476
rect 10502 14464 10508 14476
rect 10100 14436 10508 14464
rect 10100 14424 10106 14436
rect 10502 14424 10508 14436
rect 10560 14464 10566 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10560 14436 11161 14464
rect 10560 14424 10566 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 12253 14467 12311 14473
rect 12253 14433 12265 14467
rect 12299 14464 12311 14467
rect 12618 14464 12624 14476
rect 12299 14436 12624 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 14550 14464 14556 14476
rect 12768 14436 14556 14464
rect 12768 14424 12774 14436
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 16298 14464 16304 14476
rect 14967 14436 16304 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14464 16911 14467
rect 17126 14464 17132 14476
rect 16899 14436 17132 14464
rect 16899 14433 16911 14436
rect 16853 14427 16911 14433
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17218 14424 17224 14476
rect 17276 14464 17282 14476
rect 18322 14464 18328 14476
rect 17276 14436 18328 14464
rect 17276 14424 17282 14436
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 19852 14436 21097 14464
rect 19852 14424 19858 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 9306 14396 9312 14408
rect 8343 14368 9312 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10318 14396 10324 14408
rect 9907 14368 10324 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11054 14396 11060 14408
rect 11011 14368 11060 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11974 14356 11980 14408
rect 12032 14356 12038 14408
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 14090 14396 14096 14408
rect 13412 14368 14096 14396
rect 13412 14356 13418 14368
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 14332 14368 14657 14396
rect 14332 14356 14338 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 14645 14359 14703 14365
rect 18432 14368 19625 14396
rect 5350 14328 5356 14340
rect 4264 14300 5356 14328
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14260 3479 14263
rect 3605 14263 3663 14269
rect 3605 14260 3617 14263
rect 3467 14232 3617 14260
rect 3467 14229 3479 14232
rect 3421 14223 3479 14229
rect 3605 14229 3617 14232
rect 3651 14260 3663 14263
rect 3970 14260 3976 14272
rect 3651 14232 3976 14260
rect 3651 14229 3663 14232
rect 3605 14223 3663 14229
rect 3970 14220 3976 14232
rect 4028 14220 4034 14272
rect 4264 14269 4292 14300
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 5721 14331 5779 14337
rect 5721 14297 5733 14331
rect 5767 14297 5779 14331
rect 5721 14291 5779 14297
rect 4249 14263 4307 14269
rect 4249 14229 4261 14263
rect 4295 14229 4307 14263
rect 4249 14223 4307 14229
rect 4706 14220 4712 14272
rect 4764 14220 4770 14272
rect 5736 14260 5764 14291
rect 5994 14288 6000 14340
rect 6052 14328 6058 14340
rect 15194 14328 15200 14340
rect 6052 14300 6210 14328
rect 7210 14300 12434 14328
rect 6052 14288 6058 14300
rect 5902 14260 5908 14272
rect 5736 14232 5908 14260
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 6454 14220 6460 14272
rect 6512 14260 6518 14272
rect 7210 14260 7238 14300
rect 6512 14232 7238 14260
rect 6512 14220 6518 14232
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8904 14232 9045 14260
rect 8904 14220 8910 14232
rect 9033 14229 9045 14232
rect 9079 14229 9091 14263
rect 9033 14223 9091 14229
rect 9398 14220 9404 14272
rect 9456 14220 9462 14272
rect 9766 14220 9772 14272
rect 9824 14220 9830 14272
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 11020 14232 11069 14260
rect 11020 14220 11026 14232
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 12406 14260 12434 14300
rect 14016 14300 15200 14328
rect 14016 14260 14044 14300
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15470 14288 15476 14340
rect 15528 14288 15534 14340
rect 17129 14331 17187 14337
rect 16316 14300 17080 14328
rect 12406 14232 14044 14260
rect 11057 14223 11115 14229
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 16316 14260 16344 14300
rect 14884 14232 16344 14260
rect 14884 14220 14890 14232
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 17052 14260 17080 14300
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17402 14328 17408 14340
rect 17175 14300 17408 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 18138 14288 18144 14340
rect 18196 14288 18202 14340
rect 18432 14260 18460 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 20898 14356 20904 14408
rect 20956 14356 20962 14408
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14396 21051 14399
rect 21744 14396 21772 14492
rect 22002 14424 22008 14476
rect 22060 14464 22066 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22060 14436 22293 14464
rect 22060 14424 22066 14436
rect 22281 14433 22293 14436
rect 22327 14464 22339 14467
rect 23934 14464 23940 14476
rect 22327 14436 23940 14464
rect 22327 14433 22339 14436
rect 22281 14427 22339 14433
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14464 25191 14467
rect 26329 14467 26387 14473
rect 26329 14464 26341 14467
rect 25179 14436 26341 14464
rect 25179 14433 25191 14436
rect 25133 14427 25191 14433
rect 26329 14433 26341 14436
rect 26375 14464 26387 14467
rect 26602 14464 26608 14476
rect 26375 14436 26608 14464
rect 26375 14433 26387 14436
rect 26329 14427 26387 14433
rect 25148 14396 25176 14427
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 21039 14368 21772 14396
rect 23952 14368 25176 14396
rect 26145 14399 26203 14405
rect 21039 14365 21051 14368
rect 20993 14359 21051 14365
rect 20916 14328 20944 14356
rect 21545 14331 21603 14337
rect 21545 14328 21557 14331
rect 20916 14300 21557 14328
rect 21545 14297 21557 14300
rect 21591 14328 21603 14331
rect 21818 14328 21824 14340
rect 21591 14300 21824 14328
rect 21591 14297 21603 14300
rect 21545 14291 21603 14297
rect 21818 14288 21824 14300
rect 21876 14288 21882 14340
rect 21910 14288 21916 14340
rect 21968 14328 21974 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 21968 14300 22569 14328
rect 21968 14288 21974 14300
rect 22557 14297 22569 14300
rect 22603 14297 22615 14331
rect 22557 14291 22615 14297
rect 23566 14288 23572 14340
rect 23624 14288 23630 14340
rect 17052 14232 18460 14260
rect 19426 14220 19432 14272
rect 19484 14220 19490 14272
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 21634 14260 21640 14272
rect 20956 14232 21640 14260
rect 20956 14220 20962 14232
rect 21634 14220 21640 14232
rect 21692 14220 21698 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23952 14260 23980 14368
rect 26145 14365 26157 14399
rect 26191 14396 26203 14399
rect 26970 14396 26976 14408
rect 26191 14368 26976 14396
rect 26191 14365 26203 14368
rect 26145 14359 26203 14365
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 24946 14288 24952 14340
rect 25004 14288 25010 14340
rect 25041 14331 25099 14337
rect 25041 14297 25053 14331
rect 25087 14328 25099 14331
rect 25130 14328 25136 14340
rect 25087 14300 25136 14328
rect 25087 14297 25099 14300
rect 25041 14291 25099 14297
rect 25130 14288 25136 14300
rect 25188 14288 25194 14340
rect 26237 14331 26295 14337
rect 26237 14297 26249 14331
rect 26283 14328 26295 14331
rect 26326 14328 26332 14340
rect 26283 14300 26332 14328
rect 26283 14297 26295 14300
rect 26237 14291 26295 14297
rect 26326 14288 26332 14300
rect 26384 14328 26390 14340
rect 26789 14331 26847 14337
rect 26789 14328 26801 14331
rect 26384 14300 26801 14328
rect 26384 14288 26390 14300
rect 26789 14297 26801 14300
rect 26835 14297 26847 14331
rect 26789 14291 26847 14297
rect 22796 14232 23980 14260
rect 22796 14220 22802 14232
rect 24578 14220 24584 14272
rect 24636 14220 24642 14272
rect 24964 14260 24992 14288
rect 25682 14260 25688 14272
rect 24964 14232 25688 14260
rect 25682 14220 25688 14232
rect 25740 14220 25746 14272
rect 25774 14220 25780 14272
rect 25832 14220 25838 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 4706 14056 4712 14068
rect 4111 14028 4712 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 6362 14056 6368 14068
rect 5675 14028 6368 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 4525 13991 4583 13997
rect 4525 13988 4537 13991
rect 2372 13960 4537 13988
rect 2372 13948 2378 13960
rect 4525 13957 4537 13960
rect 4571 13957 4583 13991
rect 4525 13951 4583 13957
rect 5350 13948 5356 14000
rect 5408 13988 5414 14000
rect 5721 13991 5779 13997
rect 5721 13988 5733 13991
rect 5408 13960 5733 13988
rect 5408 13948 5414 13960
rect 5721 13957 5733 13960
rect 5767 13957 5779 13991
rect 6932 13988 6960 14019
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 9214 14056 9220 14068
rect 8159 14028 9220 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11112 14028 11989 14056
rect 11112 14016 11118 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 14369 14059 14427 14065
rect 13219 14028 14320 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 6932 13960 8493 13988
rect 5721 13951 5779 13957
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 9490 13948 9496 14000
rect 9548 13988 9554 14000
rect 9858 13988 9864 14000
rect 9548 13960 9864 13988
rect 9548 13948 9554 13960
rect 9858 13948 9864 13960
rect 9916 13988 9922 14000
rect 9916 13960 10074 13988
rect 9916 13948 9922 13960
rect 11606 13948 11612 14000
rect 11664 13988 11670 14000
rect 13633 13991 13691 13997
rect 13633 13988 13645 13991
rect 11664 13960 13645 13988
rect 11664 13948 11670 13960
rect 13633 13957 13645 13960
rect 13679 13957 13691 13991
rect 14292 13988 14320 14028
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 14458 14056 14464 14068
rect 14415 14028 14464 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 14734 14016 14740 14068
rect 14792 14016 14798 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 17218 14056 17224 14068
rect 15611 14028 17224 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 17368 14028 18889 14056
rect 17368 14016 17374 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 18966 14016 18972 14068
rect 19024 14056 19030 14068
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 19024 14028 20085 14056
rect 19024 14016 19030 14028
rect 20073 14025 20085 14028
rect 20119 14025 20131 14059
rect 20073 14019 20131 14025
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 21232 14028 23397 14056
rect 21232 14016 21238 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 24949 14059 25007 14065
rect 24949 14025 24961 14059
rect 24995 14056 25007 14059
rect 25774 14056 25780 14068
rect 24995 14028 25780 14056
rect 24995 14025 25007 14028
rect 24949 14019 25007 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 16666 13988 16672 14000
rect 14292 13960 16672 13988
rect 13633 13951 13691 13957
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 16761 13991 16819 13997
rect 16761 13957 16773 13991
rect 16807 13988 16819 13991
rect 17678 13988 17684 14000
rect 16807 13960 17684 13988
rect 16807 13957 16819 13960
rect 16761 13951 16819 13957
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1762 13920 1768 13932
rect 1544 13892 1768 13920
rect 1544 13880 1550 13892
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 3620 13784 3648 13883
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 3936 13892 4445 13920
rect 3936 13880 3942 13892
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 5316 13892 7389 13920
rect 5316 13880 5322 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 11940 13892 12357 13920
rect 11940 13880 11946 13892
rect 12345 13889 12357 13892
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 13170 13920 13176 13932
rect 12676 13892 13176 13920
rect 12676 13880 12682 13892
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 13538 13880 13544 13932
rect 13596 13880 13602 13932
rect 13740 13892 13952 13920
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4798 13852 4804 13864
rect 4755 13824 4804 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 5828 13784 5856 13815
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6730 13852 6736 13864
rect 6420 13824 6736 13852
rect 6420 13812 6426 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 7926 13852 7932 13864
rect 7616 13824 7932 13852
rect 7616 13812 7622 13824
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 5902 13784 5908 13796
rect 3620 13756 5396 13784
rect 5828 13756 5908 13784
rect 2130 13676 2136 13728
rect 2188 13716 2194 13728
rect 4614 13716 4620 13728
rect 2188 13688 4620 13716
rect 2188 13676 2194 13688
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 5258 13676 5264 13728
rect 5316 13676 5322 13728
rect 5368 13716 5396 13756
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 6546 13744 6552 13796
rect 6604 13744 6610 13796
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 8680 13784 8708 13815
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 9631 13824 10732 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 8628 13756 8708 13784
rect 10704 13784 10732 13824
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 10836 13824 11069 13852
rect 10836 13812 10842 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12216 13824 12449 13852
rect 12216 13812 12222 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 12894 13852 12900 13864
rect 12575 13824 12900 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 12544 13784 12572 13815
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13630 13852 13636 13864
rect 13004 13824 13636 13852
rect 10704 13756 12572 13784
rect 8628 13744 8634 13756
rect 12710 13744 12716 13796
rect 12768 13784 12774 13796
rect 13004 13784 13032 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 13740 13784 13768 13892
rect 13817 13855 13875 13861
rect 13817 13821 13829 13855
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 12768 13756 13032 13784
rect 13096 13756 13768 13784
rect 12768 13744 12774 13756
rect 6454 13716 6460 13728
rect 5368 13688 6460 13716
rect 6454 13676 6460 13688
rect 6512 13676 6518 13728
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 13096 13716 13124 13756
rect 7248 13688 13124 13716
rect 7248 13676 7254 13688
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13630 13716 13636 13728
rect 13228 13688 13636 13716
rect 13228 13676 13234 13688
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 13832 13716 13860 13815
rect 13924 13784 13952 13892
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 14148 13892 15332 13920
rect 14148 13880 14154 13892
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 14829 13855 14887 13861
rect 14829 13852 14841 13855
rect 14608 13824 14841 13852
rect 14608 13812 14614 13824
rect 14829 13821 14841 13824
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 14918 13812 14924 13864
rect 14976 13812 14982 13864
rect 15304 13796 15332 13892
rect 15562 13880 15568 13932
rect 15620 13920 15626 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15620 13892 15945 13920
rect 15620 13880 15626 13892
rect 15933 13889 15945 13892
rect 15979 13889 15991 13923
rect 16776 13920 16804 13951
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 18138 13948 18144 14000
rect 18196 13948 18202 14000
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 19484 13960 24532 13988
rect 19484 13948 19490 13960
rect 15933 13883 15991 13889
rect 16132 13892 16804 13920
rect 19613 13923 19671 13929
rect 16022 13812 16028 13864
rect 16080 13812 16086 13864
rect 16132 13796 16160 13892
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 14366 13784 14372 13796
rect 13924 13756 14372 13784
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 15470 13784 15476 13796
rect 15344 13756 15476 13784
rect 15344 13744 15350 13756
rect 15470 13744 15476 13756
rect 15528 13744 15534 13796
rect 16114 13744 16120 13796
rect 16172 13744 16178 13796
rect 16224 13784 16252 13815
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 17405 13855 17463 13861
rect 17405 13821 17417 13855
rect 17451 13852 17463 13855
rect 17494 13852 17500 13864
rect 17451 13824 17500 13852
rect 17451 13821 17463 13824
rect 17405 13815 17463 13821
rect 17494 13812 17500 13824
rect 17552 13812 17558 13864
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 19628 13852 19656 13883
rect 20438 13880 20444 13932
rect 20496 13880 20502 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 21634 13920 21640 13932
rect 20579 13892 21640 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 21818 13880 21824 13932
rect 21876 13880 21882 13932
rect 22370 13880 22376 13932
rect 22428 13920 22434 13932
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22428 13892 22569 13920
rect 22428 13880 22434 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 22695 13892 23244 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 20346 13852 20352 13864
rect 17920 13824 19656 13852
rect 19720 13824 20352 13852
rect 17920 13812 17926 13824
rect 19429 13787 19487 13793
rect 16224 13756 17264 13784
rect 17034 13716 17040 13728
rect 13832 13688 17040 13716
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 17236 13716 17264 13756
rect 19429 13753 19441 13787
rect 19475 13784 19487 13787
rect 19720 13784 19748 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 22664 13852 22692 13883
rect 20625 13815 20683 13821
rect 20824 13824 22232 13852
rect 19475 13756 19748 13784
rect 20640 13784 20668 13815
rect 20714 13784 20720 13796
rect 20640 13756 20720 13784
rect 19475 13753 19487 13756
rect 19429 13747 19487 13753
rect 20714 13744 20720 13756
rect 20772 13744 20778 13796
rect 19150 13716 19156 13728
rect 17236 13688 19156 13716
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20824 13716 20852 13824
rect 22204 13793 22232 13824
rect 22296 13824 22692 13852
rect 22189 13787 22247 13793
rect 22189 13753 22201 13787
rect 22235 13753 22247 13787
rect 22189 13747 22247 13753
rect 20220 13688 20852 13716
rect 20220 13676 20226 13688
rect 21818 13676 21824 13728
rect 21876 13716 21882 13728
rect 22296 13716 22324 13824
rect 22830 13812 22836 13864
rect 22888 13812 22894 13864
rect 23216 13852 23244 13892
rect 23382 13880 23388 13932
rect 23440 13920 23446 13932
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 23440 13892 23765 13920
rect 23440 13880 23446 13892
rect 23753 13889 23765 13892
rect 23799 13920 23811 13923
rect 24504 13920 24532 13960
rect 24578 13948 24584 14000
rect 24636 13988 24642 14000
rect 25041 13991 25099 13997
rect 25041 13988 25053 13991
rect 24636 13960 25053 13988
rect 24636 13948 24642 13960
rect 25041 13957 25053 13960
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 25130 13948 25136 14000
rect 25188 13988 25194 14000
rect 25593 13991 25651 13997
rect 25593 13988 25605 13991
rect 25188 13960 25605 13988
rect 25188 13948 25194 13960
rect 25593 13957 25605 13960
rect 25639 13957 25651 13991
rect 25593 13951 25651 13957
rect 25682 13948 25688 14000
rect 25740 13988 25746 14000
rect 25869 13991 25927 13997
rect 25869 13988 25881 13991
rect 25740 13960 25881 13988
rect 25740 13948 25746 13960
rect 25869 13957 25881 13960
rect 25915 13957 25927 13991
rect 25869 13951 25927 13957
rect 34974 13920 34980 13932
rect 23799 13892 24164 13920
rect 24504 13892 34980 13920
rect 23799 13889 23811 13892
rect 23753 13883 23811 13889
rect 23842 13852 23848 13864
rect 23216 13824 23848 13852
rect 23842 13812 23848 13824
rect 23900 13812 23906 13864
rect 24026 13812 24032 13864
rect 24084 13812 24090 13864
rect 24136 13852 24164 13892
rect 34974 13880 34980 13892
rect 35032 13880 35038 13932
rect 24136 13824 25084 13852
rect 25056 13784 25084 13824
rect 25130 13812 25136 13864
rect 25188 13852 25194 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 25188 13824 25237 13852
rect 25188 13812 25194 13824
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 26145 13855 26203 13861
rect 26145 13852 26157 13855
rect 25271 13824 26157 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 26145 13821 26157 13824
rect 26191 13821 26203 13855
rect 26145 13815 26203 13821
rect 25961 13787 26019 13793
rect 25961 13784 25973 13787
rect 25056 13756 25973 13784
rect 25961 13753 25973 13756
rect 26007 13753 26019 13787
rect 25961 13747 26019 13753
rect 21876 13688 22324 13716
rect 21876 13676 21882 13688
rect 24578 13676 24584 13728
rect 24636 13676 24642 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 3786 13512 3792 13524
rect 3384 13484 3792 13512
rect 3384 13472 3390 13484
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 4798 13512 4804 13524
rect 4080 13484 4804 13512
rect 2038 13336 2044 13388
rect 2096 13336 2102 13388
rect 1762 13268 1768 13320
rect 1820 13268 1826 13320
rect 3510 13200 3516 13252
rect 3568 13200 3574 13252
rect 4080 13240 4108 13484
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5166 13472 5172 13524
rect 5224 13512 5230 13524
rect 5626 13512 5632 13524
rect 5224 13484 5632 13512
rect 5224 13472 5230 13484
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 6052 13484 6469 13512
rect 6052 13472 6058 13484
rect 6457 13481 6469 13484
rect 6503 13512 6515 13515
rect 9766 13512 9772 13524
rect 6503 13484 9772 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 12710 13512 12716 13524
rect 11624 13484 12716 13512
rect 8386 13404 8392 13456
rect 8444 13444 8450 13456
rect 8481 13447 8539 13453
rect 8481 13444 8493 13447
rect 8444 13416 8493 13444
rect 8444 13404 8450 13416
rect 8481 13413 8493 13416
rect 8527 13444 8539 13447
rect 8570 13444 8576 13456
rect 8527 13416 8576 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 8570 13404 8576 13416
rect 8628 13444 8634 13456
rect 8628 13416 11008 13444
rect 8628 13404 8634 13416
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 5442 13376 5448 13388
rect 4212 13348 5448 13376
rect 4212 13336 4218 13348
rect 5442 13336 5448 13348
rect 5500 13376 5506 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 5500 13348 6745 13376
rect 5500 13336 5506 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 5810 13308 5816 13320
rect 5566 13280 5816 13308
rect 5810 13268 5816 13280
rect 5868 13308 5874 13320
rect 6270 13308 6276 13320
rect 5868 13280 6276 13308
rect 5868 13268 5874 13280
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 3804 13212 4108 13240
rect 4433 13243 4491 13249
rect 2406 13132 2412 13184
rect 2464 13172 2470 13184
rect 3421 13175 3479 13181
rect 3421 13172 3433 13175
rect 2464 13144 3433 13172
rect 2464 13132 2470 13144
rect 3421 13141 3433 13144
rect 3467 13172 3479 13175
rect 3804 13172 3832 13212
rect 4433 13209 4445 13243
rect 4479 13209 4491 13243
rect 6748 13240 6776 13339
rect 7558 13336 7564 13388
rect 7616 13376 7622 13388
rect 8294 13376 8300 13388
rect 7616 13348 8300 13376
rect 7616 13336 7622 13348
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 10980 13385 11008 13416
rect 11146 13404 11152 13456
rect 11204 13444 11210 13456
rect 11425 13447 11483 13453
rect 11425 13444 11437 13447
rect 11204 13416 11437 13444
rect 11204 13404 11210 13416
rect 11425 13413 11437 13416
rect 11471 13413 11483 13447
rect 11425 13407 11483 13413
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13308 10839 13311
rect 11624 13308 11652 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13688 13484 13737 13512
rect 13688 13472 13694 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15068 13484 16037 13512
rect 15068 13472 15074 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 17552 13484 18889 13512
rect 17552 13472 17558 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 18966 13472 18972 13524
rect 19024 13512 19030 13524
rect 19150 13512 19156 13524
rect 19024 13484 19156 13512
rect 19024 13472 19030 13484
rect 19150 13472 19156 13484
rect 19208 13512 19214 13524
rect 20606 13515 20664 13521
rect 20606 13512 20618 13515
rect 19208 13484 20618 13512
rect 19208 13472 19214 13484
rect 20606 13481 20618 13484
rect 20652 13481 20664 13515
rect 20606 13475 20664 13481
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22554 13512 22560 13524
rect 22143 13484 22560 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23937 13515 23995 13521
rect 23937 13512 23949 13515
rect 23348 13484 23949 13512
rect 23348 13472 23354 13484
rect 23937 13481 23949 13484
rect 23983 13481 23995 13515
rect 23937 13475 23995 13481
rect 11701 13447 11759 13453
rect 11701 13413 11713 13447
rect 11747 13444 11759 13447
rect 11882 13444 11888 13456
rect 11747 13416 11888 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 21634 13404 21640 13456
rect 21692 13444 21698 13456
rect 22833 13447 22891 13453
rect 22833 13444 22845 13447
rect 21692 13416 22845 13444
rect 21692 13404 21698 13416
rect 22833 13413 22845 13416
rect 22879 13413 22891 13447
rect 23750 13444 23756 13456
rect 22833 13407 22891 13413
rect 23308 13416 23756 13444
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 13262 13376 13268 13388
rect 12032 13348 13268 13376
rect 12032 13336 12038 13348
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15194 13376 15200 13388
rect 14599 13348 15200 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15194 13336 15200 13348
rect 15252 13376 15258 13388
rect 16390 13376 16396 13388
rect 15252 13348 16396 13376
rect 15252 13336 15258 13348
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17494 13376 17500 13388
rect 17184 13348 17500 13376
rect 17184 13336 17190 13348
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 22186 13376 22192 13388
rect 20395 13348 22192 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 23308 13385 23336 13416
rect 23750 13404 23756 13416
rect 23808 13404 23814 13456
rect 23842 13404 23848 13456
rect 23900 13444 23906 13456
rect 24121 13447 24179 13453
rect 24121 13444 24133 13447
rect 23900 13416 24133 13444
rect 23900 13404 23906 13416
rect 24121 13413 24133 13416
rect 24167 13413 24179 13447
rect 24121 13407 24179 13413
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13345 23351 13379
rect 23293 13339 23351 13345
rect 23474 13336 23480 13388
rect 23532 13336 23538 13388
rect 10827 13280 11652 13308
rect 10827 13277 10839 13280
rect 10781 13271 10839 13277
rect 7009 13243 7067 13249
rect 6748 13212 6868 13240
rect 4433 13203 4491 13209
rect 3467 13144 3832 13172
rect 3881 13175 3939 13181
rect 3467 13141 3479 13144
rect 3421 13135 3479 13141
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4246 13172 4252 13184
rect 3927 13144 4252 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 4448 13172 4476 13203
rect 6840 13184 6868 13212
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 7098 13240 7104 13252
rect 7055 13212 7104 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 7098 13200 7104 13212
rect 7156 13240 7162 13252
rect 7156 13212 7236 13240
rect 7156 13200 7162 13212
rect 5074 13172 5080 13184
rect 4448 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13172 5138 13184
rect 5810 13172 5816 13184
rect 5132 13144 5816 13172
rect 5132 13132 5138 13144
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 6178 13132 6184 13184
rect 6236 13132 6242 13184
rect 6822 13132 6828 13184
rect 6880 13132 6886 13184
rect 7208 13172 7236 13212
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 9140 13240 9168 13271
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 19978 13308 19984 13320
rect 19260 13280 19984 13308
rect 12253 13243 12311 13249
rect 7340 13212 7498 13240
rect 9140 13212 11744 13240
rect 7340 13200 7346 13212
rect 7926 13172 7932 13184
rect 7208 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9030 13132 9036 13184
rect 9088 13172 9094 13184
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9088 13144 10425 13172
rect 9088 13132 9094 13144
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 10413 13135 10471 13141
rect 10870 13132 10876 13184
rect 10928 13132 10934 13184
rect 11716 13172 11744 13212
rect 12253 13209 12265 13243
rect 12299 13240 12311 13243
rect 12342 13240 12348 13252
rect 12299 13212 12348 13240
rect 12299 13209 12311 13212
rect 12253 13203 12311 13209
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 13262 13200 13268 13252
rect 13320 13200 13326 13252
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17405 13243 17463 13249
rect 17405 13240 17417 13243
rect 17092 13212 17417 13240
rect 17092 13200 17098 13212
rect 17405 13209 17417 13212
rect 17451 13209 17463 13243
rect 17405 13203 17463 13209
rect 18138 13200 18144 13252
rect 18196 13200 18202 13252
rect 14182 13172 14188 13184
rect 11716 13144 14188 13172
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 19260 13172 19288 13280
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 22370 13268 22376 13320
rect 22428 13308 22434 13320
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 22428 13280 22477 13308
rect 22428 13268 22434 13280
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23072 13280 25452 13308
rect 23072 13268 23078 13280
rect 21082 13240 21088 13252
rect 19444 13212 21088 13240
rect 19444 13181 19472 13212
rect 21082 13200 21088 13212
rect 21140 13200 21146 13252
rect 23201 13243 23259 13249
rect 23201 13209 23213 13243
rect 23247 13240 23259 13243
rect 23247 13212 23336 13240
rect 23247 13209 23259 13212
rect 23201 13203 23259 13209
rect 15896 13144 19288 13172
rect 19337 13175 19395 13181
rect 15896 13132 15902 13144
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 19383 13144 19441 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 19429 13141 19441 13144
rect 19475 13141 19487 13175
rect 19429 13135 19487 13141
rect 20346 13132 20352 13184
rect 20404 13172 20410 13184
rect 23106 13172 23112 13184
rect 20404 13144 23112 13172
rect 20404 13132 20410 13144
rect 23106 13132 23112 13144
rect 23164 13132 23170 13184
rect 23308 13172 23336 13212
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 25424 13249 25452 13280
rect 24581 13243 24639 13249
rect 24581 13240 24593 13243
rect 23440 13212 24593 13240
rect 23440 13200 23446 13212
rect 24581 13209 24593 13212
rect 24627 13209 24639 13243
rect 24581 13203 24639 13209
rect 25409 13243 25467 13249
rect 25409 13209 25421 13243
rect 25455 13240 25467 13243
rect 26878 13240 26884 13252
rect 25455 13212 26884 13240
rect 25455 13209 25467 13212
rect 25409 13203 25467 13209
rect 26878 13200 26884 13212
rect 26936 13200 26942 13252
rect 25222 13172 25228 13184
rect 23308 13144 25228 13172
rect 25222 13132 25228 13144
rect 25280 13132 25286 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 3881 12971 3939 12977
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 7190 12968 7196 12980
rect 3927 12940 7196 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 1302 12860 1308 12912
rect 1360 12900 1366 12912
rect 1762 12900 1768 12912
rect 1360 12872 1768 12900
rect 1360 12860 1366 12872
rect 1762 12860 1768 12872
rect 1820 12900 1826 12912
rect 1820 12872 2774 12900
rect 1820 12860 1826 12872
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 2498 12832 2504 12844
rect 1903 12804 2504 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 2746 12832 2774 12872
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2746 12804 2881 12832
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 1118 12724 1124 12776
rect 1176 12764 1182 12776
rect 1581 12767 1639 12773
rect 1581 12764 1593 12767
rect 1176 12736 1593 12764
rect 1176 12724 1182 12736
rect 1581 12733 1593 12736
rect 1627 12764 1639 12767
rect 1670 12764 1676 12776
rect 1627 12736 1676 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 474 12656 480 12708
rect 532 12696 538 12708
rect 3896 12696 3924 12931
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 10594 12968 10600 12980
rect 7331 12940 10600 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 12529 12971 12587 12977
rect 12529 12968 12541 12971
rect 11020 12940 12541 12968
rect 11020 12928 11026 12940
rect 12529 12937 12541 12940
rect 12575 12937 12587 12971
rect 13630 12968 13636 12980
rect 12529 12931 12587 12937
rect 12636 12940 13636 12968
rect 4249 12903 4307 12909
rect 4249 12869 4261 12903
rect 4295 12900 4307 12903
rect 4338 12900 4344 12912
rect 4295 12872 4344 12900
rect 4295 12869 4307 12872
rect 4249 12863 4307 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 4798 12900 4804 12912
rect 4488 12872 4804 12900
rect 4488 12860 4494 12872
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 5721 12903 5779 12909
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 6454 12900 6460 12912
rect 5767 12872 6460 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 7374 12900 7380 12912
rect 6748 12872 7380 12900
rect 6748 12844 6776 12872
rect 7374 12860 7380 12872
rect 7432 12900 7438 12912
rect 8754 12900 8760 12912
rect 7432 12872 8760 12900
rect 7432 12860 7438 12872
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 10045 12903 10103 12909
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 10134 12900 10140 12912
rect 10091 12872 10140 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 12636 12900 12664 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 13722 12928 13728 12980
rect 13780 12928 13786 12980
rect 13998 12928 14004 12980
rect 14056 12968 14062 12980
rect 14182 12968 14188 12980
rect 14056 12940 14188 12968
rect 14056 12928 14062 12940
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 16080 12940 17785 12968
rect 16080 12928 16086 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 18187 12940 19104 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 11931 12872 12664 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 13170 12900 13176 12912
rect 12768 12872 13176 12900
rect 12768 12860 12774 12872
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 13354 12860 13360 12912
rect 13412 12900 13418 12912
rect 14274 12900 14280 12912
rect 13412 12872 14280 12900
rect 13412 12860 13418 12872
rect 14274 12860 14280 12872
rect 14332 12900 14338 12912
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 14332 12872 15669 12900
rect 14332 12860 14338 12872
rect 15657 12869 15669 12872
rect 15703 12869 15715 12903
rect 15657 12863 15715 12869
rect 16114 12860 16120 12912
rect 16172 12860 16178 12912
rect 16393 12903 16451 12909
rect 16393 12869 16405 12903
rect 16439 12900 16451 12903
rect 18414 12900 18420 12912
rect 16439 12872 18420 12900
rect 16439 12869 16451 12872
rect 16393 12863 16451 12869
rect 3970 12792 3976 12844
rect 4028 12832 4034 12844
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 4028 12804 4997 12832
rect 4028 12792 4034 12804
rect 4985 12801 4997 12804
rect 5031 12832 5043 12835
rect 5031 12804 5580 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5166 12764 5172 12776
rect 4856 12736 5172 12764
rect 4856 12724 4862 12736
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5552 12764 5580 12804
rect 5626 12792 5632 12844
rect 5684 12792 5690 12844
rect 6270 12832 6276 12844
rect 5736 12804 6276 12832
rect 5736 12764 5764 12804
rect 6270 12792 6276 12804
rect 6328 12832 6334 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6328 12804 6561 12832
rect 6328 12792 6334 12804
rect 6549 12801 6561 12804
rect 6595 12832 6607 12835
rect 6730 12832 6736 12844
rect 6595 12804 6736 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 6880 12804 7696 12832
rect 6880 12792 6886 12804
rect 5552 12736 5764 12764
rect 5810 12724 5816 12776
rect 5868 12764 5874 12776
rect 5905 12767 5963 12773
rect 5905 12764 5917 12767
rect 5868 12736 5917 12764
rect 5868 12724 5874 12736
rect 5905 12733 5917 12736
rect 5951 12764 5963 12767
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 5951 12736 7389 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 7377 12733 7389 12736
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 532 12668 3924 12696
rect 4433 12699 4491 12705
rect 532 12656 538 12668
rect 4433 12665 4445 12699
rect 4479 12696 4491 12699
rect 7558 12696 7564 12708
rect 4479 12668 7564 12696
rect 4479 12665 4491 12668
rect 4433 12659 4491 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 1854 12588 1860 12640
rect 1912 12628 1918 12640
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 1912 12600 3525 12628
rect 1912 12588 1918 12600
rect 3513 12597 3525 12600
rect 3559 12597 3571 12631
rect 3513 12591 3571 12597
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5442 12628 5448 12640
rect 5307 12600 5448 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 6822 12588 6828 12640
rect 6880 12588 6886 12640
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 7668 12628 7696 12804
rect 10686 12792 10692 12844
rect 10744 12792 10750 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12406 12804 12909 12832
rect 8018 12724 8024 12776
rect 8076 12724 8082 12776
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 9582 12764 9588 12776
rect 8343 12736 9588 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 12406 12764 12434 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13136 12804 14105 12832
rect 13136 12792 13142 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14792 12804 14933 12832
rect 14792 12792 14798 12804
rect 14921 12801 14933 12804
rect 14967 12832 14979 12835
rect 15102 12832 15108 12844
rect 14967 12804 15108 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 15102 12792 15108 12804
rect 15160 12832 15166 12844
rect 16408 12832 16436 12863
rect 18414 12860 18420 12872
rect 18472 12900 18478 12912
rect 18874 12900 18880 12912
rect 18472 12872 18880 12900
rect 18472 12860 18478 12872
rect 18874 12860 18880 12872
rect 18932 12900 18938 12912
rect 18969 12903 19027 12909
rect 18969 12900 18981 12903
rect 18932 12872 18981 12900
rect 18932 12860 18938 12872
rect 18969 12869 18981 12872
rect 19015 12869 19027 12903
rect 19076 12900 19104 12940
rect 19150 12928 19156 12980
rect 19208 12968 19214 12980
rect 20898 12968 20904 12980
rect 19208 12940 20904 12968
rect 19208 12928 19214 12940
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 21174 12968 21180 12980
rect 21131 12940 21180 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 21266 12928 21272 12980
rect 21324 12968 21330 12980
rect 21910 12968 21916 12980
rect 21324 12940 21916 12968
rect 21324 12928 21330 12940
rect 21910 12928 21916 12940
rect 21968 12968 21974 12980
rect 22189 12971 22247 12977
rect 22189 12968 22201 12971
rect 21968 12940 22201 12968
rect 21968 12928 21974 12940
rect 22189 12937 22201 12940
rect 22235 12968 22247 12971
rect 22235 12940 22784 12968
rect 22235 12937 22247 12940
rect 22189 12931 22247 12937
rect 20070 12900 20076 12912
rect 19076 12872 20076 12900
rect 18969 12863 19027 12869
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 22462 12900 22468 12912
rect 21100 12872 22468 12900
rect 15160 12804 16436 12832
rect 15160 12792 15166 12804
rect 17034 12792 17040 12844
rect 17092 12832 17098 12844
rect 17954 12832 17960 12844
rect 17092 12804 17960 12832
rect 17092 12792 17098 12804
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 21100 12832 21128 12872
rect 22462 12860 22468 12872
rect 22520 12860 22526 12912
rect 22756 12900 22784 12940
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 23290 12968 23296 12980
rect 22888 12940 23296 12968
rect 22888 12928 22894 12940
rect 23290 12928 23296 12940
rect 23348 12928 23354 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23532 12940 24777 12968
rect 23532 12928 23538 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 23566 12900 23572 12912
rect 22756 12872 23572 12900
rect 23566 12860 23572 12872
rect 23624 12900 23630 12912
rect 23624 12872 23782 12900
rect 23624 12860 23630 12872
rect 18279 12804 21128 12832
rect 21177 12835 21235 12841
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 21177 12801 21189 12835
rect 21223 12832 21235 12835
rect 21223 12804 22094 12832
rect 21223 12801 21235 12804
rect 21177 12795 21235 12801
rect 10192 12736 12434 12764
rect 12989 12767 13047 12773
rect 10192 12724 10198 12736
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 14369 12767 14427 12773
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 15194 12764 15200 12776
rect 14415 12736 15200 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 10226 12656 10232 12708
rect 10284 12696 10290 12708
rect 10505 12699 10563 12705
rect 10505 12696 10517 12699
rect 10284 12668 10517 12696
rect 10284 12656 10290 12668
rect 10505 12665 10517 12668
rect 10551 12665 10563 12699
rect 10505 12659 10563 12665
rect 11149 12699 11207 12705
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 12250 12696 12256 12708
rect 11195 12668 12256 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 12250 12656 12256 12668
rect 12308 12656 12314 12708
rect 7432 12600 7696 12628
rect 7432 12588 7438 12600
rect 8754 12588 8760 12640
rect 8812 12628 8818 12640
rect 9490 12628 9496 12640
rect 8812 12600 9496 12628
rect 8812 12588 8818 12600
rect 9490 12588 9496 12600
rect 9548 12628 9554 12640
rect 11241 12631 11299 12637
rect 11241 12628 11253 12631
rect 9548 12600 11253 12628
rect 9548 12588 9554 12600
rect 11241 12597 11253 12600
rect 11287 12597 11299 12631
rect 11241 12591 11299 12597
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 11388 12600 11621 12628
rect 11388 12588 11394 12600
rect 11609 12597 11621 12600
rect 11655 12628 11667 12631
rect 12158 12628 12164 12640
rect 11655 12600 12164 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 12158 12588 12164 12600
rect 12216 12628 12222 12640
rect 12894 12628 12900 12640
rect 12216 12600 12900 12628
rect 12216 12588 12222 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13004 12628 13032 12727
rect 13188 12696 13216 12727
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15344 12736 16865 12764
rect 15344 12724 15350 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 18414 12724 18420 12776
rect 18472 12724 18478 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20070 12764 20076 12776
rect 19843 12736 20076 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 15470 12696 15476 12708
rect 13188 12668 15476 12696
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 17494 12656 17500 12708
rect 17552 12696 17558 12708
rect 19812 12696 19840 12727
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 22066 12764 22094 12804
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 23014 12832 23020 12844
rect 22244 12804 23020 12832
rect 22244 12792 22250 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 22646 12764 22652 12776
rect 22066 12736 22652 12764
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 23658 12764 23664 12776
rect 23339 12736 23664 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 17552 12668 19840 12696
rect 17552 12656 17558 12668
rect 17862 12628 17868 12640
rect 13004 12600 17868 12628
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 19484 12600 20729 12628
rect 19484 12588 19490 12600
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 23658 12588 23664 12640
rect 23716 12628 23722 12640
rect 25041 12631 25099 12637
rect 25041 12628 25053 12631
rect 23716 12600 25053 12628
rect 23716 12588 23722 12600
rect 25041 12597 25053 12600
rect 25087 12597 25099 12631
rect 25041 12591 25099 12597
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3053 12427 3111 12433
rect 3053 12424 3065 12427
rect 2832 12396 3065 12424
rect 2832 12384 2838 12396
rect 3053 12393 3065 12396
rect 3099 12393 3111 12427
rect 3053 12387 3111 12393
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 3970 12424 3976 12436
rect 3559 12396 3976 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 4396 12396 4721 12424
rect 4396 12384 4402 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 4709 12387 4767 12393
rect 4798 12384 4804 12436
rect 4856 12424 4862 12436
rect 6086 12424 6092 12436
rect 4856 12396 6092 12424
rect 4856 12384 4862 12396
rect 6086 12384 6092 12396
rect 6144 12384 6150 12436
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 7742 12424 7748 12436
rect 7616 12396 7748 12424
rect 7616 12384 7622 12396
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 10870 12424 10876 12436
rect 7883 12396 10876 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 11606 12424 11612 12436
rect 11296 12396 11612 12424
rect 11296 12384 11302 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11793 12427 11851 12433
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 12526 12424 12532 12436
rect 11839 12396 12532 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 12710 12384 12716 12436
rect 12768 12424 12774 12436
rect 13722 12424 13728 12436
rect 12768 12396 13728 12424
rect 12768 12384 12774 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14240 12396 14381 12424
rect 14240 12384 14246 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 14550 12384 14556 12436
rect 14608 12424 14614 12436
rect 14608 12396 17632 12424
rect 14608 12384 14614 12396
rect 4249 12359 4307 12365
rect 4249 12325 4261 12359
rect 4295 12356 4307 12359
rect 4982 12356 4988 12368
rect 4295 12328 4988 12356
rect 4295 12325 4307 12328
rect 4249 12319 4307 12325
rect 4982 12316 4988 12328
rect 5040 12316 5046 12368
rect 7374 12316 7380 12368
rect 7432 12356 7438 12368
rect 8018 12356 8024 12368
rect 7432 12328 8024 12356
rect 7432 12316 7438 12328
rect 8018 12316 8024 12328
rect 8076 12356 8082 12368
rect 8076 12328 9352 12356
rect 8076 12316 8082 12328
rect 9324 12300 9352 12328
rect 9766 12316 9772 12368
rect 9824 12356 9830 12368
rect 9824 12328 10916 12356
rect 9824 12316 9830 12328
rect 10888 12300 10916 12328
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 13446 12356 13452 12368
rect 11020 12328 13452 12356
rect 11020 12316 11026 12328
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 15286 12356 15292 12368
rect 13556 12328 15292 12356
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 4212 12260 5365 12288
rect 4212 12248 4218 12260
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 7156 12260 8401 12288
rect 7156 12248 7162 12260
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9364 12260 9873 12288
rect 9364 12248 9370 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 10870 12248 10876 12300
rect 10928 12248 10934 12300
rect 11238 12248 11244 12300
rect 11296 12248 11302 12300
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 12158 12288 12164 12300
rect 11388 12260 12164 12288
rect 11388 12248 11394 12260
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12250 12248 12256 12300
rect 12308 12248 12314 12300
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 1578 12180 1584 12232
rect 1636 12180 1642 12232
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 4338 12220 4344 12232
rect 1903 12192 4344 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 4338 12180 4344 12192
rect 4396 12220 4402 12232
rect 4798 12220 4804 12232
rect 4396 12192 4804 12220
rect 4396 12180 4402 12192
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 4890 12180 4896 12232
rect 4948 12180 4954 12232
rect 6730 12180 6736 12232
rect 6788 12180 6794 12232
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12220 7435 12223
rect 7466 12220 7472 12232
rect 7423 12192 7472 12220
rect 7423 12189 7435 12192
rect 7377 12183 7435 12189
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 10410 12220 10416 12232
rect 8343 12192 10416 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12220 11115 12223
rect 13262 12220 13268 12232
rect 11103 12192 13268 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 13556 12220 13584 12328
rect 15286 12316 15292 12328
rect 15344 12316 15350 12368
rect 15470 12316 15476 12368
rect 15528 12356 15534 12368
rect 17604 12356 17632 12396
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18049 12427 18107 12433
rect 18049 12424 18061 12427
rect 18012 12396 18061 12424
rect 18012 12384 18018 12396
rect 18049 12393 18061 12396
rect 18095 12424 18107 12427
rect 19150 12424 19156 12436
rect 18095 12396 19156 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21821 12427 21879 12433
rect 21821 12424 21833 12427
rect 20772 12396 21833 12424
rect 20772 12384 20778 12396
rect 21821 12393 21833 12396
rect 21867 12424 21879 12427
rect 21867 12396 22094 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 19518 12356 19524 12368
rect 15528 12328 16252 12356
rect 17604 12328 19524 12356
rect 15528 12316 15534 12328
rect 16224 12300 16252 12328
rect 19518 12316 19524 12328
rect 19576 12316 19582 12368
rect 19812 12328 20208 12356
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 15838 12288 15844 12300
rect 13679 12260 15844 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 16206 12248 16212 12300
rect 16264 12288 16270 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16264 12260 16589 12288
rect 16264 12248 16270 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 18782 12288 18788 12300
rect 16577 12251 16635 12257
rect 18524 12260 18788 12288
rect 13403 12192 13584 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13780 12192 14105 12220
rect 13780 12180 13786 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 14516 12192 15485 12220
rect 14516 12180 14522 12192
rect 15473 12189 15485 12192
rect 15519 12220 15531 12223
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 15519 12192 16313 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 17710 12192 18337 12220
rect 16301 12183 16359 12189
rect 18325 12189 18337 12192
rect 18371 12220 18383 12223
rect 18524 12220 18552 12260
rect 18782 12248 18788 12260
rect 18840 12288 18846 12300
rect 19061 12291 19119 12297
rect 19061 12288 19073 12291
rect 18840 12260 19073 12288
rect 18840 12248 18846 12260
rect 19061 12257 19073 12260
rect 19107 12288 19119 12291
rect 19812 12288 19840 12328
rect 19107 12260 19840 12288
rect 19107 12257 19119 12260
rect 19061 12251 19119 12257
rect 20070 12248 20076 12300
rect 20128 12248 20134 12300
rect 20180 12288 20208 12328
rect 22066 12288 22094 12396
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 20180 12260 21588 12288
rect 22066 12260 22569 12288
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 18371 12192 18552 12220
rect 18616 12192 19533 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 2590 12112 2596 12164
rect 2648 12152 2654 12164
rect 2866 12152 2872 12164
rect 2648 12124 2872 12152
rect 2648 12112 2654 12124
rect 2866 12112 2872 12124
rect 2924 12152 2930 12164
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2924 12124 2973 12152
rect 2924 12112 2930 12124
rect 2961 12121 2973 12124
rect 3007 12121 3019 12155
rect 2961 12115 3019 12121
rect 3970 12112 3976 12164
rect 4028 12152 4034 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 4028 12124 4077 12152
rect 4028 12112 4034 12124
rect 4065 12121 4077 12124
rect 4111 12152 4123 12155
rect 5534 12152 5540 12164
rect 4111 12124 5540 12152
rect 4111 12121 4123 12124
rect 4065 12115 4123 12121
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 5629 12155 5687 12161
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 5718 12152 5724 12164
rect 5675 12124 5724 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 9122 12112 9128 12164
rect 9180 12112 9186 12164
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 9364 12124 10977 12152
rect 9364 12112 9370 12124
rect 10965 12121 10977 12124
rect 11011 12121 11023 12155
rect 10965 12115 11023 12121
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 12161 12155 12219 12161
rect 12161 12152 12173 12155
rect 11940 12124 12173 12152
rect 11940 12112 11946 12124
rect 12161 12121 12173 12124
rect 12207 12121 12219 12155
rect 12161 12115 12219 12121
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13449 12155 13507 12161
rect 13449 12152 13461 12155
rect 12952 12124 13461 12152
rect 12952 12112 12958 12124
rect 13449 12121 13461 12124
rect 13495 12121 13507 12155
rect 14550 12152 14556 12164
rect 13449 12115 13507 12121
rect 14016 12124 14556 12152
rect 6270 12044 6276 12096
rect 6328 12084 6334 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 6328 12056 8217 12084
rect 6328 12044 6334 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8846 12084 8852 12096
rect 8352 12056 8852 12084
rect 8352 12044 8358 12056
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 11974 12084 11980 12096
rect 11756 12056 11980 12084
rect 11756 12044 11762 12056
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 14016 12084 14044 12124
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 14754 12155 14812 12161
rect 14754 12121 14766 12155
rect 14800 12152 14812 12155
rect 18616 12152 18644 12192
rect 19521 12189 19533 12192
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 14800 12124 14964 12152
rect 14800 12121 14812 12124
rect 14754 12115 14812 12121
rect 14936 12096 14964 12124
rect 17880 12124 18644 12152
rect 13035 12056 14044 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 14918 12044 14924 12096
rect 14976 12084 14982 12096
rect 15933 12087 15991 12093
rect 15933 12084 15945 12087
rect 14976 12056 15945 12084
rect 14976 12044 14982 12056
rect 15933 12053 15945 12056
rect 15979 12053 15991 12087
rect 15933 12047 15991 12053
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 17880 12084 17908 12124
rect 17460 12056 17908 12084
rect 17460 12044 17466 12056
rect 18414 12044 18420 12096
rect 18472 12084 18478 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 18472 12056 18521 12084
rect 18472 12044 18478 12056
rect 18509 12053 18521 12056
rect 18555 12084 18567 12087
rect 18690 12084 18696 12096
rect 18555 12056 18696 12084
rect 18555 12053 18567 12056
rect 18509 12047 18567 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 18874 12084 18880 12096
rect 18831 12056 18880 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 18874 12044 18880 12056
rect 18932 12084 18938 12096
rect 19242 12084 19248 12096
rect 18932 12056 19248 12084
rect 18932 12044 18938 12056
rect 19242 12044 19248 12056
rect 19300 12084 19306 12096
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 19300 12056 19349 12084
rect 19300 12044 19306 12056
rect 19337 12053 19349 12056
rect 19383 12053 19395 12087
rect 19536 12084 19564 12183
rect 20346 12112 20352 12164
rect 20404 12112 20410 12164
rect 21560 12152 21588 12260
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22244 12192 22293 12220
rect 22244 12180 22250 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 23658 12180 23664 12232
rect 23716 12220 23722 12232
rect 23934 12220 23940 12232
rect 23716 12192 23940 12220
rect 23716 12180 23722 12192
rect 23934 12180 23940 12192
rect 23992 12180 23998 12232
rect 21910 12152 21916 12164
rect 21560 12138 21916 12152
rect 21574 12124 21916 12138
rect 21910 12112 21916 12124
rect 21968 12112 21974 12164
rect 25038 12152 25044 12164
rect 23860 12124 25044 12152
rect 23860 12084 23888 12124
rect 25038 12112 25044 12124
rect 25096 12112 25102 12164
rect 19536 12056 23888 12084
rect 19337 12047 19395 12053
rect 24026 12044 24032 12096
rect 24084 12044 24090 12096
rect 24489 12087 24547 12093
rect 24489 12053 24501 12087
rect 24535 12084 24547 12087
rect 24670 12084 24676 12096
rect 24535 12056 24676 12084
rect 24535 12053 24547 12056
rect 24489 12047 24547 12053
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 2225 11883 2283 11889
rect 2225 11880 2237 11883
rect 1636 11852 2237 11880
rect 1636 11840 1642 11852
rect 2225 11849 2237 11852
rect 2271 11849 2283 11883
rect 2225 11843 2283 11849
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3602 11880 3608 11892
rect 3016 11852 3608 11880
rect 3016 11840 3022 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4479 11852 5273 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5500 11852 5641 11880
rect 5500 11840 5506 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 12345 11883 12403 11889
rect 12345 11880 12357 11883
rect 6779 11852 12357 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 12345 11849 12357 11852
rect 12391 11849 12403 11883
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 12345 11843 12403 11849
rect 13096 11852 14933 11880
rect 1302 11772 1308 11824
rect 1360 11812 1366 11824
rect 3789 11815 3847 11821
rect 1360 11784 2728 11812
rect 1360 11772 1366 11784
rect 1118 11704 1124 11756
rect 1176 11744 1182 11756
rect 1394 11744 1400 11756
rect 1176 11716 1400 11744
rect 1176 11704 1182 11716
rect 1394 11704 1400 11716
rect 1452 11744 1458 11756
rect 2700 11753 2728 11784
rect 3789 11781 3801 11815
rect 3835 11812 3847 11815
rect 4614 11812 4620 11824
rect 3835 11784 4620 11812
rect 3835 11781 3847 11784
rect 3789 11775 3847 11781
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1452 11716 1593 11744
rect 1452 11704 1458 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11744 2743 11747
rect 3418 11744 3424 11756
rect 2731 11716 3424 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 3804 11676 3832 11775
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 5721 11815 5779 11821
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 6822 11812 6828 11824
rect 5767 11784 6828 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 8110 11772 8116 11824
rect 8168 11772 8174 11824
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 9490 11812 9496 11824
rect 9088 11784 9496 11812
rect 9088 11772 9094 11784
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 10594 11772 10600 11824
rect 10652 11812 10658 11824
rect 12437 11815 12495 11821
rect 12437 11812 12449 11815
rect 10652 11784 12449 11812
rect 10652 11772 10658 11784
rect 12437 11781 12449 11784
rect 12483 11781 12495 11815
rect 12437 11775 12495 11781
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 5258 11744 5264 11756
rect 4571 11716 5264 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9180 11716 9597 11744
rect 9180 11704 9186 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9692 11716 10640 11744
rect 2556 11648 3832 11676
rect 4709 11679 4767 11685
rect 2556 11636 2562 11648
rect 4709 11645 4721 11679
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 4724 11608 4752 11639
rect 5902 11636 5908 11688
rect 5960 11636 5966 11688
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 8386 11676 8392 11688
rect 7699 11648 8392 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8846 11636 8852 11688
rect 8904 11676 8910 11688
rect 9692 11676 9720 11716
rect 8904 11648 9720 11676
rect 8904 11636 8910 11648
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 9916 11648 10333 11676
rect 9916 11636 9922 11648
rect 10321 11645 10333 11648
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 9125 11611 9183 11617
rect 4724 11580 5764 11608
rect 5736 11552 5764 11580
rect 9125 11577 9137 11611
rect 9171 11608 9183 11611
rect 9582 11608 9588 11620
rect 9171 11580 9588 11608
rect 9171 11577 9183 11580
rect 9125 11571 9183 11577
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3329 11543 3387 11549
rect 3329 11540 3341 11543
rect 2832 11512 3341 11540
rect 2832 11500 2838 11512
rect 3329 11509 3341 11512
rect 3375 11509 3387 11543
rect 3329 11503 3387 11509
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 5534 11540 5540 11552
rect 4111 11512 5540 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5718 11500 5724 11552
rect 5776 11500 5782 11552
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 9398 11540 9404 11552
rect 6420 11512 9404 11540
rect 6420 11500 6426 11512
rect 9398 11500 9404 11512
rect 9456 11540 9462 11552
rect 10502 11540 10508 11552
rect 9456 11512 10508 11540
rect 9456 11500 9462 11512
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 10612 11540 10640 11716
rect 10962 11704 10968 11756
rect 11020 11704 11026 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 12066 11744 12072 11756
rect 11296 11716 12072 11744
rect 11296 11704 11302 11716
rect 12066 11704 12072 11716
rect 12124 11744 12130 11756
rect 13096 11744 13124 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 14921 11843 14979 11849
rect 17402 11840 17408 11892
rect 17460 11840 17466 11892
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 18141 11883 18199 11889
rect 18141 11880 18153 11883
rect 17920 11852 18153 11880
rect 17920 11840 17926 11852
rect 18141 11849 18153 11852
rect 18187 11849 18199 11883
rect 18141 11843 18199 11849
rect 18506 11840 18512 11892
rect 18564 11840 18570 11892
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 19337 11883 19395 11889
rect 19337 11880 19349 11883
rect 18656 11852 19349 11880
rect 18656 11840 18662 11852
rect 19337 11849 19349 11852
rect 19383 11849 19395 11883
rect 32398 11880 32404 11892
rect 19337 11843 19395 11849
rect 19536 11852 32404 11880
rect 13354 11812 13360 11824
rect 13188 11784 13360 11812
rect 13188 11753 13216 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 15286 11812 15292 11824
rect 14674 11784 15292 11812
rect 15286 11772 15292 11784
rect 15344 11772 15350 11824
rect 16025 11815 16083 11821
rect 16025 11781 16037 11815
rect 16071 11812 16083 11815
rect 18524 11812 18552 11840
rect 19153 11815 19211 11821
rect 19153 11812 19165 11815
rect 16071 11784 17724 11812
rect 18524 11784 19165 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 12124 11716 13124 11744
rect 13173 11747 13231 11753
rect 12124 11704 12130 11716
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 15930 11704 15936 11756
rect 15988 11704 15994 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 16132 11716 17325 11744
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 11848 11648 12541 11676
rect 11848 11636 11854 11648
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 15010 11676 15016 11688
rect 13495 11648 15016 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 16132 11676 16160 11716
rect 17313 11713 17325 11716
rect 17359 11744 17371 11747
rect 17696 11744 17724 11784
rect 19153 11781 19165 11784
rect 19199 11781 19211 11815
rect 19153 11775 19211 11781
rect 19426 11744 19432 11756
rect 17359 11716 17632 11744
rect 17696 11716 19432 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 15120 11648 16160 11676
rect 16209 11679 16267 11685
rect 10870 11568 10876 11620
rect 10928 11608 10934 11620
rect 11609 11611 11667 11617
rect 11609 11608 11621 11611
rect 10928 11580 11621 11608
rect 10928 11568 10934 11580
rect 11609 11577 11621 11580
rect 11655 11608 11667 11611
rect 12894 11608 12900 11620
rect 11655 11580 12900 11608
rect 11655 11577 11667 11580
rect 11609 11571 11667 11577
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 10612 11512 11989 11540
rect 11977 11509 11989 11512
rect 12023 11509 12035 11543
rect 11977 11503 12035 11509
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 15120 11540 15148 11648
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 17034 11676 17040 11688
rect 16255 11648 17040 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 17034 11636 17040 11648
rect 17092 11636 17098 11688
rect 17402 11636 17408 11688
rect 17460 11676 17466 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 17460 11648 17509 11676
rect 17460 11636 17466 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17604 11676 17632 11716
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 18414 11676 18420 11688
rect 17604 11648 18420 11676
rect 17497 11639 17555 11645
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 18690 11636 18696 11688
rect 18748 11636 18754 11688
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 19536 11676 19564 11852
rect 32398 11840 32404 11852
rect 32456 11840 32462 11892
rect 21910 11812 21916 11824
rect 21206 11784 21916 11812
rect 21910 11772 21916 11784
rect 21968 11772 21974 11824
rect 22649 11815 22707 11821
rect 22649 11781 22661 11815
rect 22695 11812 22707 11815
rect 22738 11812 22744 11824
rect 22695 11784 22744 11812
rect 22695 11781 22707 11784
rect 22649 11775 22707 11781
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 23934 11812 23940 11824
rect 23874 11784 23940 11812
rect 23934 11772 23940 11784
rect 23992 11812 23998 11824
rect 24670 11812 24676 11824
rect 23992 11784 24676 11812
rect 23992 11772 23998 11784
rect 24670 11772 24676 11784
rect 24728 11772 24734 11824
rect 18840 11648 19564 11676
rect 18840 11636 18846 11648
rect 19702 11636 19708 11688
rect 19760 11636 19766 11688
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11676 20039 11679
rect 20027 11648 22094 11676
rect 20027 11645 20039 11648
rect 19981 11639 20039 11645
rect 15565 11611 15623 11617
rect 15565 11577 15577 11611
rect 15611 11608 15623 11611
rect 19150 11608 19156 11620
rect 15611 11580 19156 11608
rect 15611 11577 15623 11580
rect 15565 11571 15623 11577
rect 19150 11568 19156 11580
rect 19208 11568 19214 11620
rect 22066 11608 22094 11648
rect 22186 11636 22192 11688
rect 22244 11676 22250 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 22244 11648 22385 11676
rect 22244 11636 22250 11648
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 24026 11676 24032 11688
rect 22373 11639 22431 11645
rect 22480 11648 24032 11676
rect 22480 11608 22508 11648
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 24121 11679 24179 11685
rect 24121 11645 24133 11679
rect 24167 11676 24179 11679
rect 25130 11676 25136 11688
rect 24167 11648 25136 11676
rect 24167 11645 24179 11648
rect 24121 11639 24179 11645
rect 22066 11580 22508 11608
rect 12308 11512 15148 11540
rect 12308 11500 12314 11512
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16114 11540 16120 11552
rect 15344 11512 16120 11540
rect 15344 11500 15350 11512
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 16942 11500 16948 11552
rect 17000 11500 17006 11552
rect 21450 11500 21456 11552
rect 21508 11500 21514 11552
rect 21634 11500 21640 11552
rect 21692 11540 21698 11552
rect 24136 11540 24164 11639
rect 25130 11636 25136 11648
rect 25188 11636 25194 11688
rect 21692 11512 24164 11540
rect 24489 11543 24547 11549
rect 21692 11500 21698 11512
rect 24489 11509 24501 11543
rect 24535 11540 24547 11543
rect 24670 11540 24676 11552
rect 24535 11512 24676 11540
rect 24535 11509 24547 11512
rect 24489 11503 24547 11509
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 1489 11339 1547 11345
rect 1489 11305 1501 11339
rect 1535 11336 1547 11339
rect 1578 11336 1584 11348
rect 1535 11308 1584 11336
rect 1535 11305 1547 11308
rect 1489 11299 1547 11305
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1719 11308 2774 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 2746 11268 2774 11308
rect 3878 11296 3884 11348
rect 3936 11296 3942 11348
rect 4890 11296 4896 11348
rect 4948 11296 4954 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 5776 11308 6561 11336
rect 5776 11296 5782 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 6788 11308 7481 11336
rect 6788 11296 6794 11308
rect 7469 11305 7481 11308
rect 7515 11336 7527 11339
rect 8110 11336 8116 11348
rect 7515 11308 8116 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 8110 11296 8116 11308
rect 8168 11336 8174 11348
rect 9125 11339 9183 11345
rect 8168 11308 8892 11336
rect 8168 11296 8174 11308
rect 4908 11268 4936 11296
rect 2746 11240 4936 11268
rect 1946 11160 1952 11212
rect 2004 11160 2010 11212
rect 4154 11160 4160 11212
rect 4212 11160 4218 11212
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5810 11200 5816 11212
rect 5123 11172 5816 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6748 11200 6776 11296
rect 8864 11280 8892 11308
rect 9125 11305 9137 11339
rect 9171 11336 9183 11339
rect 11330 11336 11336 11348
rect 9171 11308 11336 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 12400 11308 13277 11336
rect 12400 11296 12406 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 14369 11339 14427 11345
rect 13412 11308 14136 11336
rect 13412 11296 13418 11308
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7156 11240 8432 11268
rect 7156 11228 7162 11240
rect 6196 11172 6776 11200
rect 7009 11203 7067 11209
rect 2590 11092 2596 11144
rect 2648 11092 2654 11144
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 2884 11064 2912 11095
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 6196 11118 6224 11172
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7190 11200 7196 11212
rect 7055 11172 7196 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8404 11209 8432 11240
rect 8846 11228 8852 11280
rect 8904 11228 8910 11280
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 14108 11277 14136 11308
rect 14369 11305 14381 11339
rect 14415 11336 14427 11339
rect 14642 11336 14648 11348
rect 14415 11308 14648 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 14844 11308 16068 11336
rect 13541 11271 13599 11277
rect 13541 11268 13553 11271
rect 12860 11240 13553 11268
rect 12860 11228 12866 11240
rect 13541 11237 13553 11240
rect 13587 11237 13599 11271
rect 13541 11231 13599 11237
rect 14093 11271 14151 11277
rect 14093 11237 14105 11271
rect 14139 11268 14151 11271
rect 14844 11268 14872 11308
rect 14139 11240 14872 11268
rect 16040 11268 16068 11308
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 16264 11308 16497 11336
rect 16264 11296 16270 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 18877 11339 18935 11345
rect 16485 11299 16543 11305
rect 16592 11308 18460 11336
rect 16592 11268 16620 11308
rect 16040 11240 16620 11268
rect 18432 11268 18460 11308
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 18966 11336 18972 11348
rect 18923 11308 18972 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 20990 11336 20996 11348
rect 19306 11308 20996 11336
rect 19306 11268 19334 11308
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 22646 11296 22652 11348
rect 22704 11336 22710 11348
rect 23290 11336 23296 11348
rect 22704 11308 23296 11336
rect 22704 11296 22710 11308
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 18432 11240 19334 11268
rect 23017 11271 23075 11277
rect 14139 11237 14151 11240
rect 14093 11231 14151 11237
rect 23017 11237 23029 11271
rect 23063 11268 23075 11271
rect 24302 11268 24308 11280
rect 23063 11240 24308 11268
rect 23063 11237 23075 11240
rect 23017 11231 23075 11237
rect 24302 11228 24308 11240
rect 24360 11268 24366 11280
rect 24670 11268 24676 11280
rect 24360 11240 24676 11268
rect 24360 11228 24366 11240
rect 24670 11228 24676 11240
rect 24728 11268 24734 11280
rect 24728 11240 29868 11268
rect 24728 11228 24734 11240
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 7892 11172 8309 11200
rect 7892 11160 7898 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 9214 11160 9220 11212
rect 9272 11200 9278 11212
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9272 11172 9597 11200
rect 9272 11160 9278 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 9674 11160 9680 11212
rect 9732 11160 9738 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11011 11172 11805 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11793 11169 11805 11172
rect 11839 11200 11851 11203
rect 13354 11200 13360 11212
rect 11839 11172 13360 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 14182 11160 14188 11212
rect 14240 11200 14246 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14240 11172 15025 11200
rect 14240 11160 14246 11172
rect 15013 11169 15025 11172
rect 15059 11200 15071 11203
rect 18690 11200 18696 11212
rect 15059 11172 18696 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 18690 11160 18696 11172
rect 18748 11160 18754 11212
rect 26878 11160 26884 11212
rect 26936 11200 26942 11212
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 26936 11172 29745 11200
rect 26936 11160 26942 11172
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29840 11200 29868 11240
rect 32033 11203 32091 11209
rect 32033 11200 32045 11203
rect 29840 11172 32045 11200
rect 29733 11163 29791 11169
rect 7466 11132 7472 11144
rect 6380 11104 7472 11132
rect 2884 11036 5488 11064
rect 5460 10996 5488 11036
rect 6380 10996 6408 11104
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8478 11132 8484 11144
rect 8251 11104 8484 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 9916 11104 11529 11132
rect 9916 11092 9922 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 13722 11132 13728 11144
rect 12926 11104 13728 11132
rect 11517 11095 11575 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14516 11104 14749 11132
rect 14516 11092 14522 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 16114 11092 16120 11144
rect 16172 11092 16178 11144
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16908 11104 17141 11132
rect 16908 11092 16914 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 19242 11092 19248 11144
rect 19300 11132 19306 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 19300 11104 19533 11132
rect 19300 11092 19306 11104
rect 19521 11101 19533 11104
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 31128 11118 31156 11172
rect 32033 11169 32045 11172
rect 32079 11169 32091 11203
rect 32033 11163 32091 11169
rect 20901 11095 20959 11101
rect 7852 11036 9720 11064
rect 7852 11005 7880 11036
rect 5460 10968 6408 10996
rect 7837 10999 7895 11005
rect 7837 10965 7849 10999
rect 7883 10965 7895 10999
rect 9692 10996 9720 11036
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 9824 11036 10701 11064
rect 9824 11024 9830 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10689 11027 10747 11033
rect 13648 11036 14228 11064
rect 9950 10996 9956 11008
rect 9692 10968 9956 10996
rect 7837 10959 7895 10965
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 10318 10956 10324 11008
rect 10376 10956 10382 11008
rect 10778 10956 10784 11008
rect 10836 10956 10842 11008
rect 10962 10956 10968 11008
rect 11020 10996 11026 11008
rect 13648 10996 13676 11036
rect 11020 10968 13676 10996
rect 11020 10956 11026 10968
rect 13814 10956 13820 11008
rect 13872 10956 13878 11008
rect 14200 10996 14228 11036
rect 15286 10996 15292 11008
rect 14200 10968 15292 10996
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 16132 10996 16160 11092
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17405 11067 17463 11073
rect 17405 11064 17417 11067
rect 17368 11036 17417 11064
rect 17368 11024 17374 11036
rect 17405 11033 17417 11036
rect 17451 11064 17463 11067
rect 17678 11064 17684 11076
rect 17451 11036 17684 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 17678 11024 17684 11036
rect 17736 11064 17742 11076
rect 18874 11064 18880 11076
rect 17736 11036 17816 11064
rect 18630 11036 18880 11064
rect 17736 11024 17742 11036
rect 16758 10996 16764 11008
rect 16132 10968 16764 10996
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 17788 10996 17816 11036
rect 18874 11024 18880 11036
rect 18932 11024 18938 11076
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 19760 11036 20269 11064
rect 19760 11024 19766 11036
rect 20257 11033 20269 11036
rect 20303 11064 20315 11067
rect 20916 11064 20944 11095
rect 31294 11092 31300 11144
rect 31352 11132 31358 11144
rect 31757 11135 31815 11141
rect 31757 11132 31769 11135
rect 31352 11104 31769 11132
rect 31352 11092 31358 11104
rect 31757 11101 31769 11104
rect 31803 11132 31815 11135
rect 47578 11132 47584 11144
rect 31803 11104 47584 11132
rect 31803 11101 31815 11104
rect 31757 11095 31815 11101
rect 47578 11092 47584 11104
rect 47636 11092 47642 11144
rect 20303 11036 20944 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 21910 11024 21916 11076
rect 21968 11024 21974 11076
rect 27614 11024 27620 11076
rect 27672 11064 27678 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 27672 11036 30021 11064
rect 27672 11024 27678 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 21358 10996 21364 11008
rect 17788 10968 21364 10996
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1762 10752 1768 10804
rect 1820 10752 1826 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 9861 10795 9919 10801
rect 5859 10764 9076 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 1673 10727 1731 10733
rect 1673 10693 1685 10727
rect 1719 10724 1731 10727
rect 2038 10724 2044 10736
rect 1719 10696 2044 10724
rect 1719 10693 1731 10696
rect 1673 10687 1731 10693
rect 2038 10684 2044 10696
rect 2096 10684 2102 10736
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 8018 10724 8024 10736
rect 6328 10696 8024 10724
rect 6328 10684 6334 10696
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 9048 10724 9076 10764
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 14734 10792 14740 10804
rect 9907 10764 14740 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 15436 10764 15577 10792
rect 15436 10752 15442 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 15565 10755 15623 10761
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 17092 10764 19257 10792
rect 17092 10752 17098 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 21450 10792 21456 10804
rect 19245 10755 19303 10761
rect 19536 10764 21456 10792
rect 10689 10727 10747 10733
rect 10689 10724 10701 10727
rect 9048 10696 10701 10724
rect 10689 10693 10701 10696
rect 10735 10693 10747 10727
rect 10689 10687 10747 10693
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 11422 10724 11428 10736
rect 10827 10696 11428 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 11422 10684 11428 10696
rect 11480 10684 11486 10736
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12345 10727 12403 10733
rect 12345 10724 12357 10727
rect 12124 10696 12357 10724
rect 12124 10684 12130 10696
rect 12345 10693 12357 10696
rect 12391 10693 12403 10727
rect 13814 10724 13820 10736
rect 13570 10696 13820 10724
rect 12345 10687 12403 10693
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 16942 10724 16948 10736
rect 14875 10696 16948 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 658 10616 664 10668
rect 716 10656 722 10668
rect 2409 10659 2467 10665
rect 2409 10656 2421 10659
rect 716 10628 2421 10656
rect 716 10616 722 10628
rect 2409 10625 2421 10628
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 4246 10616 4252 10668
rect 4304 10656 4310 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4304 10628 4721 10656
rect 4304 10616 4310 10628
rect 4709 10625 4721 10628
rect 4755 10656 4767 10659
rect 5350 10656 5356 10668
rect 4755 10628 5356 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 7006 10616 7012 10668
rect 7064 10616 7070 10668
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 9456 10628 9505 10656
rect 9456 10616 9462 10628
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 11609 10659 11667 10665
rect 11609 10656 11621 10659
rect 9732 10628 11621 10656
rect 9732 10616 9738 10628
rect 11609 10625 11621 10628
rect 11655 10656 11667 10659
rect 11882 10656 11888 10668
rect 11655 10628 11888 10656
rect 11655 10625 11667 10628
rect 11609 10619 11667 10625
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 2087 10560 2145 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2133 10557 2145 10560
rect 2179 10588 2191 10591
rect 3234 10588 3240 10600
rect 2179 10560 3240 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 6914 10588 6920 10600
rect 3743 10560 6920 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 1489 10523 1547 10529
rect 1489 10489 1501 10523
rect 1535 10520 1547 10523
rect 2866 10520 2872 10532
rect 1535 10492 2872 10520
rect 1535 10489 1547 10492
rect 1489 10483 1547 10489
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 3436 10520 3464 10551
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7745 10591 7803 10597
rect 7515 10560 7604 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 5258 10520 5264 10532
rect 3436 10492 5264 10520
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 4338 10412 4344 10464
rect 4396 10452 4402 10464
rect 5353 10455 5411 10461
rect 5353 10452 5365 10455
rect 4396 10424 5365 10452
rect 4396 10412 4402 10424
rect 5353 10421 5365 10424
rect 5399 10421 5411 10455
rect 5353 10415 5411 10421
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6328 10424 6469 10452
rect 6328 10412 6334 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6604 10424 6837 10452
rect 6604 10412 6610 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 7576 10452 7604 10560
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8110 10588 8116 10600
rect 7791 10560 8116 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 10045 10591 10103 10597
rect 8260 10560 8800 10588
rect 8260 10548 8266 10560
rect 8772 10520 8800 10560
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 10686 10588 10692 10600
rect 10091 10560 10692 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11296 10560 12081 10588
rect 11296 10548 11302 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 14752 10588 14780 10619
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 14976 10628 15945 10656
rect 14976 10616 14982 10628
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 12492 10560 14780 10588
rect 15013 10591 15071 10597
rect 12492 10548 12498 10560
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15194 10588 15200 10600
rect 15059 10560 15200 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 10321 10523 10379 10529
rect 10321 10520 10333 10523
rect 8772 10492 10333 10520
rect 10321 10489 10333 10492
rect 10367 10489 10379 10523
rect 10321 10483 10379 10489
rect 14369 10523 14427 10529
rect 14369 10489 14381 10523
rect 14415 10520 14427 10523
rect 15654 10520 15660 10532
rect 14415 10492 15660 10520
rect 14415 10489 14427 10492
rect 14369 10483 14427 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 16040 10520 16068 10551
rect 16114 10548 16120 10600
rect 16172 10548 16178 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16356 10560 16865 10588
rect 16356 10548 16362 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 16853 10551 16911 10557
rect 17604 10560 17785 10588
rect 16040 10492 16160 10520
rect 7834 10452 7840 10464
rect 7576 10424 7840 10452
rect 6825 10415 6883 10421
rect 7834 10412 7840 10424
rect 7892 10452 7898 10464
rect 9858 10452 9864 10464
rect 7892 10424 9864 10452
rect 7892 10412 7898 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 11848 10424 13829 10452
rect 11848 10412 11854 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 16132 10452 16160 10492
rect 16482 10480 16488 10532
rect 16540 10520 16546 10532
rect 17604 10520 17632 10560
rect 17773 10557 17785 10560
rect 17819 10588 17831 10591
rect 19536 10588 19564 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21910 10752 21916 10804
rect 21968 10752 21974 10804
rect 21542 10724 21548 10736
rect 21206 10696 21548 10724
rect 21542 10684 21548 10696
rect 21600 10724 21606 10736
rect 21928 10724 21956 10752
rect 22005 10727 22063 10733
rect 22005 10724 22017 10727
rect 21600 10696 22017 10724
rect 21600 10684 21606 10696
rect 22005 10693 22017 10696
rect 22051 10693 22063 10727
rect 22005 10687 22063 10693
rect 17819 10560 19564 10588
rect 17819 10557 17831 10560
rect 17773 10551 17831 10557
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 22646 10588 22652 10600
rect 20027 10560 22652 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 16540 10492 17632 10520
rect 16540 10480 16546 10492
rect 21358 10480 21364 10532
rect 21416 10520 21422 10532
rect 21453 10523 21511 10529
rect 21453 10520 21465 10523
rect 21416 10492 21465 10520
rect 21416 10480 21422 10492
rect 21453 10489 21465 10492
rect 21499 10489 21511 10523
rect 21453 10483 21511 10489
rect 20530 10452 20536 10464
rect 16132 10424 20536 10452
rect 13817 10415 13875 10421
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2590 10248 2596 10260
rect 1995 10220 2596 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3752 10220 3801 10248
rect 3752 10208 3758 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 6288 10220 9076 10248
rect 3602 10140 3608 10192
rect 3660 10180 3666 10192
rect 6288 10180 6316 10220
rect 3660 10152 6316 10180
rect 6365 10183 6423 10189
rect 3660 10140 3666 10152
rect 6365 10149 6377 10183
rect 6411 10180 6423 10183
rect 6549 10183 6607 10189
rect 6549 10180 6561 10183
rect 6411 10152 6561 10180
rect 6411 10149 6423 10152
rect 6365 10143 6423 10149
rect 6549 10149 6561 10152
rect 6595 10180 6607 10183
rect 6730 10180 6736 10192
rect 6595 10152 6736 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 8754 10180 8760 10192
rect 8352 10152 8760 10180
rect 8352 10140 8358 10152
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 9048 10180 9076 10220
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 9674 10248 9680 10260
rect 9232 10220 9680 10248
rect 9232 10180 9260 10220
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10778 10248 10784 10260
rect 10091 10220 10784 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 11698 10248 11704 10260
rect 10888 10220 11704 10248
rect 10888 10180 10916 10220
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 14240 10220 16313 10248
rect 14240 10208 14246 10220
rect 16301 10217 16313 10220
rect 16347 10217 16359 10251
rect 16301 10211 16359 10217
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 17276 10220 18889 10248
rect 17276 10208 17282 10220
rect 18877 10217 18889 10220
rect 18923 10248 18935 10251
rect 19794 10248 19800 10260
rect 18923 10220 19800 10248
rect 18923 10217 18935 10220
rect 18877 10211 18935 10217
rect 19794 10208 19800 10220
rect 19852 10208 19858 10260
rect 21542 10208 21548 10260
rect 21600 10208 21606 10260
rect 9048 10152 9260 10180
rect 9416 10152 10916 10180
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2590 10112 2596 10124
rect 1719 10084 2596 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10081 2927 10115
rect 2869 10075 2927 10081
rect 2130 10004 2136 10056
rect 2188 10004 2194 10056
rect 2884 9976 2912 10075
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4120 10084 4537 10112
rect 4120 10072 4126 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 6825 10115 6883 10121
rect 6825 10112 6837 10115
rect 4856 10084 6837 10112
rect 4856 10072 4862 10084
rect 6825 10081 6837 10084
rect 6871 10112 6883 10115
rect 7834 10112 7840 10124
rect 6871 10084 7840 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 9416 10121 9444 10152
rect 9401 10115 9459 10121
rect 8168 10084 9352 10112
rect 8168 10072 8174 10084
rect 4246 10004 4252 10056
rect 4304 10004 4310 10056
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5684 10016 5825 10044
rect 5684 10004 5690 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 6362 10044 6368 10056
rect 5813 10007 5871 10013
rect 6288 10016 6368 10044
rect 4706 9976 4712 9988
rect 2884 9948 4712 9976
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 6288 9976 6316 10016
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 8846 10044 8852 10056
rect 8234 10016 8852 10044
rect 8846 10004 8852 10016
rect 8904 10044 8910 10056
rect 9122 10044 9128 10056
rect 8904 10016 9128 10044
rect 8904 10004 8910 10016
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9324 10044 9352 10084
rect 9401 10081 9413 10115
rect 9447 10081 9459 10115
rect 9401 10075 9459 10081
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 11974 10112 11980 10124
rect 10735 10084 11980 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 15194 10112 15200 10124
rect 14875 10084 15200 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15194 10072 15200 10084
rect 15252 10112 15258 10124
rect 16206 10112 16212 10124
rect 15252 10084 16212 10112
rect 15252 10072 15258 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 17144 10084 19441 10112
rect 10962 10044 10968 10056
rect 9324 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11238 10004 11244 10056
rect 11296 10004 11302 10056
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14516 10016 14565 10044
rect 14516 10004 14522 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17144 10053 17172 10084
rect 19429 10081 19441 10084
rect 19475 10112 19487 10115
rect 19702 10112 19708 10124
rect 19475 10084 19708 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16908 10016 17141 10044
rect 16908 10004 16914 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 21542 10044 21548 10056
rect 20772 10016 21548 10044
rect 20772 10004 20778 10016
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 5368 9948 6316 9976
rect 1489 9911 1547 9917
rect 1489 9877 1501 9911
rect 1535 9908 1547 9911
rect 2406 9908 2412 9920
rect 1535 9880 2412 9908
rect 1535 9877 1547 9880
rect 1489 9871 1547 9877
rect 2406 9868 2412 9880
rect 2464 9908 2470 9920
rect 5368 9917 5396 9948
rect 7098 9936 7104 9988
rect 7156 9936 7162 9988
rect 10505 9979 10563 9985
rect 10505 9945 10517 9979
rect 10551 9976 10563 9979
rect 11054 9976 11060 9988
rect 10551 9948 11060 9976
rect 10551 9945 10563 9948
rect 10505 9939 10563 9945
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 11517 9979 11575 9985
rect 11517 9945 11529 9979
rect 11563 9976 11575 9979
rect 11790 9976 11796 9988
rect 11563 9948 11796 9976
rect 11563 9945 11575 9948
rect 11517 9939 11575 9945
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 12802 9976 12808 9988
rect 12742 9948 12808 9976
rect 12802 9936 12808 9948
rect 12860 9976 12866 9988
rect 12860 9948 13860 9976
rect 16054 9948 16712 9976
rect 12860 9936 12866 9948
rect 13832 9920 13860 9948
rect 5353 9911 5411 9917
rect 5353 9908 5365 9911
rect 2464 9880 5365 9908
rect 2464 9868 2470 9880
rect 5353 9877 5365 9880
rect 5399 9877 5411 9911
rect 5353 9871 5411 9877
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 8754 9908 8760 9920
rect 8619 9880 8760 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 8904 9880 10425 9908
rect 8904 9868 8910 9880
rect 10413 9877 10425 9880
rect 10459 9877 10471 9911
rect 10413 9871 10471 9877
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 11940 9880 13001 9908
rect 11940 9868 11946 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14185 9911 14243 9917
rect 14185 9908 14197 9911
rect 13872 9880 14197 9908
rect 13872 9868 13878 9880
rect 14185 9877 14197 9880
rect 14231 9908 14243 9911
rect 16132 9908 16160 9948
rect 16684 9917 16712 9948
rect 17034 9936 17040 9988
rect 17092 9976 17098 9988
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 17092 9948 17417 9976
rect 17092 9936 17098 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 18874 9976 18880 9988
rect 18630 9948 18880 9976
rect 17405 9939 17463 9945
rect 14231 9880 16160 9908
rect 16669 9911 16727 9917
rect 14231 9877 14243 9880
rect 14185 9871 14243 9877
rect 16669 9877 16681 9911
rect 16715 9908 16727 9911
rect 16758 9908 16764 9920
rect 16715 9880 16764 9908
rect 16715 9877 16727 9880
rect 16669 9871 16727 9877
rect 16758 9868 16764 9880
rect 16816 9908 16822 9920
rect 16853 9911 16911 9917
rect 16853 9908 16865 9911
rect 16816 9880 16865 9908
rect 16816 9868 16822 9880
rect 16853 9877 16865 9880
rect 16899 9908 16911 9911
rect 18708 9908 18736 9948
rect 18874 9936 18880 9948
rect 18932 9936 18938 9988
rect 19242 9936 19248 9988
rect 19300 9976 19306 9988
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 19300 9948 19717 9976
rect 19300 9936 19306 9948
rect 19705 9945 19717 9948
rect 19751 9945 19763 9979
rect 21634 9976 21640 9988
rect 19705 9939 19763 9945
rect 21008 9948 21640 9976
rect 16899 9880 18736 9908
rect 19720 9908 19748 9939
rect 21008 9908 21036 9948
rect 21634 9936 21640 9948
rect 21692 9936 21698 9988
rect 19720 9880 21036 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 21174 9868 21180 9920
rect 21232 9868 21238 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9704 1639 9707
rect 2130 9704 2136 9716
rect 1627 9676 2136 9704
rect 1627 9673 1639 9676
rect 1581 9667 1639 9673
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 6270 9704 6276 9716
rect 5684 9676 6276 9704
rect 5684 9664 5690 9676
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6457 9707 6515 9713
rect 6457 9673 6469 9707
rect 6503 9704 6515 9707
rect 6730 9704 6736 9716
rect 6503 9676 6736 9704
rect 6503 9673 6515 9676
rect 6457 9667 6515 9673
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 12342 9704 12348 9716
rect 8772 9676 12348 9704
rect 1394 9596 1400 9648
rect 1452 9596 1458 9648
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 1728 9608 3249 9636
rect 1728 9596 1734 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 4062 9636 4068 9648
rect 3237 9599 3295 9605
rect 3804 9608 4068 9636
rect 1026 9528 1032 9580
rect 1084 9568 1090 9580
rect 3804 9577 3832 9608
rect 4062 9596 4068 9608
rect 4120 9636 4126 9648
rect 5721 9639 5779 9645
rect 4120 9608 5304 9636
rect 4120 9596 4126 9608
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 1084 9540 2421 9568
rect 1084 9528 1090 9540
rect 2409 9537 2421 9540
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 5166 9568 5172 9580
rect 3789 9531 3847 9537
rect 4080 9540 5172 9568
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 1903 9472 2145 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2133 9469 2145 9472
rect 2179 9500 2191 9503
rect 4080 9500 4108 9540
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 2179 9472 4108 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 4246 9460 4252 9512
rect 4304 9460 4310 9512
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9469 4583 9503
rect 5276 9500 5304 9608
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 5810 9636 5816 9648
rect 5767 9608 5816 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 8772 9636 8800 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 12860 9676 16160 9704
rect 12860 9664 12866 9676
rect 6840 9608 8800 9636
rect 6840 9577 6868 9608
rect 9122 9596 9128 9648
rect 9180 9596 9186 9648
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 10781 9639 10839 9645
rect 10781 9636 10793 9639
rect 10008 9608 10793 9636
rect 10008 9596 10014 9608
rect 10781 9605 10793 9608
rect 10827 9605 10839 9639
rect 10781 9599 10839 9605
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 13814 9636 13820 9648
rect 13202 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9636 13878 9648
rect 13909 9639 13967 9645
rect 13909 9636 13921 9639
rect 13872 9608 13921 9636
rect 13872 9596 13878 9608
rect 13909 9605 13921 9608
rect 13955 9605 13967 9639
rect 13909 9599 13967 9605
rect 14185 9639 14243 9645
rect 14185 9605 14197 9639
rect 14231 9636 14243 9639
rect 14366 9636 14372 9648
rect 14231 9608 14372 9636
rect 14231 9605 14243 9608
rect 14185 9599 14243 9605
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 16132 9636 16160 9676
rect 16206 9664 16212 9716
rect 16264 9664 16270 9716
rect 24486 9704 24492 9716
rect 16316 9676 24492 9704
rect 16316 9636 16344 9676
rect 24486 9664 24492 9676
rect 24544 9664 24550 9716
rect 16132 9608 16344 9636
rect 16758 9596 16764 9648
rect 16816 9596 16822 9648
rect 17129 9639 17187 9645
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 17218 9636 17224 9648
rect 17175 9608 17224 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 18874 9636 18880 9648
rect 18354 9608 18880 9636
rect 18874 9596 18880 9608
rect 18932 9596 18938 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 24578 9636 24584 9648
rect 19567 9608 24584 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 24578 9596 24584 9608
rect 24636 9596 24642 9648
rect 28629 9639 28687 9645
rect 28629 9605 28641 9639
rect 28675 9636 28687 9639
rect 31294 9636 31300 9648
rect 28675 9608 31300 9636
rect 28675 9605 28687 9608
rect 28629 9599 28687 9605
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 7374 9568 7380 9580
rect 6825 9531 6883 9537
rect 6932 9540 7380 9568
rect 6932 9500 6960 9540
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9732 9540 10701 9568
rect 9732 9528 9738 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 16776 9568 16804 9596
rect 15870 9540 16804 9568
rect 19429 9571 19487 9577
rect 10689 9531 10747 9537
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 20622 9568 20628 9580
rect 20211 9540 20628 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 5276 9472 6960 9500
rect 7101 9503 7159 9509
rect 4525 9463 4583 9469
rect 7101 9469 7113 9503
rect 7147 9500 7159 9503
rect 7147 9472 7512 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 3970 9432 3976 9444
rect 3651 9404 3976 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 3970 9392 3976 9404
rect 4028 9392 4034 9444
rect 4540 9432 4568 9463
rect 7374 9432 7380 9444
rect 4540 9404 7380 9432
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 7484 9432 7512 9472
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7892 9472 8125 9500
rect 7892 9460 7898 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8478 9500 8484 9512
rect 8435 9472 8484 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 8812 9472 10885 9500
rect 8812 9460 8818 9472
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11296 9472 11713 9500
rect 11296 9460 11302 9472
rect 11701 9469 11713 9472
rect 11747 9500 11759 9503
rect 14458 9500 14464 9512
rect 11747 9472 14464 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 16758 9500 16764 9512
rect 14792 9472 16764 9500
rect 14792 9460 14798 9472
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 19444 9500 19472 9531
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 23750 9528 23756 9580
rect 23808 9568 23814 9580
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 23808 9540 27537 9568
rect 23808 9528 23814 9540
rect 27525 9537 27537 9540
rect 27571 9568 27583 9571
rect 28166 9568 28172 9580
rect 27571 9540 28172 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 28166 9528 28172 9540
rect 28224 9528 28230 9580
rect 16960 9472 19472 9500
rect 19705 9503 19763 9509
rect 7926 9432 7932 9444
rect 7484 9404 7932 9432
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 13412 9404 13461 9432
rect 13412 9392 13418 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 14274 9432 14280 9444
rect 13449 9395 13507 9401
rect 13556 9404 14280 9432
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 3752 9336 5365 9364
rect 3752 9324 3758 9336
rect 5353 9333 5365 9336
rect 5399 9364 5411 9367
rect 6270 9364 6276 9376
rect 5399 9336 6276 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 8754 9364 8760 9376
rect 7156 9336 8760 9364
rect 7156 9324 7162 9336
rect 8754 9324 8760 9336
rect 8812 9364 8818 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 8812 9336 9873 9364
rect 8812 9324 8818 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9364 10379 9367
rect 13556 9364 13584 9404
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 16960 9432 16988 9472
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 21174 9500 21180 9512
rect 19751 9472 21180 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 23440 9472 27997 9500
rect 23440 9460 23446 9472
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 28644 9500 28672 9599
rect 31294 9596 31300 9608
rect 31352 9596 31358 9648
rect 27985 9463 28043 9469
rect 28184 9472 28672 9500
rect 15764 9404 16988 9432
rect 10367 9336 13584 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 13998 9324 14004 9376
rect 14056 9364 14062 9376
rect 15764 9364 15792 9404
rect 19058 9392 19064 9444
rect 19116 9392 19122 9444
rect 14056 9336 15792 9364
rect 14056 9324 14062 9336
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 16172 9336 18613 9364
rect 16172 9324 16178 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18601 9327 18659 9333
rect 27801 9367 27859 9373
rect 27801 9333 27813 9367
rect 27847 9364 27859 9367
rect 28184 9364 28212 9472
rect 27847 9336 28212 9364
rect 27847 9333 27859 9336
rect 27801 9327 27859 9333
rect 28350 9324 28356 9376
rect 28408 9364 28414 9376
rect 28445 9367 28503 9373
rect 28445 9364 28457 9367
rect 28408 9336 28457 9364
rect 28408 9324 28414 9336
rect 28445 9333 28457 9336
rect 28491 9364 28503 9367
rect 31570 9364 31576 9376
rect 28491 9336 31576 9364
rect 28491 9333 28503 9336
rect 28445 9327 28503 9333
rect 31570 9324 31576 9336
rect 31628 9324 31634 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3513 9163 3571 9169
rect 3513 9160 3525 9163
rect 3476 9132 3525 9160
rect 3476 9120 3482 9132
rect 3513 9129 3525 9132
rect 3559 9129 3571 9163
rect 3513 9123 3571 9129
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 5261 9163 5319 9169
rect 5261 9160 5273 9163
rect 4304 9132 5273 9160
rect 4304 9120 4310 9132
rect 5261 9129 5273 9132
rect 5307 9129 5319 9163
rect 5261 9123 5319 9129
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 9674 9160 9680 9172
rect 7883 9132 9680 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10134 9120 10140 9172
rect 10192 9120 10198 9172
rect 11514 9160 11520 9172
rect 10244 9132 11520 9160
rect 4522 9052 4528 9104
rect 4580 9092 4586 9104
rect 7926 9092 7932 9104
rect 4580 9064 4660 9092
rect 4580 9052 4586 9064
rect 1210 8984 1216 9036
rect 1268 9024 1274 9036
rect 2501 9027 2559 9033
rect 2501 9024 2513 9027
rect 1268 8996 2513 9024
rect 1268 8984 1274 8996
rect 2501 8993 2513 8996
rect 2547 8993 2559 9027
rect 2501 8987 2559 8993
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 9024 3479 9027
rect 3786 9024 3792 9036
rect 3467 8996 3792 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 4632 9033 4660 9064
rect 4724 9064 7932 9092
rect 4617 9027 4675 9033
rect 4617 8993 4629 9027
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 1854 8956 1860 8968
rect 1811 8928 1860 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2314 8956 2320 8968
rect 2271 8928 2320 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2240 8820 2268 8919
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 4724 8956 4752 9064
rect 7926 9052 7932 9064
rect 7984 9092 7990 9104
rect 7984 9064 8340 9092
rect 7984 9052 7990 9064
rect 6178 8984 6184 9036
rect 6236 8984 6242 9036
rect 4580 8928 4752 8956
rect 4580 8916 4586 8928
rect 5442 8916 5448 8968
rect 5500 8916 5506 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7558 8956 7564 8968
rect 7423 8928 7564 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 5920 8888 5948 8919
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8312 8956 8340 9064
rect 8478 9052 8484 9104
rect 8536 9092 8542 9104
rect 9950 9092 9956 9104
rect 8536 9064 9956 9092
rect 8536 9052 8542 9064
rect 9950 9052 9956 9064
rect 10008 9052 10014 9104
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 9024 8447 9027
rect 8754 9024 8760 9036
rect 8435 8996 8760 9024
rect 8435 8993 8447 8996
rect 8389 8987 8447 8993
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 9024 9459 9027
rect 9766 9024 9772 9036
rect 9447 8996 9772 9024
rect 9447 8993 9459 8996
rect 9401 8987 9459 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 10244 8956 10272 9132
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 14182 9160 14188 9172
rect 12406 9132 14188 9160
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 9024 10839 9027
rect 12406 9024 12434 9132
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 15930 9160 15936 9172
rect 14323 9132 15936 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16482 9160 16488 9172
rect 16132 9132 16488 9160
rect 15378 9052 15384 9104
rect 15436 9052 15442 9104
rect 16132 9092 16160 9132
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16758 9120 16764 9172
rect 16816 9160 16822 9172
rect 17402 9160 17408 9172
rect 16816 9132 17408 9160
rect 16816 9120 16822 9132
rect 17402 9120 17408 9132
rect 17460 9160 17466 9172
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 17460 9132 17785 9160
rect 17460 9120 17466 9132
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 17773 9123 17831 9129
rect 18141 9163 18199 9169
rect 18141 9129 18153 9163
rect 18187 9160 18199 9163
rect 18785 9163 18843 9169
rect 18785 9160 18797 9163
rect 18187 9132 18797 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 18785 9129 18797 9132
rect 18831 9160 18843 9163
rect 18874 9160 18880 9172
rect 18831 9132 18880 9160
rect 18831 9129 18843 9132
rect 18785 9123 18843 9129
rect 15948 9064 16160 9092
rect 10827 8996 12434 9024
rect 10827 8993 10839 8996
rect 10781 8987 10839 8993
rect 14366 8984 14372 9036
rect 14424 9024 14430 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14424 8996 14749 9024
rect 14424 8984 14430 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 9024 14979 9027
rect 15948 9024 15976 9064
rect 14967 8996 15976 9024
rect 16025 9027 16083 9033
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16850 9024 16856 9036
rect 16071 8996 16856 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 8312 8928 10272 8956
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10376 8928 11345 8956
rect 10376 8916 10382 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 18156 8956 18184 9123
rect 18874 9120 18880 9132
rect 18932 9160 18938 9172
rect 18969 9163 19027 9169
rect 18969 9160 18981 9163
rect 18932 9132 18981 9160
rect 18932 9120 18938 9132
rect 18969 9129 18981 9132
rect 19015 9160 19027 9163
rect 19426 9160 19432 9172
rect 19015 9132 19432 9160
rect 19015 9129 19027 9132
rect 18969 9123 19027 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 11655 8928 16068 8956
rect 17434 8928 18184 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 9122 8888 9128 8900
rect 5920 8860 9128 8888
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 10505 8891 10563 8897
rect 10505 8857 10517 8891
rect 10551 8888 10563 8891
rect 10962 8888 10968 8900
rect 10551 8860 10968 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 13541 8891 13599 8897
rect 13541 8857 13553 8891
rect 13587 8888 13599 8891
rect 14645 8891 14703 8897
rect 14645 8888 14657 8891
rect 13587 8860 14657 8888
rect 13587 8857 13599 8860
rect 13541 8851 13599 8857
rect 14645 8857 14657 8860
rect 14691 8857 14703 8891
rect 14645 8851 14703 8857
rect 1627 8792 2268 8820
rect 3973 8823 4031 8829
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 7282 8820 7288 8832
rect 4019 8792 7288 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 9033 8823 9091 8829
rect 9033 8789 9045 8823
rect 9079 8820 9091 8823
rect 9214 8820 9220 8832
rect 9079 8792 9220 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 9732 8792 10609 8820
rect 9732 8780 9738 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10597 8783 10655 8789
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 12584 8792 12633 8820
rect 12584 8780 12590 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 12621 8783 12679 8789
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 15562 8820 15568 8832
rect 13964 8792 15568 8820
rect 13964 8780 13970 8792
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 16040 8820 16068 8928
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 16264 8860 16313 8888
rect 16264 8848 16270 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 16301 8851 16359 8857
rect 17218 8820 17224 8832
rect 16040 8792 17224 8820
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 566 8576 572 8628
rect 624 8616 630 8628
rect 7285 8619 7343 8625
rect 624 8588 6040 8616
rect 624 8576 630 8588
rect 750 8508 756 8560
rect 808 8548 814 8560
rect 808 8520 4660 8548
rect 808 8508 814 8520
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 2774 8480 2780 8492
rect 1627 8452 2780 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 2866 8440 2872 8492
rect 2924 8440 2930 8492
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3510 8480 3516 8492
rect 3191 8452 3516 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4522 8480 4528 8492
rect 4387 8452 4528 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8381 1915 8415
rect 1857 8375 1915 8381
rect 1872 8344 1900 8375
rect 3694 8344 3700 8356
rect 1872 8316 3700 8344
rect 3694 8304 3700 8316
rect 3752 8304 3758 8356
rect 4632 8353 4660 8520
rect 5074 8508 5080 8560
rect 5132 8508 5138 8560
rect 5350 8508 5356 8560
rect 5408 8508 5414 8560
rect 6012 8489 6040 8588
rect 7285 8585 7297 8619
rect 7331 8616 7343 8619
rect 8570 8616 8576 8628
rect 7331 8588 8576 8616
rect 7331 8585 7343 8588
rect 7285 8579 7343 8585
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 12434 8616 12440 8628
rect 10183 8588 12440 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12526 8576 12532 8628
rect 12584 8576 12590 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 14918 8616 14924 8628
rect 14323 8588 14924 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16298 8616 16304 8628
rect 15979 8588 16304 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 17218 8576 17224 8628
rect 17276 8616 17282 8628
rect 32490 8616 32496 8628
rect 17276 8588 32496 8616
rect 17276 8576 17282 8588
rect 32490 8576 32496 8588
rect 32548 8576 32554 8628
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 11241 8551 11299 8557
rect 6972 8520 8708 8548
rect 6972 8508 6978 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 7742 8480 7748 8492
rect 7239 8452 7748 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 4816 8412 4844 8443
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 7926 8440 7932 8492
rect 7984 8440 7990 8492
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8570 8480 8576 8492
rect 8168 8452 8576 8480
rect 8168 8440 8174 8452
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8680 8489 8708 8520
rect 11241 8517 11253 8551
rect 11287 8548 11299 8551
rect 11422 8548 11428 8560
rect 11287 8520 11428 8548
rect 11287 8517 11299 8520
rect 11241 8511 11299 8517
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 14734 8548 14740 8560
rect 11532 8520 14740 8548
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 5350 8412 5356 8424
rect 4816 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8412 5414 8424
rect 5408 8384 5948 8412
rect 5408 8372 5414 8384
rect 4617 8347 4675 8353
rect 4617 8313 4629 8347
rect 4663 8313 4675 8347
rect 4617 8307 4675 8313
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5316 8316 5825 8344
rect 5316 8304 5322 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5920 8344 5948 8384
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7064 8384 8033 8412
rect 7064 8372 7070 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8412 8447 8415
rect 8435 8384 8616 8412
rect 8435 8381 8447 8384
rect 8389 8375 8447 8381
rect 8478 8344 8484 8356
rect 5920 8316 8484 8344
rect 5813 8307 5871 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8588 8344 8616 8384
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9030 8412 9036 8424
rect 8812 8384 9036 8412
rect 8812 8372 8818 8384
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 9677 8415 9735 8421
rect 9677 8412 9689 8415
rect 9272 8384 9689 8412
rect 9272 8372 9278 8384
rect 9677 8381 9689 8384
rect 9723 8412 9735 8415
rect 10318 8412 10324 8424
rect 9723 8384 10324 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11532 8412 11560 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 15378 8508 15384 8560
rect 15436 8548 15442 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 15436 8520 16037 8548
rect 15436 8508 15442 8520
rect 16025 8517 16037 8520
rect 16071 8517 16083 8551
rect 16025 8511 16083 8517
rect 16114 8508 16120 8560
rect 16172 8548 16178 8560
rect 17310 8548 17316 8560
rect 16172 8520 17316 8548
rect 16172 8508 16178 8520
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 11606 8440 11612 8492
rect 11664 8440 11670 8492
rect 12710 8480 12716 8492
rect 11716 8452 12716 8480
rect 10827 8384 11560 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 9858 8344 9864 8356
rect 8588 8316 9864 8344
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 10336 8344 10364 8372
rect 11716 8344 11744 8452
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13679 8452 14657 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 17126 8480 17132 8492
rect 14645 8443 14703 8449
rect 14936 8452 17132 8480
rect 12618 8372 12624 8424
rect 12676 8372 12682 8424
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8412 12863 8415
rect 12851 8384 14596 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 10336 8316 11744 8344
rect 12161 8347 12219 8353
rect 12161 8313 12173 8347
rect 12207 8344 12219 8347
rect 13906 8344 13912 8356
rect 12207 8316 13912 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 13906 8304 13912 8316
rect 13964 8304 13970 8356
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 3786 8276 3792 8288
rect 3568 8248 3792 8276
rect 3568 8236 3574 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 5960 8248 6377 8276
rect 5960 8236 5966 8248
rect 6365 8245 6377 8248
rect 6411 8276 6423 8279
rect 6454 8276 6460 8288
rect 6411 8248 6460 8276
rect 6411 8245 6423 8248
rect 6365 8239 6423 8245
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 6733 8279 6791 8285
rect 6733 8245 6745 8279
rect 6779 8276 6791 8279
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 6779 8248 7757 8276
rect 6779 8245 6791 8248
rect 6733 8239 6791 8245
rect 7745 8245 7757 8248
rect 7791 8276 7803 8279
rect 9214 8276 9220 8288
rect 7791 8248 9220 8276
rect 7791 8245 7803 8248
rect 7745 8239 7803 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 14568 8276 14596 8384
rect 14734 8372 14740 8424
rect 14792 8372 14798 8424
rect 14936 8421 14964 8452
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8381 14979 8415
rect 16114 8412 16120 8424
rect 14921 8375 14979 8381
rect 15028 8384 16120 8412
rect 15028 8276 15056 8384
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 20346 8412 20352 8424
rect 16255 8384 20352 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 15565 8347 15623 8353
rect 15565 8313 15577 8347
rect 15611 8344 15623 8347
rect 20438 8344 20444 8356
rect 15611 8316 20444 8344
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 14568 8248 15056 8276
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3694 8072 3700 8084
rect 3467 8044 3700 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 5166 8032 5172 8084
rect 5224 8032 5230 8084
rect 5350 8032 5356 8084
rect 5408 8032 5414 8084
rect 6362 8032 6368 8084
rect 6420 8032 6426 8084
rect 6546 8032 6552 8084
rect 6604 8032 6610 8084
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 7742 8032 7748 8084
rect 7800 8032 7806 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 8352 8044 9597 8072
rect 8352 8032 8358 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 12066 8072 12072 8084
rect 9824 8044 12072 8072
rect 9824 8032 9830 8044
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12434 8032 12440 8084
rect 12492 8032 12498 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13998 8072 14004 8084
rect 13035 8044 14004 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 19242 8072 19248 8084
rect 14240 8044 19248 8072
rect 14240 8032 14246 8044
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 842 7964 848 8016
rect 900 8004 906 8016
rect 3513 8007 3571 8013
rect 3513 8004 3525 8007
rect 900 7976 3525 8004
rect 900 7964 906 7976
rect 3513 7973 3525 7976
rect 3559 7973 3571 8007
rect 3513 7967 3571 7973
rect 5718 7964 5724 8016
rect 5776 7964 5782 8016
rect 6638 7964 6644 8016
rect 6696 8004 6702 8016
rect 6696 7976 9628 8004
rect 6696 7964 6702 7976
rect 1486 7896 1492 7948
rect 1544 7936 1550 7948
rect 1581 7939 1639 7945
rect 1581 7936 1593 7939
rect 1544 7908 1593 7936
rect 1544 7896 1550 7908
rect 1581 7905 1593 7908
rect 1627 7936 1639 7939
rect 3786 7936 3792 7948
rect 1627 7908 3792 7936
rect 1627 7905 1639 7908
rect 1581 7899 1639 7905
rect 3786 7896 3792 7908
rect 3844 7896 3850 7948
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 7374 7936 7380 7948
rect 7147 7908 7380 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7374 7896 7380 7908
rect 7432 7936 7438 7948
rect 8110 7936 8116 7948
rect 7432 7908 8116 7936
rect 7432 7896 7438 7908
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 9214 7936 9220 7948
rect 8803 7908 9220 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9600 7936 9628 7976
rect 9876 7976 13584 8004
rect 9876 7936 9904 7976
rect 9600 7908 9904 7936
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10008 7908 10241 7936
rect 10008 7896 10014 7908
rect 10229 7905 10241 7908
rect 10275 7936 10287 7939
rect 10870 7936 10876 7948
rect 10275 7908 10876 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 12434 7936 12440 7948
rect 11287 7908 12440 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 2498 7868 2504 7880
rect 1903 7840 2504 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3602 7868 3608 7880
rect 3099 7840 3608 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 4172 7800 4200 7831
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4304 7840 4813 7868
rect 4304 7828 4310 7840
rect 4801 7837 4813 7840
rect 4847 7868 4859 7871
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 4847 7840 5457 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 5445 7837 5457 7840
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7524 7840 7849 7868
rect 7524 7828 7530 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 10045 7871 10103 7877
rect 7837 7831 7895 7837
rect 8036 7840 9996 7868
rect 5718 7800 5724 7812
rect 992 7772 3648 7800
rect 4172 7772 5724 7800
rect 992 7760 998 7772
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 2958 7732 2964 7744
rect 2915 7704 2964 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3620 7732 3648 7772
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 8036 7800 8064 7840
rect 9968 7809 9996 7840
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 11146 7868 11152 7880
rect 10091 7840 11152 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11514 7828 11520 7880
rect 11572 7828 11578 7880
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 13556 7868 13584 7976
rect 15194 7964 15200 8016
rect 15252 7964 15258 8016
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 14182 7936 14188 7948
rect 13679 7908 14188 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 14829 7939 14887 7945
rect 14829 7905 14841 7939
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 14844 7868 14872 7899
rect 13556 7840 14872 7868
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15068 7840 15884 7868
rect 15068 7828 15074 7840
rect 6880 7772 8064 7800
rect 9953 7803 10011 7809
rect 6880 7760 6886 7772
rect 9953 7769 9965 7803
rect 9999 7769 10011 7803
rect 9953 7763 10011 7769
rect 13357 7803 13415 7809
rect 13357 7769 13369 7803
rect 13403 7800 13415 7803
rect 13538 7800 13544 7812
rect 13403 7772 13544 7800
rect 13403 7769 13415 7772
rect 13357 7763 13415 7769
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3620 7704 3985 7732
rect 3973 7701 3985 7704
rect 4019 7701 4031 7735
rect 3973 7695 4031 7701
rect 4617 7735 4675 7741
rect 4617 7701 4629 7735
rect 4663 7732 4675 7735
rect 9766 7732 9772 7744
rect 4663 7704 9772 7732
rect 4663 7701 4675 7704
rect 4617 7695 4675 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 9968 7732 9996 7763
rect 13538 7760 13544 7772
rect 13596 7760 13602 7812
rect 14734 7732 14740 7744
rect 9968 7704 14740 7732
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 15856 7741 15884 7840
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 22830 7732 22836 7744
rect 15887 7704 22836 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 22830 7692 22836 7704
rect 22888 7732 22894 7744
rect 23382 7732 23388 7744
rect 22888 7704 23388 7732
rect 22888 7692 22894 7704
rect 23382 7692 23388 7704
rect 23440 7692 23446 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3326 7528 3332 7540
rect 2915 7500 3332 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 3602 7488 3608 7540
rect 3660 7488 3666 7540
rect 4430 7528 4436 7540
rect 3712 7500 4436 7528
rect 1302 7420 1308 7472
rect 1360 7460 1366 7472
rect 1360 7432 2774 7460
rect 1360 7420 1366 7432
rect 1578 7352 1584 7404
rect 1636 7352 1642 7404
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2222 7392 2228 7404
rect 1903 7364 2228 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2746 7392 2774 7432
rect 2958 7420 2964 7472
rect 3016 7460 3022 7472
rect 3712 7460 3740 7500
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 7650 7528 7656 7540
rect 4663 7500 7656 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11885 7531 11943 7537
rect 11885 7528 11897 7531
rect 11020 7500 11897 7528
rect 11020 7488 11026 7500
rect 11885 7497 11897 7500
rect 11931 7497 11943 7531
rect 11885 7491 11943 7497
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7528 13507 7531
rect 13538 7528 13544 7540
rect 13495 7500 13544 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 27614 7528 27620 7540
rect 23992 7500 27620 7528
rect 23992 7488 23998 7500
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 3016 7432 3740 7460
rect 4172 7432 5396 7460
rect 3016 7420 3022 7432
rect 3053 7395 3111 7401
rect 3053 7392 3065 7395
rect 2746 7364 3065 7392
rect 3053 7361 3065 7364
rect 3099 7392 3111 7395
rect 3326 7392 3332 7404
rect 3099 7364 3332 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4172 7401 4200 7432
rect 5368 7404 5396 7432
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 5592 7432 10824 7460
rect 5592 7420 5598 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 4304 7364 4813 7392
rect 4304 7352 4310 7364
rect 4801 7361 4813 7364
rect 4847 7392 4859 7395
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4847 7364 5089 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5350 7352 5356 7404
rect 5408 7352 5414 7404
rect 8938 7352 8944 7404
rect 8996 7392 9002 7404
rect 10796 7401 10824 7432
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 15010 7460 15016 7472
rect 12124 7432 15016 7460
rect 12124 7420 12130 7432
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 24302 7460 24308 7472
rect 23690 7432 24308 7460
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 9309 7395 9367 7401
rect 9309 7392 9321 7395
rect 8996 7364 9321 7392
rect 8996 7352 9002 7364
rect 9309 7361 9321 7364
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 11330 7352 11336 7404
rect 11388 7392 11394 7404
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 11388 7364 12725 7392
rect 11388 7352 11394 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 11514 7324 11520 7336
rect 6512 7296 11520 7324
rect 6512 7284 6518 7296
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 22462 7284 22468 7336
rect 22520 7284 22526 7336
rect 2866 7216 2872 7268
rect 2924 7256 2930 7268
rect 3329 7259 3387 7265
rect 3329 7256 3341 7259
rect 2924 7228 3341 7256
rect 2924 7216 2930 7228
rect 3329 7225 3341 7228
rect 3375 7225 3387 7259
rect 3329 7219 3387 7225
rect 3970 7216 3976 7268
rect 4028 7216 4034 7268
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 12434 7188 12440 7200
rect 10643 7160 12440 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 12529 7191 12587 7197
rect 12529 7157 12541 7191
rect 12575 7188 12587 7191
rect 13998 7188 14004 7200
rect 12575 7160 14004 7188
rect 12575 7157 12587 7160
rect 12529 7151 12587 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 17494 7188 17500 7200
rect 14139 7160 17500 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 1489 6987 1547 6993
rect 1489 6953 1501 6987
rect 1535 6984 1547 6987
rect 1578 6984 1584 6996
rect 1535 6956 1584 6984
rect 1535 6953 1547 6956
rect 1489 6947 1547 6953
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 2593 6987 2651 6993
rect 2593 6953 2605 6987
rect 2639 6984 2651 6987
rect 2682 6984 2688 6996
rect 2639 6956 2688 6984
rect 2639 6953 2651 6956
rect 2593 6947 2651 6953
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 3237 6987 3295 6993
rect 3237 6953 3249 6987
rect 3283 6984 3295 6987
rect 5166 6984 5172 6996
rect 3283 6956 5172 6984
rect 3283 6953 3295 6956
rect 3237 6947 3295 6953
rect 5166 6944 5172 6956
rect 5224 6944 5230 6996
rect 23201 6987 23259 6993
rect 23201 6953 23213 6987
rect 23247 6984 23259 6987
rect 23934 6984 23940 6996
rect 23247 6956 23940 6984
rect 23247 6953 23259 6956
rect 23201 6947 23259 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 3878 6916 3884 6928
rect 3252 6888 3884 6916
rect 750 6808 756 6860
rect 808 6848 814 6860
rect 1581 6851 1639 6857
rect 1581 6848 1593 6851
rect 808 6820 1593 6848
rect 808 6808 814 6820
rect 1581 6817 1593 6820
rect 1627 6817 1639 6851
rect 3252 6848 3280 6888
rect 3878 6876 3884 6888
rect 3936 6876 3942 6928
rect 3973 6919 4031 6925
rect 3973 6885 3985 6919
rect 4019 6916 4031 6919
rect 4019 6888 4936 6916
rect 4019 6885 4031 6888
rect 3973 6879 4031 6885
rect 1581 6811 1639 6817
rect 2148 6820 3280 6848
rect 3344 6820 3740 6848
rect 2148 6789 2176 6820
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 3142 6780 3148 6792
rect 2823 6752 3148 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 3142 6740 3148 6752
rect 3200 6780 3206 6792
rect 3344 6780 3372 6820
rect 3200 6752 3372 6780
rect 3421 6783 3479 6789
rect 3200 6740 3206 6752
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3712 6780 3740 6820
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 3844 6820 4813 6848
rect 3844 6808 3850 6820
rect 4801 6817 4813 6820
rect 4847 6817 4859 6851
rect 4908 6848 4936 6888
rect 23750 6876 23756 6928
rect 23808 6876 23814 6928
rect 8846 6848 8852 6860
rect 4908 6820 8852 6848
rect 4801 6811 4859 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10560 6820 10609 6848
rect 10560 6808 10566 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 3970 6780 3976 6792
rect 3712 6752 3976 6780
rect 3421 6743 3479 6749
rect 3436 6712 3464 6743
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 4120 6752 4169 6780
rect 4120 6740 4126 6752
rect 4157 6749 4169 6752
rect 4203 6780 4215 6783
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 4203 6752 4445 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 21726 6740 21732 6792
rect 21784 6780 21790 6792
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 21784 6752 22937 6780
rect 21784 6740 21790 6752
rect 22925 6749 22937 6752
rect 22971 6780 22983 6783
rect 23768 6780 23796 6876
rect 22971 6752 23796 6780
rect 22971 6749 22983 6752
rect 22925 6743 22983 6749
rect 4338 6712 4344 6724
rect 3436 6684 4344 6712
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 3510 6644 3516 6656
rect 1995 6616 3516 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4028 6616 4629 6644
rect 4028 6604 4034 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 23382 6604 23388 6656
rect 23440 6604 23446 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 3326 6400 3332 6452
rect 3384 6440 3390 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 3384 6412 3985 6440
rect 3384 6400 3390 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 3973 6403 4031 6409
rect 22830 6400 22836 6452
rect 22888 6400 22894 6452
rect 12158 6372 12164 6384
rect 1872 6344 12164 6372
rect 1872 6313 1900 6344
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2832 6276 3065 6304
rect 2832 6264 2838 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 4157 6307 4215 6313
rect 4157 6304 4169 6307
rect 3752 6276 4169 6304
rect 3752 6264 3758 6276
rect 4157 6273 4169 6276
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 22424 6307 22482 6313
rect 22424 6273 22436 6307
rect 22470 6304 22482 6307
rect 22848 6304 22876 6400
rect 22470 6276 22876 6304
rect 22470 6273 22482 6276
rect 22424 6267 22482 6273
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 1360 6208 1593 6236
rect 1360 6196 1366 6208
rect 1581 6205 1593 6208
rect 1627 6236 1639 6239
rect 2866 6236 2872 6248
rect 1627 6208 2872 6236
rect 1627 6205 1639 6208
rect 1581 6199 1639 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 22511 6239 22569 6245
rect 22511 6205 22523 6239
rect 22557 6236 22569 6239
rect 24854 6236 24860 6248
rect 22557 6208 24860 6236
rect 22557 6205 22569 6208
rect 22511 6199 22569 6205
rect 24854 6196 24860 6208
rect 24912 6196 24918 6248
rect 3513 6171 3571 6177
rect 3513 6137 3525 6171
rect 3559 6168 3571 6171
rect 6086 6168 6092 6180
rect 3559 6140 6092 6168
rect 3559 6137 3571 6140
rect 3513 6131 3571 6137
rect 6086 6128 6092 6140
rect 6144 6128 6150 6180
rect 19334 6128 19340 6180
rect 19392 6168 19398 6180
rect 38746 6168 38752 6180
rect 19392 6140 38752 6168
rect 19392 6128 19398 6140
rect 38746 6128 38752 6140
rect 38804 6128 38810 6180
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6100 2927 6103
rect 4062 6100 4068 6112
rect 2915 6072 4068 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 3329 5899 3387 5905
rect 3329 5896 3341 5899
rect 2832 5868 3341 5896
rect 2832 5856 2838 5868
rect 3329 5865 3341 5868
rect 3375 5865 3387 5899
rect 3329 5859 3387 5865
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 3878 5896 3884 5908
rect 3651 5868 3884 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 18923 5868 21005 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 20993 5865 21005 5868
rect 21039 5896 21051 5899
rect 22462 5896 22468 5908
rect 21039 5868 22468 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 2869 5831 2927 5837
rect 2869 5797 2881 5831
rect 2915 5828 2927 5831
rect 9306 5828 9312 5840
rect 2915 5800 9312 5828
rect 2915 5797 2927 5800
rect 2869 5791 2927 5797
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 9582 5788 9588 5840
rect 9640 5828 9646 5840
rect 12618 5828 12624 5840
rect 9640 5800 12624 5828
rect 9640 5788 9646 5800
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 19337 5831 19395 5837
rect 19337 5797 19349 5831
rect 19383 5828 19395 5831
rect 19426 5828 19432 5840
rect 19383 5800 19432 5828
rect 19383 5797 19395 5800
rect 19337 5791 19395 5797
rect 1210 5720 1216 5772
rect 1268 5760 1274 5772
rect 1857 5763 1915 5769
rect 1268 5732 1808 5760
rect 1268 5720 1274 5732
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1780 5692 1808 5732
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 3602 5760 3608 5772
rect 1903 5732 3608 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 3602 5720 3608 5732
rect 3660 5720 3666 5772
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 14056 5732 15577 5760
rect 14056 5720 14062 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 16908 5732 17141 5760
rect 16908 5720 16914 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 2774 5692 2780 5704
rect 1780 5664 2780 5692
rect 1581 5655 1639 5661
rect 1596 5624 1624 5655
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2832 5664 3065 5692
rect 2832 5652 2838 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 12676 5664 15761 5692
rect 12676 5652 12682 5664
rect 15749 5661 15761 5664
rect 15795 5692 15807 5695
rect 19352 5692 19380 5791
rect 19426 5788 19432 5800
rect 19484 5788 19490 5840
rect 21726 5788 21732 5840
rect 21784 5788 21790 5840
rect 15795 5664 17172 5692
rect 18538 5664 19380 5692
rect 15795 5661 15807 5664
rect 15749 5655 15807 5661
rect 2958 5624 2964 5636
rect 1596 5596 2964 5624
rect 2958 5584 2964 5596
rect 3016 5584 3022 5636
rect 16209 5559 16267 5565
rect 16209 5525 16221 5559
rect 16255 5556 16267 5559
rect 17034 5556 17040 5568
rect 16255 5528 17040 5556
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 17144 5556 17172 5664
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20312 5664 20913 5692
rect 20312 5652 20318 5664
rect 20901 5661 20913 5664
rect 20947 5692 20959 5695
rect 21744 5692 21772 5788
rect 27065 5763 27123 5769
rect 27065 5729 27077 5763
rect 27111 5760 27123 5763
rect 30282 5760 30288 5772
rect 27111 5732 30288 5760
rect 27111 5729 27123 5732
rect 27065 5723 27123 5729
rect 30282 5720 30288 5732
rect 30340 5720 30346 5772
rect 20947 5664 21772 5692
rect 20947 5661 20959 5664
rect 20901 5655 20959 5661
rect 17402 5584 17408 5636
rect 17460 5584 17466 5636
rect 22186 5624 22192 5636
rect 18708 5596 22192 5624
rect 18708 5556 18736 5596
rect 22186 5584 22192 5596
rect 22244 5624 22250 5636
rect 23382 5624 23388 5636
rect 22244 5596 23388 5624
rect 22244 5584 22250 5596
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 24765 5627 24823 5633
rect 24765 5593 24777 5627
rect 24811 5593 24823 5627
rect 24765 5587 24823 5593
rect 17144 5528 18736 5556
rect 21358 5516 21364 5568
rect 21416 5516 21422 5568
rect 24780 5556 24808 5587
rect 24854 5584 24860 5636
rect 24912 5584 24918 5636
rect 25774 5584 25780 5636
rect 25832 5584 25838 5636
rect 27154 5584 27160 5636
rect 27212 5584 27218 5636
rect 28077 5627 28135 5633
rect 28077 5593 28089 5627
rect 28123 5624 28135 5627
rect 35710 5624 35716 5636
rect 28123 5596 35716 5624
rect 28123 5593 28135 5596
rect 28077 5587 28135 5593
rect 35710 5584 35716 5596
rect 35768 5584 35774 5636
rect 25498 5556 25504 5568
rect 24780 5528 25504 5556
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 2774 5312 2780 5364
rect 2832 5312 2838 5364
rect 2866 5312 2872 5364
rect 2924 5312 2930 5364
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 3016 5324 3065 5352
rect 3016 5312 3022 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 22879 5355 22937 5361
rect 22879 5321 22891 5355
rect 22925 5352 22937 5355
rect 27154 5352 27160 5364
rect 22925 5324 27160 5352
rect 22925 5321 22937 5324
rect 22879 5315 22937 5321
rect 27154 5312 27160 5324
rect 27212 5312 27218 5364
rect 28810 5244 28816 5296
rect 28868 5244 28874 5296
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1360 5188 1593 5216
rect 1360 5176 1366 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 8386 5216 8392 5228
rect 1903 5188 8392 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 12492 5188 15669 5216
rect 12492 5176 12498 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 21358 5216 21364 5228
rect 17604 5188 21364 5216
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15528 5120 15853 5148
rect 15528 5108 15534 5120
rect 15841 5117 15853 5120
rect 15887 5148 15899 5151
rect 17604 5148 17632 5188
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 22186 5225 22192 5228
rect 22164 5219 22192 5225
rect 22164 5185 22176 5219
rect 22164 5179 22192 5185
rect 22186 5176 22192 5179
rect 22244 5176 22250 5228
rect 22776 5219 22834 5225
rect 22776 5216 22788 5219
rect 22388 5188 22788 5216
rect 15887 5120 17632 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 17678 5108 17684 5160
rect 17736 5108 17742 5160
rect 21376 5148 21404 5176
rect 22388 5148 22416 5188
rect 22776 5185 22788 5188
rect 22822 5185 22834 5219
rect 22776 5179 22834 5185
rect 21376 5120 22416 5148
rect 28721 5151 28779 5157
rect 28721 5117 28733 5151
rect 28767 5148 28779 5151
rect 29638 5148 29644 5160
rect 28767 5120 29644 5148
rect 28767 5117 28779 5120
rect 28721 5111 28779 5117
rect 29638 5108 29644 5120
rect 29696 5108 29702 5160
rect 29733 5151 29791 5157
rect 29733 5117 29745 5151
rect 29779 5148 29791 5151
rect 31386 5148 31392 5160
rect 29779 5120 31392 5148
rect 29779 5117 29791 5120
rect 29733 5111 29791 5117
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 3237 5083 3295 5089
rect 3237 5080 3249 5083
rect 2746 5052 3249 5080
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 2746 5012 2774 5052
rect 3237 5049 3249 5052
rect 3283 5049 3295 5083
rect 3237 5043 3295 5049
rect 1912 4984 2774 5012
rect 16301 5015 16359 5021
rect 1912 4972 1918 4984
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 17862 5012 17868 5024
rect 16347 4984 17868 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 20530 5012 20536 5024
rect 18187 4984 20536 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 22235 5015 22293 5021
rect 22235 4981 22247 5015
rect 22281 5012 22293 5015
rect 22738 5012 22744 5024
rect 22281 4984 22744 5012
rect 22281 4981 22293 4984
rect 22235 4975 22293 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 6822 4808 6828 4820
rect 2915 4780 6828 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 17460 4780 19533 4808
rect 17460 4768 17466 4780
rect 19521 4777 19533 4780
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 20254 4768 20260 4820
rect 20312 4768 20318 4820
rect 24719 4811 24777 4817
rect 24719 4777 24731 4811
rect 24765 4808 24777 4811
rect 28810 4808 28816 4820
rect 24765 4780 28816 4808
rect 24765 4777 24777 4780
rect 24719 4771 24777 4777
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 3513 4743 3571 4749
rect 3513 4740 3525 4743
rect 1596 4712 3525 4740
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 1596 4681 1624 4712
rect 3513 4709 3525 4712
rect 3559 4709 3571 4743
rect 3513 4703 3571 4709
rect 1581 4675 1639 4681
rect 1581 4672 1593 4675
rect 1360 4644 1593 4672
rect 1360 4632 1366 4644
rect 1581 4641 1593 4644
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 10042 4672 10048 4684
rect 1903 4644 10048 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 25869 4675 25927 4681
rect 25869 4641 25881 4675
rect 25915 4672 25927 4675
rect 27522 4672 27528 4684
rect 25915 4644 27528 4672
rect 25915 4641 25927 4644
rect 25869 4635 25927 4641
rect 27522 4632 27528 4644
rect 27580 4632 27586 4684
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2924 4576 3065 4604
rect 2924 4564 2930 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 3099 4576 3341 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20254 4604 20260 4616
rect 19475 4576 20260 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 22066 4576 24628 4604
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 19889 4471 19947 4477
rect 19889 4468 19901 4471
rect 17736 4440 19901 4468
rect 17736 4428 17742 4440
rect 19889 4437 19901 4440
rect 19935 4468 19947 4471
rect 22066 4468 22094 4576
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 22738 4496 22744 4548
rect 22796 4536 22802 4548
rect 25961 4539 26019 4545
rect 25961 4536 25973 4539
rect 22796 4508 25973 4536
rect 22796 4496 22802 4508
rect 25961 4505 25973 4508
rect 26007 4505 26019 4539
rect 25961 4499 26019 4505
rect 26881 4539 26939 4545
rect 26881 4505 26893 4539
rect 26927 4536 26939 4539
rect 37458 4536 37464 4548
rect 26927 4508 37464 4536
rect 26927 4505 26939 4508
rect 26881 4499 26939 4505
rect 37458 4496 37464 4508
rect 37516 4496 37522 4548
rect 19935 4440 22094 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 1394 4224 1400 4276
rect 1452 4224 1458 4276
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1854 4128 1860 4140
rect 1452 4100 1860 4128
rect 1452 4088 1458 4100
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2547 4100 2973 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4212 4100 4261 4128
rect 4212 4088 4218 4100
rect 4249 4097 4261 4100
rect 4295 4128 4307 4131
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4295 4100 4537 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 9674 3992 9680 4004
rect 4111 3964 9680 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3605 3927 3663 3933
rect 3605 3924 3617 3927
rect 3384 3896 3617 3924
rect 3384 3884 3390 3896
rect 3605 3893 3617 3896
rect 3651 3893 3663 3927
rect 3605 3887 3663 3893
rect 15010 3884 15016 3936
rect 15068 3884 15074 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 3973 3723 4031 3729
rect 3973 3689 3985 3723
rect 4019 3720 4031 3723
rect 10594 3720 10600 3732
rect 4019 3692 10600 3720
rect 4019 3689 4031 3692
rect 3973 3683 4031 3689
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 12066 3680 12072 3732
rect 12124 3680 12130 3732
rect 2961 3655 3019 3661
rect 2961 3621 2973 3655
rect 3007 3652 3019 3655
rect 13446 3652 13452 3664
rect 3007 3624 13452 3652
rect 3007 3621 3019 3624
rect 2961 3615 3019 3621
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 31938 3612 31944 3664
rect 31996 3652 32002 3664
rect 31996 3624 39068 3652
rect 31996 3612 32002 3624
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 1581 3587 1639 3593
rect 1581 3584 1593 3587
rect 1360 3556 1593 3584
rect 1360 3544 1366 3556
rect 1581 3553 1593 3556
rect 1627 3584 1639 3587
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 1627 3556 4629 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 25774 3544 25780 3596
rect 25832 3584 25838 3596
rect 25832 3556 35894 3584
rect 25832 3544 25838 3556
rect 658 3476 664 3528
rect 716 3516 722 3528
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 716 3488 1869 3516
rect 716 3476 722 3488
rect 1857 3485 1869 3488
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3145 3519 3203 3525
rect 3145 3516 3157 3519
rect 2924 3488 3157 3516
rect 2924 3476 2930 3488
rect 3145 3485 3157 3488
rect 3191 3516 3203 3519
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3191 3488 3433 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 4120 3488 4169 3516
rect 4120 3476 4126 3488
rect 4157 3485 4169 3488
rect 4203 3516 4215 3519
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4203 3488 4445 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 12066 3516 12072 3528
rect 11563 3488 12072 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 35710 3476 35716 3528
rect 35768 3476 35774 3528
rect 35866 3516 35894 3556
rect 37829 3519 37887 3525
rect 37829 3516 37841 3519
rect 35866 3488 37841 3516
rect 37829 3485 37841 3488
rect 37875 3485 37887 3519
rect 37829 3479 37887 3485
rect 32122 3408 32128 3460
rect 32180 3448 32186 3460
rect 39040 3457 39068 3624
rect 36909 3451 36967 3457
rect 36909 3448 36921 3451
rect 32180 3420 36921 3448
rect 32180 3408 32186 3420
rect 36909 3417 36921 3420
rect 36955 3417 36967 3451
rect 36909 3411 36967 3417
rect 39025 3451 39083 3457
rect 39025 3417 39037 3451
rect 39071 3448 39083 3451
rect 49418 3448 49424 3460
rect 39071 3420 49424 3448
rect 39071 3417 39083 3420
rect 39025 3411 39083 3417
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 31754 3340 31760 3392
rect 31812 3380 31818 3392
rect 33594 3380 33600 3392
rect 31812 3352 33600 3380
rect 31812 3340 31818 3352
rect 33594 3340 33600 3352
rect 33652 3340 33658 3392
rect 36924 3380 36952 3411
rect 49418 3408 49424 3420
rect 49476 3408 49482 3460
rect 44082 3380 44088 3392
rect 36924 3352 44088 3380
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3145 4031 3179
rect 3973 3139 4031 3145
rect 3988 3108 4016 3139
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 9824 3148 14013 3176
rect 9824 3136 9830 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 14001 3139 14059 3145
rect 25498 3136 25504 3188
rect 25556 3136 25562 3188
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 28169 3179 28227 3185
rect 28169 3176 28181 3179
rect 27580 3148 28181 3176
rect 27580 3136 27586 3148
rect 28169 3145 28181 3148
rect 28215 3145 28227 3179
rect 28169 3139 28227 3145
rect 29638 3136 29644 3188
rect 29696 3176 29702 3188
rect 33505 3179 33563 3185
rect 33505 3176 33517 3179
rect 29696 3148 33517 3176
rect 29696 3136 29702 3148
rect 33505 3145 33517 3148
rect 33551 3145 33563 3179
rect 33505 3139 33563 3145
rect 33594 3136 33600 3188
rect 33652 3176 33658 3188
rect 33652 3148 38608 3176
rect 33652 3136 33658 3148
rect 10318 3108 10324 3120
rect 3988 3080 4660 3108
rect 10258 3080 10324 3108
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3040 1639 3043
rect 2774 3040 2780 3052
rect 1627 3012 2780 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3326 3040 3332 3052
rect 2915 3012 3332 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 4632 3049 4660 3080
rect 10318 3068 10324 3080
rect 10376 3108 10382 3120
rect 10781 3111 10839 3117
rect 10781 3108 10793 3111
rect 10376 3080 10793 3108
rect 10376 3068 10382 3080
rect 10781 3077 10793 3080
rect 10827 3077 10839 3111
rect 10781 3071 10839 3077
rect 12618 3068 12624 3120
rect 12676 3068 12682 3120
rect 13909 3111 13967 3117
rect 13909 3077 13921 3111
rect 13955 3108 13967 3111
rect 15470 3108 15476 3120
rect 13955 3080 15476 3108
rect 13955 3077 13967 3080
rect 13909 3071 13967 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15565 3111 15623 3117
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 17678 3108 17684 3120
rect 15611 3080 17684 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 31386 3068 31392 3120
rect 31444 3108 31450 3120
rect 31444 3080 35296 3108
rect 31444 3068 31450 3080
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3559 3012 4169 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 5307 3012 6561 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7892 3012 8769 3040
rect 7892 3000 7898 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17920 3012 18337 3040
rect 17920 3000 17926 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20530 3000 20536 3052
rect 20588 3000 20594 3052
rect 25685 3043 25743 3049
rect 25685 3009 25697 3043
rect 25731 3040 25743 3043
rect 26234 3040 26240 3052
rect 25731 3012 26240 3040
rect 25731 3009 25743 3012
rect 25685 3003 25743 3009
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 28350 3000 28356 3052
rect 28408 3000 28414 3052
rect 31018 3000 31024 3052
rect 31076 3000 31082 3052
rect 33686 3000 33692 3052
rect 33744 3000 33750 3052
rect 35268 3049 35296 3080
rect 35253 3043 35311 3049
rect 35253 3009 35265 3043
rect 35299 3009 35311 3043
rect 35253 3003 35311 3009
rect 37458 3000 37464 3052
rect 37516 3000 37522 3052
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 5626 2972 5632 2984
rect 1903 2944 5632 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 7239 2944 9045 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 17402 2972 17408 2984
rect 10551 2944 17408 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 35158 2932 35164 2984
rect 35216 2972 35222 2984
rect 38580 2981 38608 3148
rect 36449 2975 36507 2981
rect 36449 2972 36461 2975
rect 35216 2944 36461 2972
rect 35216 2932 35222 2944
rect 36449 2941 36461 2944
rect 36495 2941 36507 2975
rect 36449 2935 36507 2941
rect 38565 2975 38623 2981
rect 38565 2941 38577 2975
rect 38611 2972 38623 2975
rect 46750 2972 46756 2984
rect 38611 2944 46756 2972
rect 38611 2941 38623 2944
rect 38565 2935 38623 2941
rect 10060 2876 10916 2904
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 10060 2836 10088 2876
rect 8352 2808 10088 2836
rect 10888 2836 10916 2876
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 12492 2876 15761 2904
rect 12492 2864 12498 2876
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 30282 2864 30288 2916
rect 30340 2904 30346 2916
rect 30837 2907 30895 2913
rect 30837 2904 30849 2907
rect 30340 2876 30849 2904
rect 30340 2864 30346 2876
rect 30837 2873 30849 2876
rect 30883 2873 30895 2907
rect 36464 2904 36492 2935
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 41414 2904 41420 2916
rect 36464 2876 41420 2904
rect 30837 2867 30895 2873
rect 41414 2864 41420 2876
rect 41472 2864 41478 2916
rect 12713 2839 12771 2845
rect 12713 2836 12725 2839
rect 10888 2808 12725 2836
rect 8352 2796 8358 2808
rect 12713 2805 12725 2808
rect 12759 2805 12771 2839
rect 12713 2799 12771 2805
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17494 2836 17500 2848
rect 16899 2808 17500 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 20070 2836 20076 2848
rect 18187 2808 20076 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20349 2839 20407 2845
rect 20349 2805 20361 2839
rect 20395 2836 20407 2839
rect 21910 2836 21916 2848
rect 20395 2808 21916 2836
rect 20395 2805 20407 2808
rect 20349 2799 20407 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 9582 2632 9588 2644
rect 2915 2604 9588 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 26234 2592 26240 2644
rect 26292 2592 26298 2644
rect 28350 2592 28356 2644
rect 28408 2632 28414 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 28408 2604 28917 2632
rect 28408 2592 28414 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 28905 2595 28963 2601
rect 31018 2592 31024 2644
rect 31076 2632 31082 2644
rect 31573 2635 31631 2641
rect 31573 2632 31585 2635
rect 31076 2604 31585 2632
rect 31076 2592 31082 2604
rect 31573 2601 31585 2604
rect 31619 2601 31631 2635
rect 31573 2595 31631 2601
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 34241 2635 34299 2641
rect 34241 2632 34253 2635
rect 33744 2604 34253 2632
rect 33744 2592 33750 2604
rect 34241 2601 34253 2604
rect 34287 2601 34299 2635
rect 34241 2595 34299 2601
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 3513 2567 3571 2573
rect 3513 2564 3525 2567
rect 2832 2536 3525 2564
rect 2832 2524 2838 2536
rect 3513 2533 3525 2536
rect 3559 2533 3571 2567
rect 11606 2564 11612 2576
rect 3513 2527 3571 2533
rect 5184 2536 11612 2564
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1268 2468 1593 2496
rect 1268 2456 1274 2468
rect 1581 2465 1593 2468
rect 1627 2496 1639 2499
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 1627 2468 3801 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4120 2468 4629 2496
rect 4120 2456 4126 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 5184 2428 5212 2536
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6788 2468 7297 2496
rect 6788 2456 6794 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9456 2468 9965 2496
rect 9456 2456 9462 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12124 2468 12633 2496
rect 12124 2456 12130 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 14792 2468 15301 2496
rect 14792 2456 14798 2468
rect 15289 2465 15301 2468
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17957 2499 18015 2505
rect 17957 2496 17969 2499
rect 17460 2468 17969 2496
rect 17460 2456 17466 2468
rect 17957 2465 17969 2468
rect 18003 2465 18015 2499
rect 17957 2459 18015 2465
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22796 2468 23121 2496
rect 22796 2456 22802 2468
rect 23109 2465 23121 2468
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 31570 2456 31576 2508
rect 31628 2496 31634 2508
rect 36357 2499 36415 2505
rect 36357 2496 36369 2499
rect 31628 2468 36369 2496
rect 31628 2456 31634 2468
rect 36357 2465 36369 2468
rect 36403 2465 36415 2499
rect 36357 2459 36415 2465
rect 4387 2400 5212 2428
rect 7009 2431 7067 2437
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8294 2428 8300 2440
rect 7055 2400 8300 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 3068 2360 3096 2391
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12434 2428 12440 2440
rect 12391 2400 12440 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 15010 2388 15016 2440
rect 15068 2388 15074 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 21968 2400 22661 2428
rect 21968 2388 21974 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 22649 2391 22707 2397
rect 25424 2400 25605 2428
rect 3329 2363 3387 2369
rect 3329 2360 3341 2363
rect 1360 2332 3341 2360
rect 1360 2320 1366 2332
rect 3329 2329 3341 2332
rect 3375 2329 3387 2363
rect 3329 2323 3387 2329
rect 25424 2304 25452 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 28261 2431 28319 2437
rect 28261 2428 28273 2431
rect 25593 2391 25651 2397
rect 27908 2400 28273 2428
rect 1811 2295 1869 2301
rect 1811 2261 1823 2295
rect 1857 2292 1869 2295
rect 5994 2292 6000 2304
rect 1857 2264 6000 2292
rect 1857 2261 1869 2264
rect 1811 2255 1869 2261
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 25317 2295 25375 2301
rect 25317 2261 25329 2295
rect 25363 2292 25375 2295
rect 25406 2292 25412 2304
rect 25363 2264 25412 2292
rect 25363 2261 25375 2264
rect 25317 2255 25375 2261
rect 25406 2252 25412 2264
rect 25464 2252 25470 2304
rect 27798 2252 27804 2304
rect 27856 2292 27862 2304
rect 27908 2301 27936 2400
rect 28261 2397 28273 2400
rect 28307 2397 28319 2431
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 28261 2391 28319 2397
rect 30760 2400 30941 2428
rect 30760 2304 30788 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 30929 2391 30987 2397
rect 33428 2400 33609 2428
rect 33428 2304 33456 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36136 2400 37289 2428
rect 36136 2388 36142 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 27893 2295 27951 2301
rect 27893 2292 27905 2295
rect 27856 2264 27905 2292
rect 27856 2252 27862 2264
rect 27893 2261 27905 2264
rect 27939 2261 27951 2295
rect 27893 2255 27951 2261
rect 30653 2295 30711 2301
rect 30653 2261 30665 2295
rect 30699 2292 30711 2295
rect 30742 2292 30748 2304
rect 30699 2264 30748 2292
rect 30699 2261 30711 2264
rect 30653 2255 30711 2261
rect 30742 2252 30748 2264
rect 30800 2252 30806 2304
rect 33321 2295 33379 2301
rect 33321 2261 33333 2295
rect 33367 2292 33379 2295
rect 33410 2292 33416 2304
rect 33367 2264 33416 2292
rect 33367 2261 33379 2264
rect 33321 2255 33379 2261
rect 33410 2252 33416 2264
rect 33468 2252 33474 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 9680 25576 9732 25628
rect 21824 25576 21876 25628
rect 4804 25508 4856 25560
rect 21180 25508 21232 25560
rect 10048 25440 10100 25492
rect 28448 25440 28500 25492
rect 12072 25372 12124 25424
rect 33968 25372 34020 25424
rect 12348 25304 12400 25356
rect 26424 25304 26476 25356
rect 17776 25236 17828 25288
rect 34336 25236 34388 25288
rect 15384 25168 15436 25220
rect 33600 25168 33652 25220
rect 10600 25100 10652 25152
rect 30380 25100 30432 25152
rect 4068 25032 4120 25084
rect 8484 25032 8536 25084
rect 12716 25032 12768 25084
rect 33416 25032 33468 25084
rect 15016 24964 15068 25016
rect 30012 24964 30064 25016
rect 30564 24964 30616 25016
rect 32864 24964 32916 25016
rect 14832 24896 14884 24948
rect 39304 24896 39356 24948
rect 10784 24828 10836 24880
rect 36544 24828 36596 24880
rect 4068 24760 4120 24812
rect 8300 24760 8352 24812
rect 11704 24760 11756 24812
rect 21916 24760 21968 24812
rect 22652 24760 22704 24812
rect 28540 24760 28592 24812
rect 28632 24760 28684 24812
rect 32312 24760 32364 24812
rect 4252 24692 4304 24744
rect 6460 24624 6512 24676
rect 13636 24624 13688 24676
rect 25044 24692 25096 24744
rect 30564 24692 30616 24744
rect 17132 24624 17184 24676
rect 18604 24624 18656 24676
rect 25964 24624 26016 24676
rect 27528 24624 27580 24676
rect 31300 24624 31352 24676
rect 24124 24556 24176 24608
rect 25228 24556 25280 24608
rect 29000 24556 29052 24608
rect 29092 24556 29144 24608
rect 35532 24692 35584 24744
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 2780 24352 2832 24404
rect 5264 24352 5316 24404
rect 16488 24352 16540 24404
rect 572 24284 624 24336
rect 3516 24216 3568 24268
rect 1032 24148 1084 24200
rect 9312 24284 9364 24336
rect 7380 24216 7432 24268
rect 4252 24148 4304 24200
rect 664 24080 716 24132
rect 6828 24148 6880 24200
rect 8576 24148 8628 24200
rect 14740 24284 14792 24336
rect 10048 24148 10100 24200
rect 3700 24012 3752 24064
rect 6276 24012 6328 24064
rect 9680 24012 9732 24064
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 14372 24216 14424 24268
rect 18972 24352 19024 24404
rect 19064 24352 19116 24404
rect 18696 24216 18748 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 22100 24216 22152 24268
rect 25044 24259 25096 24268
rect 25044 24225 25053 24259
rect 25053 24225 25087 24259
rect 25087 24225 25096 24259
rect 25044 24216 25096 24225
rect 25228 24259 25280 24268
rect 25228 24225 25237 24259
rect 25237 24225 25271 24259
rect 25271 24225 25280 24259
rect 25228 24216 25280 24225
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 14556 24148 14608 24200
rect 16580 24148 16632 24200
rect 18420 24148 18472 24200
rect 19892 24148 19944 24200
rect 21916 24148 21968 24200
rect 23572 24148 23624 24200
rect 24768 24148 24820 24200
rect 13820 24080 13872 24132
rect 15292 24080 15344 24132
rect 17132 24123 17184 24132
rect 17132 24089 17141 24123
rect 17141 24089 17175 24123
rect 17175 24089 17184 24123
rect 17132 24080 17184 24089
rect 18512 24080 18564 24132
rect 19524 24080 19576 24132
rect 23940 24080 23992 24132
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 17040 24012 17092 24064
rect 20168 24012 20220 24064
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 24952 24055 25004 24064
rect 24952 24021 24961 24055
rect 24961 24021 24995 24055
rect 24995 24021 25004 24055
rect 24952 24012 25004 24021
rect 25964 24080 26016 24132
rect 26976 24352 27028 24404
rect 29460 24352 29512 24404
rect 29552 24352 29604 24404
rect 31024 24352 31076 24404
rect 31300 24352 31352 24404
rect 34796 24352 34848 24404
rect 27344 24284 27396 24336
rect 30748 24284 30800 24336
rect 33784 24284 33836 24336
rect 41512 24352 41564 24404
rect 42616 24352 42668 24404
rect 44732 24395 44784 24404
rect 44732 24361 44741 24395
rect 44741 24361 44775 24395
rect 44775 24361 44784 24395
rect 44732 24352 44784 24361
rect 35624 24284 35676 24336
rect 37096 24284 37148 24336
rect 43444 24284 43496 24336
rect 44916 24284 44968 24336
rect 27988 24148 28040 24200
rect 28448 24148 28500 24200
rect 26424 24080 26476 24132
rect 31024 24191 31076 24200
rect 31024 24157 31033 24191
rect 31033 24157 31067 24191
rect 31067 24157 31076 24191
rect 31024 24148 31076 24157
rect 31392 24148 31444 24200
rect 29920 24080 29972 24132
rect 33324 24148 33376 24200
rect 32036 24080 32088 24132
rect 35532 24216 35584 24268
rect 47676 24216 47728 24268
rect 35072 24148 35124 24200
rect 35624 24080 35676 24132
rect 36360 24148 36412 24200
rect 38476 24191 38528 24200
rect 38476 24157 38485 24191
rect 38485 24157 38519 24191
rect 38519 24157 38528 24191
rect 38476 24148 38528 24157
rect 38936 24148 38988 24200
rect 39948 24148 40000 24200
rect 40224 24148 40276 24200
rect 44180 24148 44232 24200
rect 44732 24148 44784 24200
rect 45560 24148 45612 24200
rect 45928 24191 45980 24200
rect 45928 24157 45937 24191
rect 45937 24157 45971 24191
rect 45971 24157 45980 24191
rect 45928 24148 45980 24157
rect 46020 24148 46072 24200
rect 47308 24148 47360 24200
rect 48596 24191 48648 24200
rect 48596 24157 48605 24191
rect 48605 24157 48639 24191
rect 48639 24157 48648 24191
rect 48596 24148 48648 24157
rect 43352 24080 43404 24132
rect 25872 24012 25924 24064
rect 26240 24055 26292 24064
rect 26240 24021 26249 24055
rect 26249 24021 26283 24055
rect 26283 24021 26292 24055
rect 26240 24012 26292 24021
rect 26332 24012 26384 24064
rect 27344 24012 27396 24064
rect 28356 24012 28408 24064
rect 29184 24055 29236 24064
rect 29184 24021 29193 24055
rect 29193 24021 29227 24055
rect 29227 24021 29236 24055
rect 29184 24012 29236 24021
rect 30656 24012 30708 24064
rect 33508 24012 33560 24064
rect 34152 24012 34204 24064
rect 35992 24012 36044 24064
rect 37372 24012 37424 24064
rect 38476 24012 38528 24064
rect 40684 24055 40736 24064
rect 40684 24021 40693 24055
rect 40693 24021 40727 24055
rect 40727 24021 40736 24055
rect 40684 24012 40736 24021
rect 41420 24012 41472 24064
rect 42800 24012 42852 24064
rect 45376 24055 45428 24064
rect 45376 24021 45385 24055
rect 45385 24021 45419 24055
rect 45419 24021 45428 24055
rect 45376 24012 45428 24021
rect 48688 24012 48740 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 4160 23740 4212 23792
rect 6460 23851 6512 23860
rect 6460 23817 6469 23851
rect 6469 23817 6503 23851
rect 6503 23817 6512 23851
rect 6460 23808 6512 23817
rect 9772 23808 9824 23860
rect 23940 23808 23992 23860
rect 24952 23808 25004 23860
rect 28448 23808 28500 23860
rect 7380 23740 7432 23792
rect 9956 23740 10008 23792
rect 12532 23740 12584 23792
rect 15752 23740 15804 23792
rect 756 23672 808 23724
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 7656 23672 7708 23724
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 11796 23672 11848 23724
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 17132 23740 17184 23792
rect 19248 23740 19300 23792
rect 19524 23740 19576 23792
rect 21180 23783 21232 23792
rect 21180 23749 21189 23783
rect 21189 23749 21223 23783
rect 21223 23749 21232 23783
rect 21180 23740 21232 23749
rect 23664 23740 23716 23792
rect 26424 23740 26476 23792
rect 29184 23808 29236 23860
rect 16948 23672 17000 23724
rect 17500 23672 17552 23724
rect 18696 23715 18748 23724
rect 18696 23681 18705 23715
rect 18705 23681 18739 23715
rect 18739 23681 18748 23715
rect 18696 23672 18748 23681
rect 20444 23672 20496 23724
rect 29460 23672 29512 23724
rect 30656 23783 30708 23792
rect 30656 23749 30665 23783
rect 30665 23749 30699 23783
rect 30699 23749 30708 23783
rect 30656 23740 30708 23749
rect 30748 23740 30800 23792
rect 32036 23740 32088 23792
rect 33508 23783 33560 23792
rect 33508 23749 33517 23783
rect 33517 23749 33551 23783
rect 33551 23749 33560 23783
rect 33508 23740 33560 23749
rect 33692 23783 33744 23792
rect 33692 23749 33701 23783
rect 33701 23749 33735 23783
rect 33735 23749 33744 23783
rect 33692 23740 33744 23749
rect 3976 23604 4028 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 6276 23604 6328 23656
rect 848 23536 900 23588
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 1768 23468 1820 23520
rect 7564 23604 7616 23656
rect 18328 23604 18380 23656
rect 19064 23604 19116 23656
rect 3792 23468 3844 23520
rect 9680 23468 9732 23520
rect 11520 23511 11572 23520
rect 11520 23477 11529 23511
rect 11529 23477 11563 23511
rect 11563 23477 11572 23511
rect 11520 23468 11572 23477
rect 11888 23511 11940 23520
rect 11888 23477 11897 23511
rect 11897 23477 11931 23511
rect 11931 23477 11940 23511
rect 11888 23468 11940 23477
rect 17040 23536 17092 23588
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 24400 23604 24452 23656
rect 25872 23604 25924 23656
rect 27160 23647 27212 23656
rect 27160 23613 27169 23647
rect 27169 23613 27203 23647
rect 27203 23613 27212 23647
rect 27160 23604 27212 23613
rect 27436 23647 27488 23656
rect 27436 23613 27445 23647
rect 27445 23613 27479 23647
rect 27479 23613 27488 23647
rect 27436 23604 27488 23613
rect 32220 23672 32272 23724
rect 32312 23715 32364 23724
rect 32312 23681 32321 23715
rect 32321 23681 32355 23715
rect 32355 23681 32364 23715
rect 32312 23672 32364 23681
rect 34796 23808 34848 23860
rect 39304 23851 39356 23860
rect 39304 23817 39313 23851
rect 39313 23817 39347 23851
rect 39347 23817 39356 23851
rect 39304 23808 39356 23817
rect 39948 23808 40000 23860
rect 45928 23808 45980 23860
rect 47308 23808 47360 23860
rect 47676 23808 47728 23860
rect 35992 23783 36044 23792
rect 35992 23749 36001 23783
rect 36001 23749 36035 23783
rect 36035 23749 36044 23783
rect 35992 23740 36044 23749
rect 36176 23783 36228 23792
rect 36176 23749 36185 23783
rect 36185 23749 36219 23783
rect 36219 23749 36228 23783
rect 36176 23740 36228 23749
rect 38476 23783 38528 23792
rect 38476 23749 38485 23783
rect 38485 23749 38519 23783
rect 38519 23749 38528 23783
rect 38476 23740 38528 23749
rect 38660 23783 38712 23792
rect 38660 23749 38669 23783
rect 38669 23749 38703 23783
rect 38703 23749 38712 23783
rect 38660 23740 38712 23749
rect 40684 23740 40736 23792
rect 34520 23672 34572 23724
rect 36820 23715 36872 23724
rect 36820 23681 36829 23715
rect 36829 23681 36863 23715
rect 36863 23681 36872 23715
rect 36820 23672 36872 23681
rect 37096 23672 37148 23724
rect 39580 23672 39632 23724
rect 44088 23740 44140 23792
rect 42616 23715 42668 23724
rect 42616 23681 42625 23715
rect 42625 23681 42659 23715
rect 42659 23681 42668 23715
rect 42616 23672 42668 23681
rect 26332 23536 26384 23588
rect 14280 23468 14332 23520
rect 16580 23468 16632 23520
rect 17684 23468 17736 23520
rect 18696 23468 18748 23520
rect 20076 23468 20128 23520
rect 20536 23468 20588 23520
rect 21640 23511 21692 23520
rect 21640 23477 21649 23511
rect 21649 23477 21683 23511
rect 21683 23477 21692 23511
rect 21640 23468 21692 23477
rect 23756 23511 23808 23520
rect 23756 23477 23765 23511
rect 23765 23477 23799 23511
rect 23799 23477 23808 23511
rect 23756 23468 23808 23477
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 28540 23536 28592 23588
rect 29460 23536 29512 23588
rect 28908 23511 28960 23520
rect 28908 23477 28917 23511
rect 28917 23477 28951 23511
rect 28951 23477 28960 23511
rect 28908 23468 28960 23477
rect 30104 23511 30156 23520
rect 30104 23477 30113 23511
rect 30113 23477 30147 23511
rect 30147 23477 30156 23511
rect 30104 23468 30156 23477
rect 30380 23468 30432 23520
rect 43812 23672 43864 23724
rect 44640 23672 44692 23724
rect 46664 23672 46716 23724
rect 47768 23672 47820 23724
rect 48320 23672 48372 23724
rect 48688 23715 48740 23724
rect 48688 23681 48697 23715
rect 48697 23681 48731 23715
rect 48731 23681 48740 23715
rect 48688 23672 48740 23681
rect 31024 23536 31076 23588
rect 31852 23511 31904 23520
rect 31852 23477 31861 23511
rect 31861 23477 31895 23511
rect 31895 23477 31904 23511
rect 31852 23468 31904 23477
rect 32772 23468 32824 23520
rect 34060 23468 34112 23520
rect 35440 23511 35492 23520
rect 35440 23477 35449 23511
rect 35449 23477 35483 23511
rect 35483 23477 35492 23511
rect 35440 23468 35492 23477
rect 37004 23468 37056 23520
rect 44916 23536 44968 23588
rect 40592 23511 40644 23520
rect 40592 23477 40601 23511
rect 40601 23477 40635 23511
rect 40635 23477 40644 23511
rect 40592 23468 40644 23477
rect 44364 23511 44416 23520
rect 44364 23477 44373 23511
rect 44373 23477 44407 23511
rect 44407 23477 44416 23511
rect 44364 23468 44416 23477
rect 45008 23511 45060 23520
rect 45008 23477 45017 23511
rect 45017 23477 45051 23511
rect 45051 23477 45060 23511
rect 45008 23468 45060 23477
rect 45744 23511 45796 23520
rect 45744 23477 45753 23511
rect 45753 23477 45787 23511
rect 45787 23477 45796 23511
rect 45744 23468 45796 23477
rect 46940 23511 46992 23520
rect 46940 23477 46949 23511
rect 46949 23477 46983 23511
rect 46983 23477 46992 23511
rect 46940 23468 46992 23477
rect 48688 23468 48740 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 3608 23307 3660 23316
rect 3608 23273 3617 23307
rect 3617 23273 3651 23307
rect 3651 23273 3660 23307
rect 3608 23264 3660 23273
rect 3700 23264 3752 23316
rect 7748 23264 7800 23316
rect 12256 23264 12308 23316
rect 13820 23264 13872 23316
rect 8760 23196 8812 23248
rect 19064 23196 19116 23248
rect 23296 23264 23348 23316
rect 23848 23264 23900 23316
rect 4068 23128 4120 23180
rect 4988 23128 5040 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 12440 23128 12492 23180
rect 13268 23171 13320 23180
rect 13268 23137 13277 23171
rect 13277 23137 13311 23171
rect 13311 23137 13320 23171
rect 13268 23128 13320 23137
rect 15844 23128 15896 23180
rect 17408 23128 17460 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 23756 23196 23808 23248
rect 20720 23128 20772 23180
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 7196 23103 7248 23112
rect 7196 23069 7205 23103
rect 7205 23069 7239 23103
rect 7239 23069 7248 23103
rect 7196 23060 7248 23069
rect 8944 23060 8996 23112
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 4528 23035 4580 23044
rect 4528 23001 4537 23035
rect 4537 23001 4571 23035
rect 4571 23001 4580 23035
rect 4528 22992 4580 23001
rect 4804 22992 4856 23044
rect 9496 22992 9548 23044
rect 4160 22967 4212 22976
rect 4160 22933 4169 22967
rect 4169 22933 4203 22967
rect 4203 22933 4212 22967
rect 4160 22924 4212 22933
rect 7104 22924 7156 22976
rect 9036 22967 9088 22976
rect 9036 22933 9045 22967
rect 9045 22933 9079 22967
rect 9079 22933 9088 22967
rect 12256 22992 12308 23044
rect 9036 22924 9088 22933
rect 11520 22924 11572 22976
rect 11980 22924 12032 22976
rect 12624 22924 12676 22976
rect 12808 22924 12860 22976
rect 13636 22992 13688 23044
rect 14372 23035 14424 23044
rect 14372 23001 14381 23035
rect 14381 23001 14415 23035
rect 14415 23001 14424 23035
rect 14372 22992 14424 23001
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15476 23060 15528 23069
rect 16856 23060 16908 23112
rect 18512 23060 18564 23112
rect 19800 23060 19852 23112
rect 21732 23060 21784 23112
rect 23664 23060 23716 23112
rect 28540 23264 28592 23316
rect 29000 23307 29052 23316
rect 29000 23273 29009 23307
rect 29009 23273 29043 23307
rect 29043 23273 29052 23307
rect 29000 23264 29052 23273
rect 29460 23264 29512 23316
rect 29828 23264 29880 23316
rect 30104 23264 30156 23316
rect 31852 23264 31904 23316
rect 32220 23264 32272 23316
rect 33876 23264 33928 23316
rect 38568 23264 38620 23316
rect 44180 23264 44232 23316
rect 44640 23307 44692 23316
rect 44640 23273 44649 23307
rect 44649 23273 44683 23307
rect 44683 23273 44692 23307
rect 44640 23264 44692 23273
rect 48596 23264 48648 23316
rect 27252 23171 27304 23180
rect 27252 23137 27261 23171
rect 27261 23137 27295 23171
rect 27295 23137 27304 23171
rect 27252 23128 27304 23137
rect 28908 23128 28960 23180
rect 32496 23196 32548 23248
rect 37096 23196 37148 23248
rect 29368 23060 29420 23112
rect 16948 22992 17000 23044
rect 17040 22992 17092 23044
rect 20352 23035 20404 23044
rect 20352 23001 20361 23035
rect 20361 23001 20395 23035
rect 20395 23001 20404 23035
rect 20352 22992 20404 23001
rect 21640 22992 21692 23044
rect 30748 23128 30800 23180
rect 31944 23128 31996 23180
rect 36820 23128 36872 23180
rect 40592 23128 40644 23180
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 32404 23060 32456 23112
rect 32680 23060 32732 23112
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 17224 22924 17276 22976
rect 22284 22924 22336 22976
rect 23388 22924 23440 22976
rect 24124 22924 24176 22976
rect 24676 22924 24728 22976
rect 25872 22924 25924 22976
rect 26792 22924 26844 22976
rect 26976 22924 27028 22976
rect 29920 22992 29972 23044
rect 31484 22992 31536 23044
rect 33140 23103 33192 23112
rect 33140 23069 33149 23103
rect 33149 23069 33183 23103
rect 33183 23069 33192 23103
rect 33140 23060 33192 23069
rect 33876 23060 33928 23112
rect 34152 23060 34204 23112
rect 35440 23060 35492 23112
rect 35716 23060 35768 23112
rect 40316 23103 40368 23112
rect 40316 23069 40325 23103
rect 40325 23069 40359 23103
rect 40359 23069 40368 23103
rect 40316 23060 40368 23069
rect 43260 23060 43312 23112
rect 44364 23060 44416 23112
rect 32036 22924 32088 22976
rect 32588 22967 32640 22976
rect 32588 22933 32597 22967
rect 32597 22933 32631 22967
rect 32631 22933 32640 22967
rect 32588 22924 32640 22933
rect 32956 22967 33008 22976
rect 32956 22933 32965 22967
rect 32965 22933 32999 22967
rect 32999 22933 33008 22967
rect 32956 22924 33008 22933
rect 33508 22992 33560 23044
rect 35624 23035 35676 23044
rect 35624 23001 35633 23035
rect 35633 23001 35667 23035
rect 35667 23001 35676 23035
rect 35624 22992 35676 23001
rect 47860 23060 47912 23112
rect 48504 23060 48556 23112
rect 37464 22924 37516 22976
rect 38752 22967 38804 22976
rect 38752 22933 38761 22967
rect 38761 22933 38795 22967
rect 38795 22933 38804 22967
rect 38752 22924 38804 22933
rect 48412 22992 48464 23044
rect 46848 22967 46900 22976
rect 46848 22933 46857 22967
rect 46857 22933 46891 22967
rect 46891 22933 46900 22967
rect 46848 22924 46900 22933
rect 47492 22924 47544 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 14464 22720 14516 22772
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 20352 22720 20404 22772
rect 25136 22720 25188 22772
rect 26332 22720 26384 22772
rect 26424 22763 26476 22772
rect 26424 22729 26433 22763
rect 26433 22729 26467 22763
rect 26467 22729 26476 22763
rect 26424 22720 26476 22729
rect 27528 22720 27580 22772
rect 3792 22627 3844 22636
rect 3792 22593 3801 22627
rect 3801 22593 3835 22627
rect 3835 22593 3844 22627
rect 3792 22584 3844 22593
rect 2872 22516 2924 22568
rect 3332 22516 3384 22568
rect 6368 22584 6420 22636
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 7012 22652 7064 22704
rect 6828 22584 6880 22636
rect 7840 22584 7892 22636
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 10968 22652 11020 22704
rect 12808 22652 12860 22704
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 16672 22652 16724 22704
rect 18512 22652 18564 22704
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 12256 22584 12308 22636
rect 13820 22584 13872 22636
rect 15016 22627 15068 22636
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 19432 22584 19484 22636
rect 20076 22652 20128 22704
rect 21640 22652 21692 22704
rect 23664 22652 23716 22704
rect 24676 22652 24728 22704
rect 26608 22652 26660 22704
rect 26792 22695 26844 22704
rect 26792 22661 26801 22695
rect 26801 22661 26835 22695
rect 26835 22661 26844 22695
rect 26792 22652 26844 22661
rect 22836 22584 22888 22636
rect 25504 22584 25556 22636
rect 26976 22584 27028 22636
rect 28356 22652 28408 22704
rect 28540 22652 28592 22704
rect 30748 22720 30800 22772
rect 31024 22763 31076 22772
rect 31024 22729 31033 22763
rect 31033 22729 31067 22763
rect 31067 22729 31076 22763
rect 31024 22720 31076 22729
rect 29368 22652 29420 22704
rect 30840 22652 30892 22704
rect 32956 22720 33008 22772
rect 33416 22720 33468 22772
rect 34520 22720 34572 22772
rect 37464 22763 37516 22772
rect 37464 22729 37473 22763
rect 37473 22729 37507 22763
rect 37507 22729 37516 22763
rect 37464 22720 37516 22729
rect 40868 22720 40920 22772
rect 31392 22652 31444 22704
rect 36544 22695 36596 22704
rect 36544 22661 36553 22695
rect 36553 22661 36587 22695
rect 36587 22661 36596 22695
rect 36544 22652 36596 22661
rect 43260 22763 43312 22772
rect 43260 22729 43269 22763
rect 43269 22729 43303 22763
rect 43303 22729 43312 22763
rect 43260 22720 43312 22729
rect 47768 22763 47820 22772
rect 47768 22729 47777 22763
rect 47777 22729 47811 22763
rect 47811 22729 47820 22763
rect 47768 22720 47820 22729
rect 3700 22448 3752 22500
rect 4620 22448 4672 22500
rect 5724 22448 5776 22500
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 8760 22516 8812 22568
rect 11980 22516 12032 22568
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 9588 22448 9640 22500
rect 10876 22448 10928 22500
rect 13268 22516 13320 22568
rect 16856 22559 16908 22568
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 18604 22516 18656 22568
rect 20536 22516 20588 22568
rect 21732 22516 21784 22568
rect 23388 22559 23440 22568
rect 23388 22525 23397 22559
rect 23397 22525 23431 22559
rect 23431 22525 23440 22559
rect 23388 22516 23440 22525
rect 23756 22516 23808 22568
rect 24032 22516 24084 22568
rect 27252 22516 27304 22568
rect 29920 22584 29972 22636
rect 5356 22380 5408 22432
rect 11336 22380 11388 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 13452 22380 13504 22432
rect 19156 22380 19208 22432
rect 20168 22380 20220 22432
rect 20352 22380 20404 22432
rect 20720 22380 20772 22432
rect 23572 22380 23624 22432
rect 23940 22380 23992 22432
rect 26056 22448 26108 22500
rect 27528 22448 27580 22500
rect 28356 22559 28408 22568
rect 28356 22525 28365 22559
rect 28365 22525 28399 22559
rect 28399 22525 28408 22559
rect 28356 22516 28408 22525
rect 29000 22516 29052 22568
rect 31024 22584 31076 22636
rect 31760 22584 31812 22636
rect 32220 22584 32272 22636
rect 32496 22584 32548 22636
rect 33416 22584 33468 22636
rect 34244 22627 34296 22636
rect 34244 22593 34253 22627
rect 34253 22593 34287 22627
rect 34287 22593 34296 22627
rect 34244 22584 34296 22593
rect 34520 22627 34572 22636
rect 34520 22593 34529 22627
rect 34529 22593 34563 22627
rect 34563 22593 34572 22627
rect 34520 22584 34572 22593
rect 34704 22584 34756 22636
rect 35716 22584 35768 22636
rect 29644 22448 29696 22500
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 25688 22380 25740 22432
rect 28264 22380 28316 22432
rect 28356 22380 28408 22432
rect 29828 22380 29880 22432
rect 30564 22491 30616 22500
rect 30564 22457 30573 22491
rect 30573 22457 30607 22491
rect 30607 22457 30616 22491
rect 30564 22448 30616 22457
rect 31852 22448 31904 22500
rect 32036 22448 32088 22500
rect 41420 22584 41472 22636
rect 42800 22584 42852 22636
rect 46848 22584 46900 22636
rect 48320 22627 48372 22636
rect 48320 22593 48329 22627
rect 48329 22593 48363 22627
rect 48363 22593 48372 22627
rect 48320 22584 48372 22593
rect 49056 22627 49108 22636
rect 49056 22593 49065 22627
rect 49065 22593 49099 22627
rect 49099 22593 49108 22627
rect 49056 22584 49108 22593
rect 32128 22380 32180 22432
rect 34520 22380 34572 22432
rect 39580 22423 39632 22432
rect 39580 22389 39589 22423
rect 39589 22389 39623 22423
rect 39623 22389 39632 22423
rect 39580 22380 39632 22389
rect 40684 22423 40736 22432
rect 40684 22389 40693 22423
rect 40693 22389 40727 22423
rect 40727 22389 40736 22423
rect 40684 22380 40736 22389
rect 41328 22423 41380 22432
rect 41328 22389 41337 22423
rect 41337 22389 41371 22423
rect 41371 22389 41380 22423
rect 41328 22380 41380 22389
rect 48504 22423 48556 22432
rect 48504 22389 48513 22423
rect 48513 22389 48547 22423
rect 48547 22389 48556 22423
rect 48504 22380 48556 22389
rect 49240 22423 49292 22432
rect 49240 22389 49249 22423
rect 49249 22389 49283 22423
rect 49283 22389 49292 22423
rect 49240 22380 49292 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 3700 22176 3752 22228
rect 3424 22108 3476 22160
rect 4160 22108 4212 22160
rect 1308 22040 1360 22092
rect 4068 22040 4120 22092
rect 3792 21972 3844 22024
rect 4252 21972 4304 22024
rect 11888 22176 11940 22228
rect 11980 22176 12032 22228
rect 14556 22176 14608 22228
rect 16396 22176 16448 22228
rect 23388 22176 23440 22228
rect 6736 22108 6788 22160
rect 9036 22151 9088 22160
rect 9036 22117 9045 22151
rect 9045 22117 9079 22151
rect 9079 22117 9088 22151
rect 9036 22108 9088 22117
rect 11060 22108 11112 22160
rect 11336 22108 11388 22160
rect 18512 22108 18564 22160
rect 19064 22108 19116 22160
rect 21732 22108 21784 22160
rect 21824 22108 21876 22160
rect 22284 22151 22336 22160
rect 22284 22117 22293 22151
rect 22293 22117 22327 22151
rect 22327 22117 22336 22151
rect 22284 22108 22336 22117
rect 6644 21972 6696 22024
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 8392 21972 8444 22024
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 10048 22040 10100 22092
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 15108 22040 15160 22092
rect 19432 22040 19484 22092
rect 23572 22040 23624 22092
rect 26056 22176 26108 22228
rect 26240 22176 26292 22228
rect 27528 22219 27580 22228
rect 27528 22185 27537 22219
rect 27537 22185 27571 22219
rect 27571 22185 27580 22219
rect 27528 22176 27580 22185
rect 24308 22108 24360 22160
rect 24768 22040 24820 22092
rect 27252 22108 27304 22160
rect 29828 22219 29880 22228
rect 29828 22185 29837 22219
rect 29837 22185 29871 22219
rect 29871 22185 29880 22219
rect 29828 22176 29880 22185
rect 28264 22108 28316 22160
rect 31944 22176 31996 22228
rect 26056 22040 26108 22092
rect 28448 22040 28500 22092
rect 10416 21972 10468 22024
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 14556 21972 14608 22024
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 15384 21972 15436 22024
rect 18512 21972 18564 22024
rect 18880 21972 18932 22024
rect 12716 21904 12768 21956
rect 17500 21904 17552 21956
rect 6092 21879 6144 21888
rect 6092 21845 6101 21879
rect 6101 21845 6135 21879
rect 6135 21845 6144 21879
rect 6092 21836 6144 21845
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9956 21836 10008 21888
rect 10508 21836 10560 21888
rect 10784 21836 10836 21888
rect 11520 21836 11572 21888
rect 14648 21836 14700 21888
rect 14924 21879 14976 21888
rect 14924 21845 14933 21879
rect 14933 21845 14967 21879
rect 14967 21845 14976 21879
rect 14924 21836 14976 21845
rect 18788 21836 18840 21888
rect 19340 21836 19392 21888
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 20260 21904 20312 21956
rect 24676 21972 24728 22024
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 28632 21972 28684 22024
rect 29184 22083 29236 22092
rect 29184 22049 29193 22083
rect 29193 22049 29227 22083
rect 29227 22049 29236 22083
rect 29184 22040 29236 22049
rect 29552 21972 29604 22024
rect 30748 22083 30800 22092
rect 30748 22049 30757 22083
rect 30757 22049 30791 22083
rect 30791 22049 30800 22083
rect 30748 22040 30800 22049
rect 31208 22108 31260 22160
rect 35440 22176 35492 22228
rect 42800 22176 42852 22228
rect 49240 22176 49292 22228
rect 32128 22108 32180 22160
rect 32588 22108 32640 22160
rect 32680 22108 32732 22160
rect 37648 22108 37700 22160
rect 32036 22083 32088 22092
rect 32036 22049 32045 22083
rect 32045 22049 32079 22083
rect 32079 22049 32088 22083
rect 32036 22040 32088 22049
rect 32220 22083 32272 22092
rect 32220 22049 32229 22083
rect 32229 22049 32263 22083
rect 32263 22049 32272 22083
rect 32220 22040 32272 22049
rect 22928 21904 22980 21956
rect 22192 21836 22244 21888
rect 23296 21879 23348 21888
rect 23296 21845 23305 21879
rect 23305 21845 23339 21879
rect 23339 21845 23348 21879
rect 23296 21836 23348 21845
rect 24952 21947 25004 21956
rect 24952 21913 24961 21947
rect 24961 21913 24995 21947
rect 24995 21913 25004 21947
rect 24952 21904 25004 21913
rect 26056 21947 26108 21956
rect 26056 21913 26065 21947
rect 26065 21913 26099 21947
rect 26099 21913 26108 21947
rect 26056 21904 26108 21913
rect 26516 21904 26568 21956
rect 28908 21904 28960 21956
rect 25688 21836 25740 21888
rect 25964 21836 26016 21888
rect 28724 21836 28776 21888
rect 29368 21836 29420 21888
rect 29644 21904 29696 21956
rect 30380 21836 30432 21888
rect 31392 21947 31444 21956
rect 31392 21913 31401 21947
rect 31401 21913 31435 21947
rect 31435 21913 31444 21947
rect 31392 21904 31444 21913
rect 32036 21904 32088 21956
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 32864 22015 32916 22024
rect 32864 21981 32873 22015
rect 32873 21981 32907 22015
rect 32907 21981 32916 22015
rect 32864 21972 32916 21981
rect 38752 22040 38804 22092
rect 48412 22151 48464 22160
rect 48412 22117 48421 22151
rect 48421 22117 48455 22151
rect 48455 22117 48464 22151
rect 48412 22108 48464 22117
rect 34060 21972 34112 22024
rect 35164 21972 35216 22024
rect 35440 21972 35492 22024
rect 37280 21972 37332 22024
rect 48688 21972 48740 22024
rect 49056 22015 49108 22024
rect 49056 21981 49065 22015
rect 49065 21981 49099 22015
rect 49099 21981 49108 22015
rect 49056 21972 49108 21981
rect 34980 21947 35032 21956
rect 34980 21913 34989 21947
rect 34989 21913 35023 21947
rect 35023 21913 35032 21947
rect 34980 21904 35032 21913
rect 36452 21904 36504 21956
rect 40316 21904 40368 21956
rect 33600 21836 33652 21888
rect 35072 21879 35124 21888
rect 35072 21845 35081 21879
rect 35081 21845 35115 21879
rect 35115 21845 35124 21879
rect 35072 21836 35124 21845
rect 35624 21879 35676 21888
rect 35624 21845 35633 21879
rect 35633 21845 35667 21879
rect 35667 21845 35676 21879
rect 35624 21836 35676 21845
rect 36268 21879 36320 21888
rect 36268 21845 36277 21879
rect 36277 21845 36311 21879
rect 36311 21845 36320 21879
rect 36268 21836 36320 21845
rect 37464 21879 37516 21888
rect 37464 21845 37473 21879
rect 37473 21845 37507 21879
rect 37507 21845 37516 21879
rect 37464 21836 37516 21845
rect 37556 21836 37608 21888
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 3424 21632 3476 21684
rect 3608 21632 3660 21684
rect 4252 21632 4304 21684
rect 9220 21632 9272 21684
rect 9404 21675 9456 21684
rect 9404 21641 9413 21675
rect 9413 21641 9447 21675
rect 9447 21641 9456 21675
rect 9404 21632 9456 21641
rect 10692 21632 10744 21684
rect 10968 21675 11020 21684
rect 10968 21641 10977 21675
rect 10977 21641 11011 21675
rect 11011 21641 11020 21675
rect 10968 21632 11020 21641
rect 15936 21632 15988 21684
rect 16028 21675 16080 21684
rect 16028 21641 16037 21675
rect 16037 21641 16071 21675
rect 16071 21641 16080 21675
rect 16028 21632 16080 21641
rect 16212 21632 16264 21684
rect 5816 21564 5868 21616
rect 6276 21564 6328 21616
rect 7564 21564 7616 21616
rect 1124 21428 1176 21480
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 7104 21496 7156 21548
rect 1952 21428 2004 21480
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 5540 21428 5592 21480
rect 6460 21428 6512 21480
rect 6184 21360 6236 21412
rect 3332 21292 3384 21344
rect 3608 21292 3660 21344
rect 5540 21292 5592 21344
rect 6460 21335 6512 21344
rect 6460 21301 6469 21335
rect 6469 21301 6503 21335
rect 6503 21301 6512 21335
rect 6460 21292 6512 21301
rect 7104 21335 7156 21344
rect 7104 21301 7113 21335
rect 7113 21301 7147 21335
rect 7147 21301 7156 21335
rect 7104 21292 7156 21301
rect 9036 21496 9088 21548
rect 10140 21496 10192 21548
rect 7932 21428 7984 21480
rect 10324 21496 10376 21548
rect 10876 21428 10928 21480
rect 12716 21564 12768 21616
rect 13452 21564 13504 21616
rect 13820 21564 13872 21616
rect 14648 21564 14700 21616
rect 20812 21675 20864 21684
rect 20812 21641 20821 21675
rect 20821 21641 20855 21675
rect 20855 21641 20864 21675
rect 20812 21632 20864 21641
rect 21640 21632 21692 21684
rect 21732 21632 21784 21684
rect 23388 21632 23440 21684
rect 24400 21632 24452 21684
rect 25964 21675 26016 21684
rect 25964 21641 25973 21675
rect 25973 21641 26007 21675
rect 26007 21641 26016 21675
rect 25964 21632 26016 21641
rect 26608 21632 26660 21684
rect 27620 21675 27672 21684
rect 27620 21641 27629 21675
rect 27629 21641 27663 21675
rect 27663 21641 27672 21675
rect 27620 21632 27672 21641
rect 35624 21632 35676 21684
rect 12532 21496 12584 21548
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 23572 21564 23624 21616
rect 23940 21564 23992 21616
rect 24124 21564 24176 21616
rect 10416 21360 10468 21412
rect 18604 21496 18656 21548
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 8944 21292 8996 21344
rect 11152 21292 11204 21344
rect 11520 21292 11572 21344
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 15568 21403 15620 21412
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 16672 21360 16724 21412
rect 18604 21360 18656 21412
rect 12808 21292 12860 21344
rect 14004 21292 14056 21344
rect 15016 21292 15068 21344
rect 18696 21292 18748 21344
rect 18972 21471 19024 21480
rect 18972 21437 18981 21471
rect 18981 21437 19015 21471
rect 19015 21437 19024 21471
rect 18972 21428 19024 21437
rect 19064 21428 19116 21480
rect 20812 21496 20864 21548
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 26516 21496 26568 21548
rect 24676 21428 24728 21480
rect 29000 21564 29052 21616
rect 29184 21564 29236 21616
rect 31760 21564 31812 21616
rect 31852 21564 31904 21616
rect 35440 21607 35492 21616
rect 35440 21573 35449 21607
rect 35449 21573 35483 21607
rect 35483 21573 35492 21607
rect 35440 21564 35492 21573
rect 27804 21471 27856 21480
rect 27804 21437 27813 21471
rect 27813 21437 27847 21471
rect 27847 21437 27856 21471
rect 27804 21428 27856 21437
rect 28356 21428 28408 21480
rect 20260 21360 20312 21412
rect 22744 21360 22796 21412
rect 19432 21292 19484 21344
rect 19708 21292 19760 21344
rect 25872 21360 25924 21412
rect 26056 21360 26108 21412
rect 27896 21360 27948 21412
rect 25228 21292 25280 21344
rect 25688 21292 25740 21344
rect 27620 21292 27672 21344
rect 30380 21360 30432 21412
rect 32128 21428 32180 21480
rect 32404 21539 32456 21548
rect 32404 21505 32413 21539
rect 32413 21505 32447 21539
rect 32447 21505 32456 21539
rect 32404 21496 32456 21505
rect 32772 21496 32824 21548
rect 33416 21496 33468 21548
rect 47584 21496 47636 21548
rect 37372 21428 37424 21480
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 31392 21360 31444 21412
rect 32312 21360 32364 21412
rect 33876 21360 33928 21412
rect 30196 21335 30248 21344
rect 30196 21301 30205 21335
rect 30205 21301 30239 21335
rect 30239 21301 30248 21335
rect 30196 21292 30248 21301
rect 30656 21335 30708 21344
rect 30656 21301 30665 21335
rect 30665 21301 30699 21335
rect 30699 21301 30708 21335
rect 30656 21292 30708 21301
rect 31576 21292 31628 21344
rect 32036 21292 32088 21344
rect 32404 21292 32456 21344
rect 32772 21292 32824 21344
rect 33968 21292 34020 21344
rect 34980 21292 35032 21344
rect 47584 21335 47636 21344
rect 47584 21301 47593 21335
rect 47593 21301 47627 21335
rect 47627 21301 47636 21335
rect 47584 21292 47636 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 3424 21131 3476 21140
rect 3424 21097 3433 21131
rect 3433 21097 3467 21131
rect 3467 21097 3476 21131
rect 3424 21088 3476 21097
rect 4068 21020 4120 21072
rect 4252 20995 4304 21004
rect 4252 20961 4261 20995
rect 4261 20961 4295 20995
rect 4295 20961 4304 20995
rect 4252 20952 4304 20961
rect 7288 20952 7340 21004
rect 1860 20884 1912 20936
rect 3332 20884 3384 20936
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 2780 20859 2832 20868
rect 2780 20825 2789 20859
rect 2789 20825 2823 20859
rect 2823 20825 2832 20859
rect 2780 20816 2832 20825
rect 5264 20816 5316 20868
rect 6184 20816 6236 20868
rect 7472 21088 7524 21140
rect 7564 21020 7616 21072
rect 7748 20952 7800 21004
rect 11796 21020 11848 21072
rect 13820 21088 13872 21140
rect 14464 21088 14516 21140
rect 16580 21088 16632 21140
rect 14924 21020 14976 21072
rect 7472 20884 7524 20936
rect 9680 20995 9732 21004
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9680 20952 9732 20961
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 11704 20884 11756 20936
rect 11980 20927 12032 20936
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 15016 20952 15068 21004
rect 17224 21020 17276 21072
rect 16212 20995 16264 21004
rect 16212 20961 16221 20995
rect 16221 20961 16255 20995
rect 16255 20961 16264 20995
rect 16212 20952 16264 20961
rect 16396 20995 16448 21004
rect 16396 20961 16405 20995
rect 16405 20961 16439 20995
rect 16439 20961 16448 20995
rect 16396 20952 16448 20961
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 18788 20995 18840 21004
rect 18788 20961 18797 20995
rect 18797 20961 18831 20995
rect 18831 20961 18840 20995
rect 18788 20952 18840 20961
rect 21640 21063 21692 21072
rect 21640 21029 21649 21063
rect 21649 21029 21683 21063
rect 21683 21029 21692 21063
rect 21640 21020 21692 21029
rect 22284 21088 22336 21140
rect 23480 21020 23532 21072
rect 23756 21088 23808 21140
rect 26056 21088 26108 21140
rect 26516 21088 26568 21140
rect 28908 21088 28960 21140
rect 29736 21088 29788 21140
rect 31852 21088 31904 21140
rect 33324 21088 33376 21140
rect 49056 21088 49108 21140
rect 19708 20995 19760 21004
rect 19708 20961 19717 20995
rect 19717 20961 19751 20995
rect 19751 20961 19760 20995
rect 19708 20952 19760 20961
rect 20076 20952 20128 21004
rect 22652 20952 22704 21004
rect 23572 20952 23624 21004
rect 24400 21020 24452 21072
rect 25780 21020 25832 21072
rect 23848 20995 23900 21004
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 25320 20995 25372 21004
rect 25320 20961 25329 20995
rect 25329 20961 25363 20995
rect 25363 20961 25372 20995
rect 25320 20952 25372 20961
rect 26056 20995 26108 21004
rect 26056 20961 26065 20995
rect 26065 20961 26099 20995
rect 26099 20961 26108 20995
rect 26056 20952 26108 20961
rect 27804 21020 27856 21072
rect 35716 21020 35768 21072
rect 27712 20952 27764 21004
rect 29920 20952 29972 21004
rect 30012 20995 30064 21004
rect 30012 20961 30021 20995
rect 30021 20961 30055 20995
rect 30055 20961 30064 20995
rect 30012 20952 30064 20961
rect 30104 20952 30156 21004
rect 32588 20952 32640 21004
rect 34152 20952 34204 21004
rect 15200 20884 15252 20936
rect 17500 20884 17552 20936
rect 18880 20884 18932 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 23296 20884 23348 20936
rect 28448 20884 28500 20936
rect 29828 20884 29880 20936
rect 32128 20884 32180 20936
rect 10324 20816 10376 20868
rect 11336 20859 11388 20868
rect 11336 20825 11345 20859
rect 11345 20825 11379 20859
rect 11379 20825 11388 20859
rect 11336 20816 11388 20825
rect 17868 20816 17920 20868
rect 5908 20748 5960 20800
rect 7564 20791 7616 20800
rect 7564 20757 7573 20791
rect 7573 20757 7607 20791
rect 7607 20757 7616 20791
rect 7564 20748 7616 20757
rect 8852 20748 8904 20800
rect 11428 20791 11480 20800
rect 11428 20757 11437 20791
rect 11437 20757 11471 20791
rect 11471 20757 11480 20791
rect 11428 20748 11480 20757
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 14740 20748 14792 20800
rect 15752 20791 15804 20800
rect 15752 20757 15761 20791
rect 15761 20757 15795 20791
rect 15795 20757 15804 20791
rect 15752 20748 15804 20757
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 17040 20748 17092 20800
rect 19984 20816 20036 20868
rect 20996 20816 21048 20868
rect 21640 20816 21692 20868
rect 22376 20816 22428 20868
rect 23388 20816 23440 20868
rect 26240 20816 26292 20868
rect 26424 20816 26476 20868
rect 18328 20748 18380 20800
rect 20536 20748 20588 20800
rect 22284 20748 22336 20800
rect 22652 20748 22704 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 23756 20748 23808 20800
rect 30656 20816 30708 20868
rect 27896 20748 27948 20800
rect 29000 20748 29052 20800
rect 32036 20859 32088 20868
rect 32036 20825 32045 20859
rect 32045 20825 32079 20859
rect 32079 20825 32088 20859
rect 32036 20816 32088 20825
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 34060 20791 34112 20800
rect 34060 20757 34069 20791
rect 34069 20757 34103 20791
rect 34103 20757 34112 20791
rect 34060 20748 34112 20757
rect 46204 20748 46256 20800
rect 47492 20748 47544 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 6920 20544 6972 20596
rect 4620 20476 4672 20528
rect 9496 20544 9548 20596
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 940 20340 992 20392
rect 6000 20408 6052 20460
rect 6092 20408 6144 20460
rect 2044 20383 2096 20392
rect 2044 20349 2053 20383
rect 2053 20349 2087 20383
rect 2087 20349 2096 20383
rect 2044 20340 2096 20349
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 7564 20408 7616 20460
rect 10140 20476 10192 20528
rect 11796 20519 11848 20528
rect 11796 20485 11805 20519
rect 11805 20485 11839 20519
rect 11839 20485 11848 20519
rect 11796 20476 11848 20485
rect 12440 20476 12492 20528
rect 13544 20476 13596 20528
rect 14004 20519 14056 20528
rect 14004 20485 14013 20519
rect 14013 20485 14047 20519
rect 14047 20485 14056 20519
rect 14004 20476 14056 20485
rect 14464 20476 14516 20528
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 16948 20544 17000 20596
rect 18880 20587 18932 20596
rect 18880 20553 18889 20587
rect 18889 20553 18923 20587
rect 18923 20553 18932 20587
rect 18880 20544 18932 20553
rect 19432 20544 19484 20596
rect 7288 20340 7340 20392
rect 6092 20272 6144 20324
rect 6184 20272 6236 20324
rect 7472 20272 7524 20324
rect 8944 20340 8996 20392
rect 9128 20272 9180 20324
rect 3884 20204 3936 20256
rect 4068 20204 4120 20256
rect 7288 20204 7340 20256
rect 8208 20204 8260 20256
rect 8392 20204 8444 20256
rect 10968 20340 11020 20392
rect 15200 20340 15252 20392
rect 16672 20408 16724 20460
rect 15476 20315 15528 20324
rect 15476 20281 15485 20315
rect 15485 20281 15519 20315
rect 15519 20281 15528 20315
rect 15476 20272 15528 20281
rect 9680 20204 9732 20256
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 11336 20204 11388 20256
rect 12532 20247 12584 20256
rect 12532 20213 12541 20247
rect 12541 20213 12575 20247
rect 12575 20213 12584 20247
rect 12532 20204 12584 20213
rect 13452 20247 13504 20256
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 13636 20247 13688 20256
rect 13636 20213 13645 20247
rect 13645 20213 13679 20247
rect 13679 20213 13688 20247
rect 13636 20204 13688 20213
rect 13728 20204 13780 20256
rect 17592 20408 17644 20460
rect 16948 20272 17000 20324
rect 17960 20340 18012 20392
rect 20996 20476 21048 20528
rect 21916 20476 21968 20528
rect 23388 20587 23440 20596
rect 23388 20553 23397 20587
rect 23397 20553 23431 20587
rect 23431 20553 23440 20587
rect 23388 20544 23440 20553
rect 24952 20544 25004 20596
rect 25504 20544 25556 20596
rect 26056 20544 26108 20596
rect 27068 20544 27120 20596
rect 30840 20544 30892 20596
rect 31668 20544 31720 20596
rect 31760 20544 31812 20596
rect 32128 20544 32180 20596
rect 32220 20544 32272 20596
rect 26424 20519 26476 20528
rect 26424 20485 26433 20519
rect 26433 20485 26467 20519
rect 26467 20485 26476 20519
rect 26424 20476 26476 20485
rect 29092 20476 29144 20528
rect 37464 20476 37516 20528
rect 23204 20408 23256 20460
rect 26332 20408 26384 20460
rect 27344 20408 27396 20460
rect 31944 20408 31996 20460
rect 19616 20272 19668 20324
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 20628 20340 20680 20392
rect 24676 20340 24728 20392
rect 25688 20272 25740 20324
rect 28356 20383 28408 20392
rect 22744 20204 22796 20256
rect 26516 20204 26568 20256
rect 27712 20204 27764 20256
rect 28356 20349 28365 20383
rect 28365 20349 28399 20383
rect 28399 20349 28408 20383
rect 28356 20340 28408 20349
rect 30196 20340 30248 20392
rect 30288 20340 30340 20392
rect 31024 20272 31076 20324
rect 31944 20272 31996 20324
rect 28356 20204 28408 20256
rect 30564 20247 30616 20256
rect 30564 20213 30573 20247
rect 30573 20213 30607 20247
rect 30607 20213 30616 20247
rect 30564 20204 30616 20213
rect 30932 20204 30984 20256
rect 31576 20247 31628 20256
rect 31576 20213 31585 20247
rect 31585 20213 31619 20247
rect 31619 20213 31628 20247
rect 31576 20204 31628 20213
rect 31760 20247 31812 20256
rect 31760 20213 31769 20247
rect 31769 20213 31803 20247
rect 31803 20213 31812 20247
rect 31760 20204 31812 20213
rect 32128 20247 32180 20256
rect 32128 20213 32137 20247
rect 32137 20213 32171 20247
rect 32171 20213 32180 20247
rect 32128 20204 32180 20213
rect 32496 20247 32548 20256
rect 32496 20213 32505 20247
rect 32505 20213 32539 20247
rect 32539 20213 32548 20247
rect 32496 20204 32548 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 3424 20000 3476 20052
rect 5264 20000 5316 20052
rect 6276 20043 6328 20052
rect 6276 20009 6285 20043
rect 6285 20009 6319 20043
rect 6319 20009 6328 20043
rect 6276 20000 6328 20009
rect 7748 20000 7800 20052
rect 8300 20000 8352 20052
rect 5448 19864 5500 19916
rect 8944 19864 8996 19916
rect 4252 19796 4304 19848
rect 10048 20000 10100 20052
rect 11796 20000 11848 20052
rect 12440 19932 12492 19984
rect 2872 19728 2924 19780
rect 3516 19728 3568 19780
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 3884 19703 3936 19712
rect 3884 19669 3893 19703
rect 3893 19669 3927 19703
rect 3927 19669 3936 19703
rect 3884 19660 3936 19669
rect 5080 19728 5132 19780
rect 5264 19728 5316 19780
rect 6644 19660 6696 19712
rect 7472 19728 7524 19780
rect 10416 19796 10468 19848
rect 12072 19864 12124 19916
rect 12716 19864 12768 19916
rect 11244 19796 11296 19848
rect 13360 20000 13412 20052
rect 17960 20000 18012 20052
rect 19892 20000 19944 20052
rect 20720 20000 20772 20052
rect 14280 19975 14332 19984
rect 14280 19941 14289 19975
rect 14289 19941 14323 19975
rect 14323 19941 14332 19975
rect 14280 19932 14332 19941
rect 14464 19975 14516 19984
rect 14464 19941 14473 19975
rect 14473 19941 14507 19975
rect 14507 19941 14516 19975
rect 14464 19932 14516 19941
rect 17040 19932 17092 19984
rect 17224 19975 17276 19984
rect 17224 19941 17233 19975
rect 17233 19941 17267 19975
rect 17267 19941 17276 19975
rect 17224 19932 17276 19941
rect 15476 19864 15528 19916
rect 16028 19864 16080 19916
rect 19340 19932 19392 19984
rect 27804 20000 27856 20052
rect 29736 20043 29788 20052
rect 29736 20009 29745 20043
rect 29745 20009 29779 20043
rect 29779 20009 29788 20043
rect 29736 20000 29788 20009
rect 29920 20000 29972 20052
rect 31024 20000 31076 20052
rect 35164 20000 35216 20052
rect 49240 20000 49292 20052
rect 18972 19864 19024 19916
rect 19432 19864 19484 19916
rect 19616 19864 19668 19916
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 21548 19864 21600 19916
rect 23848 19907 23900 19916
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 26148 19864 26200 19916
rect 26516 19864 26568 19916
rect 8576 19660 8628 19712
rect 10140 19728 10192 19780
rect 12716 19728 12768 19780
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 18328 19796 18380 19848
rect 19064 19796 19116 19848
rect 19708 19796 19760 19848
rect 22376 19796 22428 19848
rect 24952 19796 25004 19848
rect 25780 19796 25832 19848
rect 27620 19864 27672 19916
rect 29000 19796 29052 19848
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 41328 19796 41380 19848
rect 14832 19728 14884 19780
rect 11152 19660 11204 19712
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 13268 19660 13320 19712
rect 13820 19703 13872 19712
rect 13820 19669 13829 19703
rect 13829 19669 13863 19703
rect 13863 19669 13872 19703
rect 13820 19660 13872 19669
rect 14464 19660 14516 19712
rect 16672 19728 16724 19780
rect 19984 19728 20036 19780
rect 20996 19728 21048 19780
rect 23572 19728 23624 19780
rect 25504 19728 25556 19780
rect 26424 19728 26476 19780
rect 26608 19728 26660 19780
rect 16396 19660 16448 19712
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 19892 19660 19944 19712
rect 20076 19660 20128 19712
rect 20720 19660 20772 19712
rect 22376 19660 22428 19712
rect 23296 19703 23348 19712
rect 23296 19669 23305 19703
rect 23305 19669 23339 19703
rect 23339 19669 23348 19703
rect 23296 19660 23348 19669
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 23848 19660 23900 19712
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 29828 19728 29880 19780
rect 27804 19660 27856 19712
rect 29092 19660 29144 19712
rect 30196 19660 30248 19712
rect 30748 19703 30800 19712
rect 30748 19669 30757 19703
rect 30757 19669 30791 19703
rect 30791 19669 30800 19703
rect 30748 19660 30800 19669
rect 31024 19660 31076 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 4344 19431 4396 19440
rect 4344 19397 4353 19431
rect 4353 19397 4387 19431
rect 4387 19397 4396 19431
rect 4344 19388 4396 19397
rect 5448 19456 5500 19508
rect 5724 19499 5776 19508
rect 5724 19465 5733 19499
rect 5733 19465 5767 19499
rect 5767 19465 5776 19499
rect 5724 19456 5776 19465
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 4896 19320 4948 19372
rect 5724 19320 5776 19372
rect 6460 19456 6512 19508
rect 10324 19456 10376 19508
rect 11888 19456 11940 19508
rect 14556 19456 14608 19508
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 16580 19456 16632 19508
rect 16948 19456 17000 19508
rect 17040 19456 17092 19508
rect 7104 19388 7156 19440
rect 8484 19388 8536 19440
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 2688 19184 2740 19236
rect 6644 19320 6696 19372
rect 8760 19320 8812 19372
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 11612 19320 11664 19372
rect 11980 19388 12032 19440
rect 12072 19388 12124 19440
rect 13268 19388 13320 19440
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 19432 19456 19484 19508
rect 23296 19456 23348 19508
rect 26240 19456 26292 19508
rect 27712 19499 27764 19508
rect 27712 19465 27721 19499
rect 27721 19465 27755 19499
rect 27755 19465 27764 19499
rect 27712 19456 27764 19465
rect 19340 19388 19392 19440
rect 13912 19320 13964 19372
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 13636 19252 13688 19304
rect 14004 19252 14056 19304
rect 14924 19295 14976 19304
rect 14924 19261 14933 19295
rect 14933 19261 14967 19295
rect 14967 19261 14976 19295
rect 14924 19252 14976 19261
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 15844 19320 15896 19372
rect 5724 19116 5776 19168
rect 8300 19184 8352 19236
rect 9496 19184 9548 19236
rect 11704 19184 11756 19236
rect 13360 19184 13412 19236
rect 13820 19227 13872 19236
rect 13820 19193 13829 19227
rect 13829 19193 13863 19227
rect 13863 19193 13872 19227
rect 13820 19184 13872 19193
rect 6920 19116 6972 19168
rect 10876 19116 10928 19168
rect 10968 19116 11020 19168
rect 14372 19227 14424 19236
rect 14372 19193 14381 19227
rect 14381 19193 14415 19227
rect 14415 19193 14424 19227
rect 14372 19184 14424 19193
rect 15108 19184 15160 19236
rect 16304 19252 16356 19304
rect 16856 19252 16908 19304
rect 17408 19363 17460 19372
rect 17408 19329 17417 19363
rect 17417 19329 17451 19363
rect 17451 19329 17460 19363
rect 17408 19320 17460 19329
rect 17868 19320 17920 19372
rect 19064 19320 19116 19372
rect 20076 19388 20128 19440
rect 21088 19320 21140 19372
rect 21732 19388 21784 19440
rect 22652 19388 22704 19440
rect 23480 19388 23532 19440
rect 25320 19388 25372 19440
rect 28172 19388 28224 19440
rect 21548 19320 21600 19372
rect 23756 19320 23808 19372
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 20628 19252 20680 19304
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 16764 19184 16816 19236
rect 20996 19184 21048 19236
rect 23848 19252 23900 19304
rect 24860 19252 24912 19304
rect 15016 19116 15068 19168
rect 17868 19116 17920 19168
rect 18788 19116 18840 19168
rect 21180 19116 21232 19168
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 22100 19116 22152 19168
rect 27344 19320 27396 19372
rect 30380 19456 30432 19508
rect 34704 19456 34756 19508
rect 29092 19388 29144 19440
rect 31024 19388 31076 19440
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 26976 19295 27028 19304
rect 26976 19261 26985 19295
rect 26985 19261 27019 19295
rect 27019 19261 27028 19295
rect 26976 19252 27028 19261
rect 27160 19252 27212 19304
rect 30656 19363 30708 19372
rect 30656 19329 30665 19363
rect 30665 19329 30699 19363
rect 30699 19329 30708 19363
rect 30656 19320 30708 19329
rect 27988 19252 28040 19304
rect 25320 19184 25372 19236
rect 25412 19184 25464 19236
rect 30472 19252 30524 19304
rect 23388 19116 23440 19168
rect 23572 19116 23624 19168
rect 26792 19116 26844 19168
rect 27528 19116 27580 19168
rect 28172 19116 28224 19168
rect 28632 19116 28684 19168
rect 30288 19116 30340 19168
rect 30932 19159 30984 19168
rect 30932 19125 30941 19159
rect 30941 19125 30975 19159
rect 30975 19125 30984 19159
rect 30932 19116 30984 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 1400 18776 1452 18828
rect 9772 18912 9824 18964
rect 11060 18912 11112 18964
rect 9128 18844 9180 18896
rect 10140 18844 10192 18896
rect 8484 18776 8536 18828
rect 10232 18776 10284 18828
rect 11060 18776 11112 18828
rect 11244 18776 11296 18828
rect 4252 18708 4304 18760
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 9772 18708 9824 18760
rect 10876 18708 10928 18760
rect 15016 18912 15068 18964
rect 13728 18844 13780 18896
rect 14464 18844 14516 18896
rect 13544 18819 13596 18828
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 14832 18776 14884 18828
rect 4988 18640 5040 18692
rect 6184 18640 6236 18692
rect 6460 18640 6512 18692
rect 7104 18683 7156 18692
rect 7104 18649 7113 18683
rect 7113 18649 7147 18683
rect 7147 18649 7156 18683
rect 7104 18640 7156 18649
rect 7564 18640 7616 18692
rect 2504 18572 2556 18624
rect 3608 18615 3660 18624
rect 3608 18581 3617 18615
rect 3617 18581 3651 18615
rect 3651 18581 3660 18615
rect 3608 18572 3660 18581
rect 5080 18572 5132 18624
rect 8852 18640 8904 18692
rect 10048 18640 10100 18692
rect 12808 18683 12860 18692
rect 12808 18649 12817 18683
rect 12817 18649 12851 18683
rect 12851 18649 12860 18683
rect 12808 18640 12860 18649
rect 22008 18912 22060 18964
rect 22652 18912 22704 18964
rect 23296 18912 23348 18964
rect 25412 18912 25464 18964
rect 25504 18912 25556 18964
rect 17592 18844 17644 18896
rect 21088 18844 21140 18896
rect 22468 18844 22520 18896
rect 26700 18844 26752 18896
rect 46940 18912 46992 18964
rect 16212 18776 16264 18828
rect 16672 18776 16724 18828
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 18604 18819 18656 18828
rect 18604 18785 18613 18819
rect 18613 18785 18647 18819
rect 18647 18785 18656 18819
rect 18604 18776 18656 18785
rect 16764 18708 16816 18760
rect 19708 18776 19760 18828
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 21824 18776 21876 18828
rect 15016 18640 15068 18692
rect 15476 18683 15528 18692
rect 15476 18649 15485 18683
rect 15485 18649 15519 18683
rect 15519 18649 15528 18683
rect 15476 18640 15528 18649
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 10508 18572 10560 18624
rect 11704 18572 11756 18624
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 14832 18572 14884 18624
rect 15292 18572 15344 18624
rect 16396 18572 16448 18624
rect 20076 18640 20128 18692
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17960 18572 18012 18624
rect 18696 18572 18748 18624
rect 19340 18615 19392 18624
rect 19340 18581 19349 18615
rect 19349 18581 19383 18615
rect 19383 18581 19392 18615
rect 19340 18572 19392 18581
rect 20812 18615 20864 18624
rect 20812 18581 20821 18615
rect 20821 18581 20855 18615
rect 20855 18581 20864 18615
rect 20812 18572 20864 18581
rect 21732 18640 21784 18692
rect 23664 18776 23716 18828
rect 25780 18776 25832 18828
rect 29828 18776 29880 18828
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 23848 18708 23900 18760
rect 26792 18708 26844 18760
rect 27620 18751 27672 18760
rect 27620 18717 27629 18751
rect 27629 18717 27663 18751
rect 27663 18717 27672 18751
rect 27620 18708 27672 18717
rect 27712 18708 27764 18760
rect 30564 18708 30616 18760
rect 22100 18572 22152 18624
rect 23848 18572 23900 18624
rect 24032 18572 24084 18624
rect 25688 18683 25740 18692
rect 25688 18649 25697 18683
rect 25697 18649 25731 18683
rect 25731 18649 25740 18683
rect 25688 18640 25740 18649
rect 29092 18640 29144 18692
rect 30932 18640 30984 18692
rect 29644 18572 29696 18624
rect 29736 18615 29788 18624
rect 29736 18581 29745 18615
rect 29745 18581 29779 18615
rect 29779 18581 29788 18615
rect 29736 18572 29788 18581
rect 30104 18615 30156 18624
rect 30104 18581 30113 18615
rect 30113 18581 30147 18615
rect 30147 18581 30156 18615
rect 30104 18572 30156 18581
rect 43444 18572 43496 18624
rect 48504 18572 48556 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 5908 18300 5960 18352
rect 5632 18275 5684 18284
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 3700 18164 3752 18216
rect 3424 18096 3476 18148
rect 5356 18164 5408 18216
rect 5724 18207 5776 18216
rect 5724 18173 5733 18207
rect 5733 18173 5767 18207
rect 5767 18173 5776 18207
rect 5724 18164 5776 18173
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 6368 18164 6420 18216
rect 7748 18343 7800 18352
rect 7748 18309 7757 18343
rect 7757 18309 7791 18343
rect 7791 18309 7800 18343
rect 7748 18300 7800 18309
rect 8392 18232 8444 18284
rect 8300 18164 8352 18216
rect 8576 18232 8628 18284
rect 12808 18300 12860 18352
rect 13728 18368 13780 18420
rect 16672 18368 16724 18420
rect 21088 18368 21140 18420
rect 21180 18368 21232 18420
rect 9956 18232 10008 18284
rect 12072 18232 12124 18284
rect 4988 18096 5040 18148
rect 6644 18096 6696 18148
rect 7564 18096 7616 18148
rect 9128 18096 9180 18148
rect 6736 18028 6788 18080
rect 7288 18028 7340 18080
rect 8208 18028 8260 18080
rect 8300 18028 8352 18080
rect 9312 18028 9364 18080
rect 9496 18096 9548 18148
rect 11428 18164 11480 18216
rect 11796 18164 11848 18216
rect 12624 18232 12676 18284
rect 14556 18300 14608 18352
rect 15016 18300 15068 18352
rect 16028 18232 16080 18284
rect 16488 18275 16540 18284
rect 16488 18241 16497 18275
rect 16497 18241 16531 18275
rect 16531 18241 16540 18275
rect 16488 18232 16540 18241
rect 16672 18232 16724 18284
rect 20996 18300 21048 18352
rect 22836 18343 22888 18352
rect 22836 18309 22845 18343
rect 22845 18309 22879 18343
rect 22879 18309 22888 18343
rect 22836 18300 22888 18309
rect 19340 18232 19392 18284
rect 9864 18028 9916 18080
rect 10600 18028 10652 18080
rect 11888 18028 11940 18080
rect 12256 18096 12308 18148
rect 15108 18164 15160 18216
rect 15016 18139 15068 18148
rect 15016 18105 15025 18139
rect 15025 18105 15059 18139
rect 15059 18105 15068 18139
rect 15016 18096 15068 18105
rect 16948 18164 17000 18216
rect 17500 18207 17552 18216
rect 17500 18173 17509 18207
rect 17509 18173 17543 18207
rect 17543 18173 17552 18207
rect 17500 18164 17552 18173
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 20076 18207 20128 18216
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20996 18164 21048 18216
rect 21732 18232 21784 18284
rect 23388 18300 23440 18352
rect 23848 18300 23900 18352
rect 24768 18300 24820 18352
rect 26700 18368 26752 18420
rect 30104 18368 30156 18420
rect 30472 18368 30524 18420
rect 25320 18343 25372 18352
rect 25320 18309 25329 18343
rect 25329 18309 25363 18343
rect 25363 18309 25372 18343
rect 25320 18300 25372 18309
rect 26056 18343 26108 18352
rect 26056 18309 26065 18343
rect 26065 18309 26099 18343
rect 26099 18309 26108 18343
rect 26056 18300 26108 18309
rect 28632 18300 28684 18352
rect 29092 18300 29144 18352
rect 43352 18300 43404 18352
rect 27804 18232 27856 18284
rect 29644 18232 29696 18284
rect 19984 18096 20036 18148
rect 12716 18028 12768 18080
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 14556 18028 14608 18080
rect 15660 18028 15712 18080
rect 17868 18028 17920 18080
rect 18328 18028 18380 18080
rect 22836 18164 22888 18216
rect 26240 18164 26292 18216
rect 27068 18164 27120 18216
rect 30380 18096 30432 18148
rect 45008 18164 45060 18216
rect 39580 18096 39632 18148
rect 24676 18028 24728 18080
rect 26700 18071 26752 18080
rect 26700 18037 26709 18071
rect 26709 18037 26743 18071
rect 26743 18037 26752 18071
rect 26700 18028 26752 18037
rect 27344 18028 27396 18080
rect 29828 18071 29880 18080
rect 29828 18037 29837 18071
rect 29837 18037 29871 18071
rect 29871 18037 29880 18071
rect 29828 18028 29880 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 8392 17824 8444 17876
rect 8576 17824 8628 17876
rect 9404 17824 9456 17876
rect 10324 17824 10376 17876
rect 1860 17756 1912 17808
rect 6644 17799 6696 17808
rect 6644 17765 6653 17799
rect 6653 17765 6687 17799
rect 6687 17765 6696 17799
rect 6644 17756 6696 17765
rect 7104 17756 7156 17808
rect 7840 17799 7892 17808
rect 7840 17765 7849 17799
rect 7849 17765 7883 17799
rect 7883 17765 7892 17799
rect 7840 17756 7892 17765
rect 16120 17824 16172 17876
rect 9036 17688 9088 17740
rect 3608 17620 3660 17672
rect 3884 17620 3936 17672
rect 4160 17620 4212 17672
rect 4620 17620 4672 17672
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 1216 17552 1268 17604
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 3424 17527 3476 17536
rect 3424 17493 3433 17527
rect 3433 17493 3467 17527
rect 3467 17493 3476 17527
rect 3424 17484 3476 17493
rect 3792 17527 3844 17536
rect 3792 17493 3801 17527
rect 3801 17493 3835 17527
rect 3835 17493 3844 17527
rect 3792 17484 3844 17493
rect 6184 17552 6236 17604
rect 7288 17552 7340 17604
rect 8576 17552 8628 17604
rect 7472 17484 7524 17536
rect 7564 17484 7616 17536
rect 10876 17756 10928 17808
rect 11888 17756 11940 17808
rect 13636 17756 13688 17808
rect 15292 17756 15344 17808
rect 16764 17824 16816 17876
rect 17132 17824 17184 17876
rect 17684 17756 17736 17808
rect 9680 17688 9732 17740
rect 10140 17688 10192 17740
rect 14372 17688 14424 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 16948 17688 17000 17740
rect 17040 17688 17092 17740
rect 20076 17756 20128 17808
rect 21824 17756 21876 17808
rect 26240 17824 26292 17876
rect 27344 17867 27396 17876
rect 27344 17833 27368 17867
rect 27368 17833 27396 17867
rect 27344 17824 27396 17833
rect 27436 17824 27488 17876
rect 29000 17824 29052 17876
rect 29092 17867 29144 17876
rect 29092 17833 29101 17867
rect 29101 17833 29135 17867
rect 29135 17833 29144 17867
rect 29092 17824 29144 17833
rect 31944 17867 31996 17876
rect 31944 17833 31953 17867
rect 31953 17833 31987 17867
rect 31987 17833 31996 17867
rect 31944 17824 31996 17833
rect 24308 17756 24360 17808
rect 28448 17756 28500 17808
rect 20444 17688 20496 17740
rect 24492 17688 24544 17740
rect 24676 17688 24728 17740
rect 25780 17688 25832 17740
rect 27804 17688 27856 17740
rect 30196 17731 30248 17740
rect 30196 17697 30205 17731
rect 30205 17697 30239 17731
rect 30239 17697 30248 17731
rect 30196 17688 30248 17697
rect 30380 17756 30432 17808
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 13360 17620 13412 17672
rect 9404 17552 9456 17604
rect 10324 17484 10376 17536
rect 12164 17552 12216 17604
rect 12256 17595 12308 17604
rect 12256 17561 12265 17595
rect 12265 17561 12299 17595
rect 12299 17561 12308 17595
rect 12256 17552 12308 17561
rect 11336 17484 11388 17536
rect 11888 17484 11940 17536
rect 14924 17620 14976 17672
rect 15384 17620 15436 17672
rect 17684 17620 17736 17672
rect 20904 17620 20956 17672
rect 21732 17663 21784 17672
rect 21732 17629 21741 17663
rect 21741 17629 21775 17663
rect 21775 17629 21784 17663
rect 21732 17620 21784 17629
rect 22008 17620 22060 17672
rect 16304 17552 16356 17604
rect 14464 17527 14516 17536
rect 14464 17493 14473 17527
rect 14473 17493 14507 17527
rect 14507 17493 14516 17527
rect 14464 17484 14516 17493
rect 14924 17527 14976 17536
rect 14924 17493 14933 17527
rect 14933 17493 14967 17527
rect 14967 17493 14976 17527
rect 14924 17484 14976 17493
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 16396 17484 16448 17536
rect 18328 17484 18380 17536
rect 18696 17527 18748 17536
rect 18696 17493 18705 17527
rect 18705 17493 18739 17527
rect 18739 17493 18748 17527
rect 18696 17484 18748 17493
rect 18880 17552 18932 17604
rect 21272 17552 21324 17604
rect 23204 17552 23256 17604
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 21640 17484 21692 17536
rect 25412 17552 25464 17604
rect 26700 17552 26752 17604
rect 24400 17527 24452 17536
rect 24400 17493 24409 17527
rect 24409 17493 24443 17527
rect 24443 17493 24452 17527
rect 30748 17552 30800 17604
rect 24400 17484 24452 17493
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 31944 17620 31996 17672
rect 37556 17552 37608 17604
rect 28816 17484 28868 17493
rect 30932 17527 30984 17536
rect 30932 17493 30941 17527
rect 30941 17493 30975 17527
rect 30975 17493 30984 17527
rect 30932 17484 30984 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 4436 17255 4488 17264
rect 4436 17221 4445 17255
rect 4445 17221 4479 17255
rect 4479 17221 4488 17255
rect 4436 17212 4488 17221
rect 7380 17280 7432 17332
rect 8576 17280 8628 17332
rect 9588 17280 9640 17332
rect 10416 17280 10468 17332
rect 11612 17280 11664 17332
rect 1308 17076 1360 17128
rect 5356 17144 5408 17196
rect 6092 17144 6144 17196
rect 6460 17144 6512 17196
rect 7840 17144 7892 17196
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 5356 17008 5408 17060
rect 7932 17076 7984 17128
rect 8852 17076 8904 17128
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 9772 17076 9824 17128
rect 10324 17144 10376 17196
rect 10784 17187 10836 17196
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 10784 17144 10836 17153
rect 11336 17144 11388 17196
rect 12532 17144 12584 17196
rect 13084 17280 13136 17332
rect 13636 17280 13688 17332
rect 13728 17323 13780 17332
rect 13728 17289 13737 17323
rect 13737 17289 13771 17323
rect 13771 17289 13780 17323
rect 13728 17280 13780 17289
rect 18328 17212 18380 17264
rect 20076 17212 20128 17264
rect 13452 17144 13504 17196
rect 15292 17144 15344 17196
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 17132 17144 17184 17196
rect 17224 17187 17276 17196
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 20168 17144 20220 17196
rect 20904 17144 20956 17196
rect 10048 17119 10100 17128
rect 10048 17085 10057 17119
rect 10057 17085 10091 17119
rect 10091 17085 10100 17119
rect 10048 17076 10100 17085
rect 13084 17119 13136 17128
rect 13084 17085 13093 17119
rect 13093 17085 13127 17119
rect 13127 17085 13136 17119
rect 13084 17076 13136 17085
rect 13820 17076 13872 17128
rect 6460 17051 6512 17060
rect 6460 17017 6469 17051
rect 6469 17017 6503 17051
rect 6503 17017 6512 17051
rect 6460 17008 6512 17017
rect 6828 17051 6880 17060
rect 6828 17017 6837 17051
rect 6837 17017 6871 17051
rect 6871 17017 6880 17051
rect 6828 17008 6880 17017
rect 15476 17076 15528 17128
rect 15844 17076 15896 17128
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 9036 16940 9088 16992
rect 10232 16940 10284 16992
rect 10876 16940 10928 16992
rect 11704 16940 11756 16992
rect 12808 16940 12860 16992
rect 15752 16940 15804 16992
rect 16120 17051 16172 17060
rect 16120 17017 16129 17051
rect 16129 17017 16163 17051
rect 16163 17017 16172 17051
rect 16120 17008 16172 17017
rect 17040 17008 17092 17060
rect 19708 17076 19760 17128
rect 20628 17076 20680 17128
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 21456 17280 21508 17332
rect 24400 17280 24452 17332
rect 24768 17280 24820 17332
rect 21640 17212 21692 17264
rect 23296 17212 23348 17264
rect 24032 17212 24084 17264
rect 24308 17255 24360 17264
rect 24308 17221 24317 17255
rect 24317 17221 24351 17255
rect 24351 17221 24360 17255
rect 28816 17280 28868 17332
rect 29092 17280 29144 17332
rect 30196 17280 30248 17332
rect 37004 17280 37056 17332
rect 24308 17212 24360 17221
rect 26700 17212 26752 17264
rect 30748 17212 30800 17264
rect 22836 17144 22888 17196
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 27804 17187 27856 17196
rect 27804 17153 27813 17187
rect 27813 17153 27847 17187
rect 27847 17153 27856 17187
rect 27804 17144 27856 17153
rect 16764 16940 16816 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 17500 16940 17552 16992
rect 21272 17008 21324 17060
rect 21640 17076 21692 17128
rect 24492 17076 24544 17128
rect 27712 17076 27764 17128
rect 30380 17076 30432 17128
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 20812 16940 20864 16992
rect 22652 16940 22704 16992
rect 23296 16983 23348 16992
rect 23296 16949 23305 16983
rect 23305 16949 23339 16983
rect 23339 16949 23348 16983
rect 23296 16940 23348 16949
rect 24676 16940 24728 16992
rect 25136 16940 25188 16992
rect 26700 16983 26752 16992
rect 26700 16949 26709 16983
rect 26709 16949 26743 16983
rect 26743 16949 26752 16983
rect 26700 16940 26752 16949
rect 27160 16940 27212 16992
rect 42800 16940 42852 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 848 16736 900 16788
rect 1124 16736 1176 16788
rect 3608 16779 3660 16788
rect 3608 16745 3617 16779
rect 3617 16745 3651 16779
rect 3651 16745 3660 16779
rect 3608 16736 3660 16745
rect 3976 16736 4028 16788
rect 5356 16736 5408 16788
rect 5816 16736 5868 16788
rect 4252 16668 4304 16720
rect 7564 16736 7616 16788
rect 572 16600 624 16652
rect 848 16600 900 16652
rect 2228 16600 2280 16652
rect 5908 16600 5960 16652
rect 6000 16600 6052 16652
rect 8116 16736 8168 16788
rect 11612 16736 11664 16788
rect 12532 16779 12584 16788
rect 8116 16600 8168 16652
rect 8576 16668 8628 16720
rect 9496 16668 9548 16720
rect 9772 16668 9824 16720
rect 9864 16668 9916 16720
rect 10416 16600 10468 16652
rect 10876 16668 10928 16720
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 12348 16711 12400 16720
rect 12348 16677 12357 16711
rect 12357 16677 12391 16711
rect 12391 16677 12400 16711
rect 12348 16668 12400 16677
rect 1308 16464 1360 16516
rect 5080 16532 5132 16584
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 9772 16532 9824 16584
rect 11888 16643 11940 16652
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 7288 16464 7340 16516
rect 2596 16396 2648 16448
rect 6460 16396 6512 16448
rect 6828 16396 6880 16448
rect 6920 16396 6972 16448
rect 9036 16464 9088 16516
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 8208 16396 8260 16405
rect 9312 16464 9364 16516
rect 9864 16464 9916 16516
rect 12532 16532 12584 16584
rect 16212 16736 16264 16788
rect 16304 16736 16356 16788
rect 16764 16736 16816 16788
rect 19708 16736 19760 16788
rect 21180 16736 21232 16788
rect 30932 16736 30984 16788
rect 18328 16668 18380 16720
rect 22284 16668 22336 16720
rect 14464 16600 14516 16652
rect 16304 16600 16356 16652
rect 17224 16600 17276 16652
rect 20444 16600 20496 16652
rect 20720 16600 20772 16652
rect 25872 16668 25924 16720
rect 25964 16711 26016 16720
rect 25964 16677 25973 16711
rect 25973 16677 26007 16711
rect 26007 16677 26016 16711
rect 25964 16668 26016 16677
rect 22836 16600 22888 16652
rect 25136 16643 25188 16652
rect 25136 16609 25145 16643
rect 25145 16609 25179 16643
rect 25179 16609 25188 16643
rect 25136 16600 25188 16609
rect 25780 16600 25832 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27160 16643 27212 16652
rect 27160 16609 27169 16643
rect 27169 16609 27203 16643
rect 27203 16609 27212 16643
rect 27160 16600 27212 16609
rect 28816 16600 28868 16652
rect 31944 16600 31996 16652
rect 15292 16532 15344 16584
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 9588 16396 9640 16448
rect 9772 16439 9824 16448
rect 9772 16405 9781 16439
rect 9781 16405 9815 16439
rect 9815 16405 9824 16439
rect 9772 16396 9824 16405
rect 10508 16396 10560 16448
rect 11244 16439 11296 16448
rect 11244 16405 11253 16439
rect 11253 16405 11287 16439
rect 11287 16405 11296 16439
rect 11244 16396 11296 16405
rect 11704 16439 11756 16448
rect 11704 16405 11713 16439
rect 11713 16405 11747 16439
rect 11747 16405 11756 16439
rect 11704 16396 11756 16405
rect 11888 16464 11940 16516
rect 12348 16464 12400 16516
rect 12808 16464 12860 16516
rect 12164 16396 12216 16448
rect 16672 16464 16724 16516
rect 16948 16464 17000 16516
rect 17224 16464 17276 16516
rect 18328 16532 18380 16584
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 23296 16532 23348 16584
rect 24308 16532 24360 16584
rect 25044 16532 25096 16584
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 14832 16396 14884 16448
rect 15200 16396 15252 16448
rect 16120 16396 16172 16448
rect 16212 16439 16264 16448
rect 16212 16405 16221 16439
rect 16221 16405 16255 16439
rect 16255 16405 16264 16439
rect 16212 16396 16264 16405
rect 16764 16396 16816 16448
rect 19340 16464 19392 16516
rect 20168 16464 20220 16516
rect 21456 16507 21508 16516
rect 21456 16473 21465 16507
rect 21465 16473 21499 16507
rect 21499 16473 21508 16507
rect 21456 16464 21508 16473
rect 23848 16464 23900 16516
rect 24124 16464 24176 16516
rect 17684 16396 17736 16448
rect 18512 16396 18564 16448
rect 18604 16396 18656 16448
rect 20720 16396 20772 16448
rect 22468 16396 22520 16448
rect 23756 16396 23808 16448
rect 25044 16439 25096 16448
rect 25044 16405 25053 16439
rect 25053 16405 25087 16439
rect 25087 16405 25096 16439
rect 25044 16396 25096 16405
rect 25964 16396 26016 16448
rect 27712 16532 27764 16584
rect 28448 16464 28500 16516
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 7196 16192 7248 16244
rect 4344 16167 4396 16176
rect 4344 16133 4353 16167
rect 4353 16133 4387 16167
rect 4387 16133 4396 16167
rect 4344 16124 4396 16133
rect 1308 15988 1360 16040
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 6000 16056 6052 16108
rect 8852 16192 8904 16244
rect 9680 16192 9732 16244
rect 4712 15988 4764 16040
rect 5908 16031 5960 16040
rect 5908 15997 5917 16031
rect 5917 15997 5951 16031
rect 5951 15997 5960 16031
rect 5908 15988 5960 15997
rect 6552 15988 6604 16040
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 8392 16124 8444 16176
rect 11152 16192 11204 16244
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 12256 16192 12308 16244
rect 14740 16192 14792 16244
rect 10784 16124 10836 16176
rect 12532 16124 12584 16176
rect 16488 16124 16540 16176
rect 16948 16167 17000 16176
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 7932 16056 7984 16108
rect 8484 16099 8536 16108
rect 8484 16065 8493 16099
rect 8493 16065 8527 16099
rect 8527 16065 8536 16099
rect 8484 16056 8536 16065
rect 9864 16056 9916 16108
rect 6184 15920 6236 15972
rect 7472 15920 7524 15972
rect 8392 15988 8444 16040
rect 10140 16056 10192 16108
rect 10692 16056 10744 16108
rect 10876 16056 10928 16108
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 13360 16056 13412 16108
rect 14924 16056 14976 16108
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 13544 15988 13596 16040
rect 10968 15963 11020 15972
rect 10968 15929 10977 15963
rect 10977 15929 11011 15963
rect 11011 15929 11020 15963
rect 10968 15920 11020 15929
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 5816 15852 5868 15904
rect 7932 15852 7984 15904
rect 11428 15852 11480 15904
rect 12624 15852 12676 15904
rect 13636 15852 13688 15904
rect 14740 15852 14792 15904
rect 16396 16056 16448 16108
rect 16948 16133 16957 16167
rect 16957 16133 16991 16167
rect 16991 16133 17000 16167
rect 16948 16124 17000 16133
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 18604 16192 18656 16244
rect 18696 16192 18748 16244
rect 20812 16192 20864 16244
rect 21272 16235 21324 16244
rect 21272 16201 21281 16235
rect 21281 16201 21315 16235
rect 21315 16201 21324 16235
rect 21272 16192 21324 16201
rect 16672 16056 16724 16108
rect 17224 15988 17276 16040
rect 17316 15988 17368 16040
rect 19156 16056 19208 16108
rect 19708 16099 19760 16108
rect 19708 16065 19717 16099
rect 19717 16065 19751 16099
rect 19751 16065 19760 16099
rect 24952 16192 25004 16244
rect 25228 16124 25280 16176
rect 19708 16056 19760 16065
rect 22560 16056 22612 16108
rect 24308 16099 24360 16108
rect 24308 16065 24317 16099
rect 24317 16065 24351 16099
rect 24351 16065 24360 16099
rect 24308 16056 24360 16065
rect 24676 16056 24728 16108
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 26240 16056 26292 16108
rect 26700 16056 26752 16108
rect 15200 15852 15252 15904
rect 16212 15852 16264 15904
rect 17500 15920 17552 15972
rect 21272 15988 21324 16040
rect 21364 15988 21416 16040
rect 21916 15988 21968 16040
rect 23480 15988 23532 16040
rect 23848 15988 23900 16040
rect 24032 15988 24084 16040
rect 24768 15988 24820 16040
rect 27160 15988 27212 16040
rect 26148 15920 26200 15972
rect 29736 15920 29788 15972
rect 22652 15852 22704 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 2872 15648 2924 15700
rect 3976 15580 4028 15632
rect 1308 15512 1360 15564
rect 3700 15512 3752 15564
rect 5356 15580 5408 15632
rect 7840 15623 7892 15632
rect 7840 15589 7849 15623
rect 7849 15589 7883 15623
rect 7883 15589 7892 15623
rect 7840 15580 7892 15589
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 3424 15444 3476 15496
rect 5540 15512 5592 15564
rect 5816 15555 5868 15564
rect 5816 15521 5825 15555
rect 5825 15521 5859 15555
rect 5859 15521 5868 15555
rect 5816 15512 5868 15521
rect 6736 15512 6788 15564
rect 6920 15555 6972 15564
rect 6920 15521 6929 15555
rect 6929 15521 6963 15555
rect 6963 15521 6972 15555
rect 6920 15512 6972 15521
rect 8760 15648 8812 15700
rect 8392 15555 8444 15564
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 12808 15648 12860 15700
rect 10324 15580 10376 15632
rect 12072 15623 12124 15632
rect 12072 15589 12081 15623
rect 12081 15589 12115 15623
rect 12115 15589 12124 15623
rect 12072 15580 12124 15589
rect 12164 15580 12216 15632
rect 15844 15691 15896 15700
rect 15844 15657 15853 15691
rect 15853 15657 15887 15691
rect 15887 15657 15896 15691
rect 15844 15648 15896 15657
rect 19616 15648 19668 15700
rect 21916 15648 21968 15700
rect 23848 15648 23900 15700
rect 24676 15648 24728 15700
rect 10692 15512 10744 15564
rect 12900 15512 12952 15564
rect 13360 15512 13412 15564
rect 14096 15555 14148 15564
rect 14096 15521 14105 15555
rect 14105 15521 14139 15555
rect 14139 15521 14148 15555
rect 14096 15512 14148 15521
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 16120 15512 16172 15564
rect 5908 15444 5960 15496
rect 6644 15444 6696 15496
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 14740 15444 14792 15496
rect 16212 15444 16264 15496
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 5356 15308 5408 15360
rect 5816 15308 5868 15360
rect 6000 15308 6052 15360
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 6460 15308 6512 15360
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 7564 15308 7616 15360
rect 8484 15376 8536 15428
rect 11152 15376 11204 15428
rect 12256 15376 12308 15428
rect 9496 15308 9548 15360
rect 9864 15308 9916 15360
rect 9956 15351 10008 15360
rect 9956 15317 9965 15351
rect 9965 15317 9999 15351
rect 9999 15317 10008 15351
rect 9956 15308 10008 15317
rect 11612 15308 11664 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 13728 15308 13780 15360
rect 14188 15308 14240 15360
rect 14648 15308 14700 15360
rect 15476 15351 15528 15360
rect 15476 15317 15485 15351
rect 15485 15317 15519 15351
rect 15519 15317 15528 15351
rect 19432 15512 19484 15564
rect 20628 15512 20680 15564
rect 20996 15512 21048 15564
rect 26332 15580 26384 15632
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 20168 15444 20220 15496
rect 25780 15555 25832 15564
rect 25780 15521 25789 15555
rect 25789 15521 25823 15555
rect 25823 15521 25832 15555
rect 25780 15512 25832 15521
rect 22928 15444 22980 15496
rect 25596 15487 25648 15496
rect 25596 15453 25605 15487
rect 25605 15453 25639 15487
rect 25639 15453 25648 15487
rect 25596 15444 25648 15453
rect 26976 15444 27028 15496
rect 17316 15419 17368 15428
rect 17316 15385 17325 15419
rect 17325 15385 17359 15419
rect 17359 15385 17368 15419
rect 17316 15376 17368 15385
rect 17776 15376 17828 15428
rect 19984 15376 20036 15428
rect 15476 15308 15528 15317
rect 16396 15308 16448 15360
rect 17408 15308 17460 15360
rect 19156 15308 19208 15360
rect 21456 15308 21508 15360
rect 21916 15308 21968 15360
rect 23940 15419 23992 15428
rect 23940 15385 23949 15419
rect 23949 15385 23983 15419
rect 23983 15385 23992 15419
rect 23940 15376 23992 15385
rect 43444 15376 43496 15428
rect 23388 15308 23440 15360
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 26332 15308 26384 15360
rect 46204 15308 46256 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 572 15104 624 15156
rect 1124 15104 1176 15156
rect 3516 15147 3568 15156
rect 3516 15113 3525 15147
rect 3525 15113 3559 15147
rect 3559 15113 3568 15147
rect 3516 15104 3568 15113
rect 4712 15104 4764 15156
rect 7472 15104 7524 15156
rect 8484 15104 8536 15156
rect 9220 15104 9272 15156
rect 11244 15104 11296 15156
rect 12716 15104 12768 15156
rect 13268 15104 13320 15156
rect 15476 15104 15528 15156
rect 18420 15147 18472 15156
rect 18420 15113 18429 15147
rect 18429 15113 18463 15147
rect 18463 15113 18472 15147
rect 18420 15104 18472 15113
rect 22100 15104 22152 15156
rect 22928 15104 22980 15156
rect 23296 15104 23348 15156
rect 24952 15104 25004 15156
rect 6000 15036 6052 15088
rect 6276 15036 6328 15088
rect 1124 14900 1176 14952
rect 3516 14968 3568 15020
rect 3884 14968 3936 15020
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 6184 14968 6236 15020
rect 8392 15036 8444 15088
rect 9036 15036 9088 15088
rect 9772 15036 9824 15088
rect 10232 15036 10284 15088
rect 10784 15079 10836 15088
rect 10784 15045 10793 15079
rect 10793 15045 10827 15079
rect 10827 15045 10836 15079
rect 10784 15036 10836 15045
rect 10968 15036 11020 15088
rect 14740 15036 14792 15088
rect 14924 15036 14976 15088
rect 17776 15036 17828 15088
rect 18144 15036 18196 15088
rect 20720 15036 20772 15088
rect 22560 15036 22612 15088
rect 7288 14968 7340 15020
rect 6276 14900 6328 14952
rect 7196 14832 7248 14884
rect 7932 14943 7984 14952
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 8576 15011 8628 15020
rect 8576 14977 8585 15011
rect 8585 14977 8619 15011
rect 8619 14977 8628 15011
rect 8576 14968 8628 14977
rect 8852 14968 8904 15020
rect 8392 14832 8444 14884
rect 8484 14832 8536 14884
rect 4896 14764 4948 14816
rect 5080 14764 5132 14816
rect 6920 14764 6972 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 12624 14968 12676 15020
rect 12900 14968 12952 15020
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 14372 14968 14424 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 19524 14968 19576 15020
rect 9680 14832 9732 14884
rect 10784 14832 10836 14884
rect 13268 14900 13320 14952
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 10232 14764 10284 14816
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 10508 14764 10560 14816
rect 11060 14764 11112 14816
rect 12716 14764 12768 14816
rect 14280 14900 14332 14952
rect 16856 14900 16908 14952
rect 18972 14900 19024 14952
rect 20628 14968 20680 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 23388 14968 23440 15020
rect 23940 14968 23992 15020
rect 26240 14968 26292 15020
rect 13820 14764 13872 14816
rect 16764 14832 16816 14884
rect 16304 14807 16356 14816
rect 16304 14773 16313 14807
rect 16313 14773 16347 14807
rect 16347 14773 16356 14807
rect 16304 14764 16356 14773
rect 16396 14764 16448 14816
rect 17592 14764 17644 14816
rect 18972 14764 19024 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 19800 14832 19852 14884
rect 23572 14900 23624 14952
rect 21916 14832 21968 14884
rect 23664 14832 23716 14884
rect 24860 14832 24912 14884
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 3884 14560 3936 14612
rect 6460 14560 6512 14612
rect 6736 14560 6788 14612
rect 10968 14560 11020 14612
rect 1308 14424 1360 14476
rect 5080 14424 5132 14476
rect 6828 14492 6880 14544
rect 6184 14424 6236 14476
rect 7564 14424 7616 14476
rect 7840 14424 7892 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 5172 14356 5224 14408
rect 5448 14399 5500 14408
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 8392 14492 8444 14544
rect 13360 14560 13412 14612
rect 13544 14560 13596 14612
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 14924 14560 14976 14612
rect 18696 14560 18748 14612
rect 22376 14560 22428 14612
rect 26976 14603 27028 14612
rect 26976 14569 26985 14603
rect 26985 14569 27019 14603
rect 27019 14569 27028 14603
rect 26976 14560 27028 14569
rect 18144 14492 18196 14544
rect 21732 14535 21784 14544
rect 21732 14501 21741 14535
rect 21741 14501 21775 14535
rect 21775 14501 21784 14535
rect 21732 14492 21784 14501
rect 23664 14492 23716 14544
rect 25780 14492 25832 14544
rect 9680 14424 9732 14476
rect 9772 14424 9824 14476
rect 10048 14424 10100 14476
rect 10508 14424 10560 14476
rect 12624 14424 12676 14476
rect 12716 14424 12768 14476
rect 14556 14424 14608 14476
rect 16304 14424 16356 14476
rect 17132 14424 17184 14476
rect 17224 14424 17276 14476
rect 18328 14424 18380 14476
rect 19800 14424 19852 14476
rect 9312 14356 9364 14408
rect 10324 14356 10376 14408
rect 11060 14356 11112 14408
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 13360 14356 13412 14408
rect 14096 14356 14148 14408
rect 14280 14356 14332 14408
rect 3976 14220 4028 14272
rect 5356 14288 5408 14340
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 6000 14288 6052 14340
rect 5908 14220 5960 14272
rect 6460 14220 6512 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 8852 14220 8904 14272
rect 9404 14263 9456 14272
rect 9404 14229 9413 14263
rect 9413 14229 9447 14263
rect 9447 14229 9456 14263
rect 9404 14220 9456 14229
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 9772 14220 9824 14229
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 10968 14220 11020 14272
rect 15200 14288 15252 14340
rect 15476 14288 15528 14340
rect 14832 14220 14884 14272
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 17408 14288 17460 14340
rect 18144 14288 18196 14340
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 22008 14424 22060 14476
rect 23940 14424 23992 14476
rect 26608 14424 26660 14476
rect 21824 14288 21876 14340
rect 21916 14288 21968 14340
rect 23572 14288 23624 14340
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 20904 14220 20956 14272
rect 21640 14220 21692 14272
rect 22744 14220 22796 14272
rect 26976 14356 27028 14408
rect 24952 14331 25004 14340
rect 24952 14297 24961 14331
rect 24961 14297 24995 14331
rect 24995 14297 25004 14331
rect 24952 14288 25004 14297
rect 25136 14288 25188 14340
rect 26332 14288 26384 14340
rect 24584 14263 24636 14272
rect 24584 14229 24593 14263
rect 24593 14229 24627 14263
rect 24627 14229 24636 14263
rect 24584 14220 24636 14229
rect 25688 14220 25740 14272
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 4712 14016 4764 14068
rect 6368 14016 6420 14068
rect 2320 13948 2372 14000
rect 5356 13948 5408 14000
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 9220 14016 9272 14068
rect 11060 14016 11112 14068
rect 8576 13991 8628 14000
rect 8576 13957 8585 13991
rect 8585 13957 8619 13991
rect 8619 13957 8628 13991
rect 8576 13948 8628 13957
rect 9496 13948 9548 14000
rect 9864 13948 9916 14000
rect 11612 13991 11664 14000
rect 11612 13957 11621 13991
rect 11621 13957 11655 13991
rect 11655 13957 11664 13991
rect 11612 13948 11664 13957
rect 14464 14016 14516 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 17224 14016 17276 14068
rect 17316 14016 17368 14068
rect 18972 14016 19024 14068
rect 21180 14016 21232 14068
rect 25780 14016 25832 14068
rect 16672 13948 16724 14000
rect 1492 13880 1544 13932
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 1308 13812 1360 13864
rect 3884 13880 3936 13932
rect 5264 13880 5316 13932
rect 11888 13880 11940 13932
rect 12624 13880 12676 13932
rect 13176 13880 13228 13932
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 4804 13812 4856 13864
rect 6368 13855 6420 13864
rect 6368 13821 6377 13855
rect 6377 13821 6411 13855
rect 6411 13821 6420 13855
rect 6368 13812 6420 13821
rect 6736 13812 6788 13864
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 7932 13812 7984 13864
rect 2136 13676 2188 13728
rect 4620 13676 4672 13728
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 5908 13744 5960 13796
rect 6552 13787 6604 13796
rect 6552 13753 6561 13787
rect 6561 13753 6595 13787
rect 6595 13753 6604 13787
rect 6552 13744 6604 13753
rect 8576 13744 8628 13796
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 10784 13812 10836 13864
rect 12164 13812 12216 13864
rect 12900 13812 12952 13864
rect 12716 13744 12768 13796
rect 13636 13812 13688 13864
rect 6460 13676 6512 13728
rect 7196 13676 7248 13728
rect 13176 13676 13228 13728
rect 13636 13676 13688 13728
rect 14096 13880 14148 13932
rect 14556 13812 14608 13864
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 15568 13880 15620 13932
rect 17684 13948 17736 14000
rect 18144 13948 18196 14000
rect 19432 13948 19484 14000
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 14372 13744 14424 13796
rect 15292 13744 15344 13796
rect 15476 13744 15528 13796
rect 16120 13744 16172 13796
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17500 13812 17552 13864
rect 17868 13812 17920 13864
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 21640 13880 21692 13932
rect 21824 13923 21876 13932
rect 21824 13889 21833 13923
rect 21833 13889 21867 13923
rect 21867 13889 21876 13923
rect 21824 13880 21876 13889
rect 22376 13880 22428 13932
rect 17040 13676 17092 13728
rect 20352 13812 20404 13864
rect 20720 13744 20772 13796
rect 19156 13676 19208 13728
rect 20168 13676 20220 13728
rect 21824 13676 21876 13728
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 23388 13880 23440 13932
rect 24584 13948 24636 14000
rect 25136 13948 25188 14000
rect 25688 13948 25740 14000
rect 23848 13855 23900 13864
rect 23848 13821 23857 13855
rect 23857 13821 23891 13855
rect 23891 13821 23900 13855
rect 23848 13812 23900 13821
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 34980 13880 35032 13932
rect 25136 13812 25188 13864
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 3332 13472 3384 13524
rect 3792 13472 3844 13524
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 3516 13243 3568 13252
rect 3516 13209 3525 13243
rect 3525 13209 3559 13243
rect 3559 13209 3568 13243
rect 3516 13200 3568 13209
rect 4804 13472 4856 13524
rect 5172 13472 5224 13524
rect 5632 13472 5684 13524
rect 6000 13472 6052 13524
rect 9772 13472 9824 13524
rect 8392 13404 8444 13456
rect 8576 13404 8628 13456
rect 4160 13379 4212 13388
rect 4160 13345 4169 13379
rect 4169 13345 4203 13379
rect 4203 13345 4212 13379
rect 4160 13336 4212 13345
rect 5448 13336 5500 13388
rect 5816 13268 5868 13320
rect 6276 13268 6328 13320
rect 2412 13132 2464 13184
rect 7564 13336 7616 13388
rect 8300 13336 8352 13388
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 11152 13404 11204 13456
rect 12716 13472 12768 13524
rect 13636 13472 13688 13524
rect 15016 13472 15068 13524
rect 17500 13472 17552 13524
rect 18972 13472 19024 13524
rect 19156 13472 19208 13524
rect 22560 13472 22612 13524
rect 23296 13472 23348 13524
rect 11888 13404 11940 13456
rect 21640 13404 21692 13456
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 13268 13336 13320 13388
rect 15200 13336 15252 13388
rect 16396 13336 16448 13388
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 17132 13379 17184 13388
rect 17132 13345 17141 13379
rect 17141 13345 17175 13379
rect 17175 13345 17184 13379
rect 17132 13336 17184 13345
rect 17500 13336 17552 13388
rect 22192 13336 22244 13388
rect 23756 13404 23808 13456
rect 23848 13404 23900 13456
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23480 13336 23532 13345
rect 4252 13132 4304 13184
rect 7104 13200 7156 13252
rect 5080 13132 5132 13184
rect 5816 13132 5868 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 6828 13132 6880 13184
rect 7288 13200 7340 13252
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 7932 13132 7984 13184
rect 9036 13132 9088 13184
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 12348 13200 12400 13252
rect 13268 13200 13320 13252
rect 15292 13200 15344 13252
rect 17040 13200 17092 13252
rect 18144 13200 18196 13252
rect 14188 13132 14240 13184
rect 15844 13132 15896 13184
rect 19984 13268 20036 13320
rect 22376 13268 22428 13320
rect 23020 13268 23072 13320
rect 21088 13200 21140 13252
rect 20352 13132 20404 13184
rect 23112 13132 23164 13184
rect 23388 13200 23440 13252
rect 26884 13200 26936 13252
rect 25228 13132 25280 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 7196 12971 7248 12980
rect 1308 12860 1360 12912
rect 1768 12860 1820 12912
rect 2504 12792 2556 12844
rect 1124 12724 1176 12776
rect 1676 12724 1728 12776
rect 480 12656 532 12708
rect 7196 12937 7205 12971
rect 7205 12937 7239 12971
rect 7239 12937 7248 12971
rect 7196 12928 7248 12937
rect 10600 12928 10652 12980
rect 10968 12928 11020 12980
rect 4344 12860 4396 12912
rect 4436 12860 4488 12912
rect 4804 12860 4856 12912
rect 6460 12860 6512 12912
rect 7380 12860 7432 12912
rect 8760 12860 8812 12912
rect 10140 12860 10192 12912
rect 13636 12928 13688 12980
rect 13728 12971 13780 12980
rect 13728 12937 13737 12971
rect 13737 12937 13771 12971
rect 13771 12937 13780 12971
rect 13728 12928 13780 12937
rect 14004 12928 14056 12980
rect 14188 12971 14240 12980
rect 14188 12937 14197 12971
rect 14197 12937 14231 12971
rect 14231 12937 14240 12971
rect 14188 12928 14240 12937
rect 16028 12928 16080 12980
rect 12716 12860 12768 12912
rect 13176 12860 13228 12912
rect 13360 12860 13412 12912
rect 14280 12860 14332 12912
rect 16120 12903 16172 12912
rect 16120 12869 16129 12903
rect 16129 12869 16163 12903
rect 16163 12869 16172 12903
rect 16120 12860 16172 12869
rect 3976 12792 4028 12844
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 5172 12724 5224 12776
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 6276 12792 6328 12844
rect 6736 12792 6788 12844
rect 6828 12792 6880 12844
rect 5816 12724 5868 12776
rect 7564 12656 7616 12708
rect 1860 12588 1912 12640
rect 5448 12588 5500 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7380 12588 7432 12640
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 9588 12724 9640 12776
rect 10140 12724 10192 12776
rect 13084 12792 13136 12844
rect 14740 12792 14792 12844
rect 15108 12792 15160 12844
rect 18420 12860 18472 12912
rect 18880 12860 18932 12912
rect 19156 12928 19208 12980
rect 20904 12928 20956 12980
rect 21180 12928 21232 12980
rect 21272 12928 21324 12980
rect 21916 12928 21968 12980
rect 20076 12860 20128 12912
rect 17040 12792 17092 12844
rect 17960 12792 18012 12844
rect 22468 12860 22520 12912
rect 22836 12928 22888 12980
rect 23296 12928 23348 12980
rect 23480 12928 23532 12980
rect 23572 12860 23624 12912
rect 10232 12656 10284 12708
rect 12256 12656 12308 12708
rect 8760 12588 8812 12640
rect 9496 12588 9548 12640
rect 11336 12588 11388 12640
rect 12164 12588 12216 12640
rect 12900 12588 12952 12640
rect 15200 12724 15252 12776
rect 15292 12724 15344 12776
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 15476 12656 15528 12708
rect 17500 12656 17552 12708
rect 20076 12724 20128 12776
rect 21456 12724 21508 12776
rect 22192 12792 22244 12844
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 22652 12724 22704 12776
rect 23664 12724 23716 12776
rect 17868 12588 17920 12640
rect 19432 12588 19484 12640
rect 23664 12588 23716 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 2780 12384 2832 12436
rect 3976 12384 4028 12436
rect 4344 12384 4396 12436
rect 4804 12384 4856 12436
rect 6092 12384 6144 12436
rect 7564 12384 7616 12436
rect 7748 12384 7800 12436
rect 10876 12384 10928 12436
rect 11244 12384 11296 12436
rect 11612 12384 11664 12436
rect 12532 12384 12584 12436
rect 12716 12384 12768 12436
rect 13728 12384 13780 12436
rect 14188 12384 14240 12436
rect 14556 12384 14608 12436
rect 4988 12316 5040 12368
rect 7380 12316 7432 12368
rect 8024 12316 8076 12368
rect 9772 12316 9824 12368
rect 10968 12316 11020 12368
rect 13452 12316 13504 12368
rect 4160 12248 4212 12300
rect 7104 12248 7156 12300
rect 9312 12248 9364 12300
rect 10876 12248 10928 12300
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 11336 12248 11388 12300
rect 12164 12248 12216 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 4344 12180 4396 12232
rect 4804 12180 4856 12232
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 6736 12180 6788 12232
rect 7472 12180 7524 12232
rect 10416 12180 10468 12232
rect 13268 12180 13320 12232
rect 15292 12316 15344 12368
rect 15476 12316 15528 12368
rect 17960 12384 18012 12436
rect 19156 12384 19208 12436
rect 20720 12384 20772 12436
rect 19524 12316 19576 12368
rect 15844 12248 15896 12300
rect 16212 12248 16264 12300
rect 13728 12180 13780 12232
rect 14464 12180 14516 12232
rect 18788 12248 18840 12300
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 2596 12112 2648 12164
rect 2872 12112 2924 12164
rect 3976 12112 4028 12164
rect 5540 12112 5592 12164
rect 5724 12112 5776 12164
rect 9128 12155 9180 12164
rect 9128 12121 9137 12155
rect 9137 12121 9171 12155
rect 9171 12121 9180 12155
rect 9128 12112 9180 12121
rect 9312 12112 9364 12164
rect 11888 12112 11940 12164
rect 12900 12112 12952 12164
rect 6276 12044 6328 12096
rect 8300 12044 8352 12096
rect 8852 12044 8904 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 11704 12044 11756 12096
rect 11980 12044 12032 12096
rect 14556 12112 14608 12164
rect 14924 12044 14976 12096
rect 17408 12044 17460 12096
rect 18420 12044 18472 12096
rect 18696 12044 18748 12096
rect 18880 12044 18932 12096
rect 19248 12044 19300 12096
rect 20352 12155 20404 12164
rect 20352 12121 20361 12155
rect 20361 12121 20395 12155
rect 20395 12121 20404 12155
rect 20352 12112 20404 12121
rect 22192 12180 22244 12232
rect 23664 12180 23716 12232
rect 23940 12180 23992 12232
rect 21916 12112 21968 12164
rect 25044 12112 25096 12164
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 24676 12044 24728 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 1584 11840 1636 11892
rect 2964 11840 3016 11892
rect 3608 11840 3660 11892
rect 5448 11840 5500 11892
rect 1308 11772 1360 11824
rect 1124 11704 1176 11756
rect 1400 11704 1452 11756
rect 3424 11704 3476 11756
rect 2504 11636 2556 11688
rect 4620 11772 4672 11824
rect 6828 11772 6880 11824
rect 8116 11772 8168 11824
rect 9036 11772 9088 11824
rect 9496 11772 9548 11824
rect 10600 11772 10652 11824
rect 5264 11704 5316 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 9128 11704 9180 11756
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 8392 11636 8444 11688
rect 8852 11636 8904 11688
rect 9864 11636 9916 11688
rect 9588 11568 9640 11620
rect 2780 11500 2832 11552
rect 5540 11500 5592 11552
rect 5724 11500 5776 11552
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 9404 11500 9456 11552
rect 10508 11500 10560 11552
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 11244 11704 11296 11756
rect 12072 11704 12124 11756
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 17868 11840 17920 11892
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 18604 11883 18656 11892
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 13360 11772 13412 11824
rect 15292 11772 15344 11824
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 11796 11636 11848 11688
rect 15016 11636 15068 11688
rect 10876 11568 10928 11620
rect 12900 11568 12952 11620
rect 12256 11500 12308 11552
rect 17040 11636 17092 11688
rect 17408 11636 17460 11688
rect 19432 11704 19484 11756
rect 18420 11636 18472 11688
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 18788 11636 18840 11688
rect 32404 11840 32456 11892
rect 21916 11815 21968 11824
rect 21916 11781 21925 11815
rect 21925 11781 21959 11815
rect 21959 11781 21968 11815
rect 21916 11772 21968 11781
rect 22744 11772 22796 11824
rect 23940 11772 23992 11824
rect 24676 11772 24728 11824
rect 19708 11679 19760 11688
rect 19708 11645 19717 11679
rect 19717 11645 19751 11679
rect 19751 11645 19760 11679
rect 19708 11636 19760 11645
rect 19156 11568 19208 11620
rect 22192 11636 22244 11688
rect 24032 11636 24084 11688
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 16120 11500 16172 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 21640 11500 21692 11552
rect 25136 11636 25188 11688
rect 24676 11500 24728 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 1584 11296 1636 11348
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 4896 11296 4948 11348
rect 5724 11296 5776 11348
rect 6736 11296 6788 11348
rect 8116 11296 8168 11348
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 4160 11203 4212 11212
rect 4160 11169 4169 11203
rect 4169 11169 4203 11203
rect 4203 11169 4212 11203
rect 4160 11160 4212 11169
rect 5816 11160 5868 11212
rect 11336 11296 11388 11348
rect 12348 11296 12400 11348
rect 13360 11296 13412 11348
rect 7104 11228 7156 11280
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 7196 11160 7248 11212
rect 7840 11160 7892 11212
rect 8852 11228 8904 11280
rect 12808 11228 12860 11280
rect 14648 11296 14700 11348
rect 16212 11296 16264 11348
rect 18972 11296 19024 11348
rect 20996 11296 21048 11348
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 23296 11296 23348 11348
rect 24308 11228 24360 11280
rect 24676 11228 24728 11280
rect 9220 11160 9272 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 13360 11160 13412 11212
rect 14188 11160 14240 11212
rect 18696 11160 18748 11212
rect 26884 11160 26936 11212
rect 7472 11092 7524 11144
rect 8484 11092 8536 11144
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 9864 11092 9916 11144
rect 13728 11092 13780 11144
rect 14464 11092 14516 11144
rect 16120 11092 16172 11144
rect 16856 11092 16908 11144
rect 19248 11092 19300 11144
rect 9772 11024 9824 11076
rect 9956 10956 10008 11008
rect 10324 10999 10376 11008
rect 10324 10965 10333 10999
rect 10333 10965 10367 10999
rect 10367 10965 10376 10999
rect 10324 10956 10376 10965
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 10968 10956 11020 11008
rect 13820 10999 13872 11008
rect 13820 10965 13829 10999
rect 13829 10965 13863 10999
rect 13863 10965 13872 10999
rect 13820 10956 13872 10965
rect 15292 10956 15344 11008
rect 17316 11024 17368 11076
rect 17684 11024 17736 11076
rect 16764 10999 16816 11008
rect 16764 10965 16773 10999
rect 16773 10965 16807 10999
rect 16807 10965 16816 10999
rect 16764 10956 16816 10965
rect 18880 11024 18932 11076
rect 19708 11024 19760 11076
rect 31300 11092 31352 11144
rect 47584 11092 47636 11144
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 21916 11024 21968 11076
rect 27620 11024 27672 11076
rect 21364 10956 21416 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 2044 10684 2096 10736
rect 6276 10684 6328 10736
rect 8024 10684 8076 10736
rect 14740 10752 14792 10804
rect 15384 10752 15436 10804
rect 17040 10752 17092 10804
rect 11428 10684 11480 10736
rect 12072 10684 12124 10736
rect 13820 10684 13872 10736
rect 16948 10684 17000 10736
rect 664 10616 716 10668
rect 4252 10616 4304 10668
rect 5356 10616 5408 10668
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 8852 10616 8904 10668
rect 9404 10616 9456 10668
rect 9680 10616 9732 10668
rect 11888 10616 11940 10668
rect 3240 10548 3292 10600
rect 2872 10480 2924 10532
rect 6920 10548 6972 10600
rect 5264 10480 5316 10532
rect 4344 10412 4396 10464
rect 6276 10412 6328 10464
rect 6552 10412 6604 10464
rect 8116 10548 8168 10600
rect 8208 10548 8260 10600
rect 10692 10548 10744 10600
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 11244 10548 11296 10600
rect 12440 10548 12492 10600
rect 14924 10616 14976 10668
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 18880 10616 18932 10668
rect 15200 10548 15252 10600
rect 15660 10480 15712 10532
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 16304 10548 16356 10600
rect 7840 10412 7892 10464
rect 9864 10412 9916 10464
rect 11796 10412 11848 10464
rect 16488 10480 16540 10532
rect 21456 10752 21508 10804
rect 21916 10795 21968 10804
rect 21916 10761 21925 10795
rect 21925 10761 21959 10795
rect 21959 10761 21968 10795
rect 21916 10752 21968 10761
rect 21548 10684 21600 10736
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 22652 10548 22704 10600
rect 21364 10480 21416 10532
rect 20536 10412 20588 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 2596 10208 2648 10260
rect 3700 10208 3752 10260
rect 3608 10140 3660 10192
rect 6736 10140 6788 10192
rect 8300 10140 8352 10192
rect 8760 10140 8812 10192
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9680 10208 9732 10260
rect 10784 10208 10836 10260
rect 11704 10208 11756 10260
rect 14188 10208 14240 10260
rect 17224 10208 17276 10260
rect 19800 10208 19852 10260
rect 21548 10251 21600 10260
rect 21548 10217 21557 10251
rect 21557 10217 21591 10251
rect 21591 10217 21600 10251
rect 21548 10208 21600 10217
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 4068 10072 4120 10124
rect 4804 10072 4856 10124
rect 7840 10072 7892 10124
rect 8116 10072 8168 10124
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 5632 10004 5684 10056
rect 4712 9936 4764 9988
rect 6368 10004 6420 10056
rect 8852 10004 8904 10056
rect 9128 10004 9180 10056
rect 11980 10072 12032 10124
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 15200 10072 15252 10124
rect 16212 10072 16264 10124
rect 10968 10004 11020 10056
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 14464 10004 14516 10056
rect 16856 10004 16908 10056
rect 19708 10072 19760 10124
rect 20720 10004 20772 10056
rect 21548 10004 21600 10056
rect 2412 9868 2464 9920
rect 7104 9979 7156 9988
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 11060 9936 11112 9988
rect 11796 9936 11848 9988
rect 12808 9936 12860 9988
rect 8760 9868 8812 9920
rect 8852 9868 8904 9920
rect 11888 9868 11940 9920
rect 13820 9868 13872 9920
rect 17040 9936 17092 9988
rect 16764 9868 16816 9920
rect 18880 9936 18932 9988
rect 19248 9936 19300 9988
rect 21640 9979 21692 9988
rect 21640 9945 21649 9979
rect 21649 9945 21683 9979
rect 21683 9945 21692 9979
rect 21640 9936 21692 9945
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 2136 9664 2188 9716
rect 5632 9664 5684 9716
rect 6276 9664 6328 9716
rect 6736 9664 6788 9716
rect 1400 9639 1452 9648
rect 1400 9605 1409 9639
rect 1409 9605 1443 9639
rect 1443 9605 1452 9639
rect 1400 9596 1452 9605
rect 1676 9596 1728 9648
rect 1032 9528 1084 9580
rect 4068 9596 4120 9648
rect 5172 9528 5224 9580
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 12348 9664 12400 9716
rect 12808 9664 12860 9716
rect 9128 9596 9180 9648
rect 9956 9596 10008 9648
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14372 9596 14424 9648
rect 16212 9707 16264 9716
rect 16212 9673 16221 9707
rect 16221 9673 16255 9707
rect 16255 9673 16264 9707
rect 16212 9664 16264 9673
rect 24492 9664 24544 9716
rect 16764 9596 16816 9648
rect 17224 9596 17276 9648
rect 18880 9596 18932 9648
rect 24584 9596 24636 9648
rect 7380 9528 7432 9580
rect 9680 9528 9732 9580
rect 3976 9392 4028 9444
rect 7380 9392 7432 9444
rect 7840 9460 7892 9512
rect 8484 9460 8536 9512
rect 8760 9460 8812 9512
rect 11244 9460 11296 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 16764 9460 16816 9512
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 20628 9528 20680 9580
rect 23756 9528 23808 9580
rect 28172 9528 28224 9580
rect 7932 9392 7984 9444
rect 13360 9392 13412 9444
rect 3700 9324 3752 9376
rect 6276 9324 6328 9376
rect 7104 9324 7156 9376
rect 8760 9324 8812 9376
rect 14280 9392 14332 9444
rect 21180 9460 21232 9512
rect 23388 9460 23440 9512
rect 31300 9596 31352 9648
rect 14004 9324 14056 9376
rect 19064 9435 19116 9444
rect 19064 9401 19073 9435
rect 19073 9401 19107 9435
rect 19107 9401 19116 9435
rect 19064 9392 19116 9401
rect 16120 9324 16172 9376
rect 28356 9324 28408 9376
rect 31576 9324 31628 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 3424 9120 3476 9172
rect 4252 9120 4304 9172
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 9680 9120 9732 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 4528 9095 4580 9104
rect 4528 9061 4537 9095
rect 4537 9061 4571 9095
rect 4571 9061 4580 9095
rect 4528 9052 4580 9061
rect 1216 8984 1268 9036
rect 3792 8984 3844 9036
rect 1860 8916 1912 8968
rect 2320 8916 2372 8968
rect 4528 8916 4580 8968
rect 7932 9052 7984 9104
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 7564 8916 7616 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8484 9052 8536 9104
rect 9956 9052 10008 9104
rect 8760 8984 8812 9036
rect 9772 8984 9824 9036
rect 11520 9120 11572 9172
rect 14188 9120 14240 9172
rect 15936 9120 15988 9172
rect 15384 9095 15436 9104
rect 15384 9061 15393 9095
rect 15393 9061 15427 9095
rect 15427 9061 15436 9095
rect 15384 9052 15436 9061
rect 16488 9120 16540 9172
rect 16764 9120 16816 9172
rect 17408 9120 17460 9172
rect 14372 8984 14424 9036
rect 16856 8984 16908 9036
rect 10324 8916 10376 8968
rect 18880 9120 18932 9172
rect 19432 9120 19484 9172
rect 9128 8848 9180 8900
rect 10968 8848 11020 8900
rect 7288 8780 7340 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 9220 8780 9272 8832
rect 9680 8780 9732 8832
rect 12532 8780 12584 8832
rect 13912 8780 13964 8832
rect 15568 8780 15620 8832
rect 16212 8848 16264 8900
rect 17224 8780 17276 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 572 8576 624 8628
rect 756 8508 808 8560
rect 2780 8440 2832 8492
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3516 8440 3568 8492
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 4528 8440 4580 8492
rect 3700 8304 3752 8356
rect 5080 8551 5132 8560
rect 5080 8517 5089 8551
rect 5089 8517 5123 8551
rect 5123 8517 5132 8551
rect 5080 8508 5132 8517
rect 5356 8551 5408 8560
rect 5356 8517 5365 8551
rect 5365 8517 5399 8551
rect 5399 8517 5408 8551
rect 5356 8508 5408 8517
rect 8576 8576 8628 8628
rect 12440 8576 12492 8628
rect 12532 8619 12584 8628
rect 12532 8585 12541 8619
rect 12541 8585 12575 8619
rect 12575 8585 12584 8619
rect 12532 8576 12584 8585
rect 14924 8576 14976 8628
rect 16304 8576 16356 8628
rect 17224 8576 17276 8628
rect 32496 8576 32548 8628
rect 6920 8508 6972 8560
rect 7748 8440 7800 8492
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 8116 8440 8168 8492
rect 8576 8440 8628 8492
rect 11428 8508 11480 8560
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 5356 8372 5408 8424
rect 5264 8304 5316 8356
rect 7012 8372 7064 8424
rect 8484 8304 8536 8356
rect 8760 8372 8812 8424
rect 9036 8372 9088 8424
rect 9220 8372 9272 8424
rect 10324 8372 10376 8424
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 14740 8508 14792 8560
rect 15384 8508 15436 8560
rect 16120 8508 16172 8560
rect 17316 8508 17368 8560
rect 11612 8483 11664 8492
rect 11612 8449 11621 8483
rect 11621 8449 11655 8483
rect 11655 8449 11664 8483
rect 11612 8440 11664 8449
rect 9864 8347 9916 8356
rect 9864 8313 9873 8347
rect 9873 8313 9907 8347
rect 9907 8313 9916 8347
rect 9864 8304 9916 8313
rect 12716 8440 12768 8492
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 13912 8304 13964 8356
rect 3516 8236 3568 8288
rect 3792 8236 3844 8288
rect 5908 8236 5960 8288
rect 6460 8236 6512 8288
rect 9220 8236 9272 8288
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 17132 8440 17184 8492
rect 16120 8372 16172 8424
rect 20352 8372 20404 8424
rect 20444 8304 20496 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 3700 8032 3752 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 5356 8075 5408 8084
rect 5356 8041 5365 8075
rect 5365 8041 5399 8075
rect 5399 8041 5408 8075
rect 5356 8032 5408 8041
rect 6368 8075 6420 8084
rect 6368 8041 6377 8075
rect 6377 8041 6411 8075
rect 6411 8041 6420 8075
rect 6368 8032 6420 8041
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 8300 8032 8352 8084
rect 9772 8032 9824 8084
rect 12072 8032 12124 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 14004 8032 14056 8084
rect 14188 8075 14240 8084
rect 14188 8041 14197 8075
rect 14197 8041 14231 8075
rect 14231 8041 14240 8075
rect 14188 8032 14240 8041
rect 19248 8032 19300 8084
rect 848 7964 900 8016
rect 5724 8007 5776 8016
rect 5724 7973 5733 8007
rect 5733 7973 5767 8007
rect 5767 7973 5776 8007
rect 5724 7964 5776 7973
rect 6644 7964 6696 8016
rect 1492 7896 1544 7948
rect 3792 7896 3844 7948
rect 7380 7896 7432 7948
rect 8116 7896 8168 7948
rect 9220 7896 9272 7948
rect 9956 7896 10008 7948
rect 10876 7896 10928 7948
rect 12440 7896 12492 7948
rect 2504 7828 2556 7880
rect 3608 7828 3660 7880
rect 940 7760 992 7812
rect 4252 7828 4304 7880
rect 7472 7828 7524 7880
rect 2964 7692 3016 7744
rect 5724 7760 5776 7812
rect 6828 7760 6880 7812
rect 11152 7828 11204 7880
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 15200 8007 15252 8016
rect 15200 7973 15209 8007
rect 15209 7973 15243 8007
rect 15243 7973 15252 8007
rect 15200 7964 15252 7973
rect 14188 7896 14240 7948
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 9772 7692 9824 7744
rect 13544 7760 13596 7812
rect 14740 7692 14792 7744
rect 22836 7692 22888 7744
rect 23388 7692 23440 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 3332 7488 3384 7540
rect 3608 7531 3660 7540
rect 3608 7497 3617 7531
rect 3617 7497 3651 7531
rect 3651 7497 3660 7531
rect 3608 7488 3660 7497
rect 1308 7420 1360 7472
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 2228 7352 2280 7404
rect 2964 7420 3016 7472
rect 4436 7488 4488 7540
rect 7656 7488 7708 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 10968 7488 11020 7540
rect 13544 7488 13596 7540
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 27620 7488 27672 7540
rect 3332 7352 3384 7404
rect 5540 7420 5592 7472
rect 4252 7352 4304 7404
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 8944 7352 8996 7404
rect 12072 7420 12124 7472
rect 15016 7420 15068 7472
rect 24308 7463 24360 7472
rect 24308 7429 24317 7463
rect 24317 7429 24351 7463
rect 24351 7429 24360 7463
rect 24308 7420 24360 7429
rect 11336 7352 11388 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 6460 7284 6512 7336
rect 11520 7284 11572 7336
rect 22468 7327 22520 7336
rect 22468 7293 22477 7327
rect 22477 7293 22511 7327
rect 22511 7293 22520 7327
rect 22468 7284 22520 7293
rect 2872 7216 2924 7268
rect 3976 7259 4028 7268
rect 3976 7225 3985 7259
rect 3985 7225 4019 7259
rect 4019 7225 4028 7259
rect 3976 7216 4028 7225
rect 12440 7148 12492 7200
rect 14004 7148 14056 7200
rect 17500 7148 17552 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 1584 6944 1636 6996
rect 2688 6944 2740 6996
rect 5172 6944 5224 6996
rect 23940 6944 23992 6996
rect 756 6808 808 6860
rect 3884 6876 3936 6928
rect 3148 6740 3200 6792
rect 3792 6808 3844 6860
rect 23756 6919 23808 6928
rect 23756 6885 23765 6919
rect 23765 6885 23799 6919
rect 23799 6885 23808 6919
rect 23756 6876 23808 6885
rect 8852 6808 8904 6860
rect 10508 6808 10560 6860
rect 3976 6740 4028 6792
rect 4068 6740 4120 6792
rect 21732 6740 21784 6792
rect 4344 6672 4396 6724
rect 3516 6604 3568 6656
rect 3976 6604 4028 6656
rect 23388 6647 23440 6656
rect 23388 6613 23397 6647
rect 23397 6613 23431 6647
rect 23431 6613 23440 6647
rect 23388 6604 23440 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 3332 6400 3384 6452
rect 22836 6443 22888 6452
rect 22836 6409 22845 6443
rect 22845 6409 22879 6443
rect 22879 6409 22888 6443
rect 22836 6400 22888 6409
rect 12164 6332 12216 6384
rect 2780 6264 2832 6316
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 1308 6196 1360 6248
rect 2872 6196 2924 6248
rect 24860 6196 24912 6248
rect 6092 6128 6144 6180
rect 19340 6128 19392 6180
rect 38752 6128 38804 6180
rect 4068 6060 4120 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 2780 5856 2832 5908
rect 3884 5856 3936 5908
rect 22468 5856 22520 5908
rect 9312 5788 9364 5840
rect 9588 5788 9640 5840
rect 12624 5788 12676 5840
rect 1216 5720 1268 5772
rect 1308 5652 1360 5704
rect 3608 5720 3660 5772
rect 14004 5720 14056 5772
rect 16856 5720 16908 5772
rect 2780 5652 2832 5704
rect 12624 5652 12676 5704
rect 19432 5788 19484 5840
rect 21732 5831 21784 5840
rect 21732 5797 21741 5831
rect 21741 5797 21775 5831
rect 21775 5797 21784 5831
rect 21732 5788 21784 5797
rect 2964 5584 3016 5636
rect 17040 5516 17092 5568
rect 20260 5652 20312 5704
rect 30288 5720 30340 5772
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 22192 5584 22244 5636
rect 23388 5584 23440 5636
rect 21364 5559 21416 5568
rect 21364 5525 21373 5559
rect 21373 5525 21407 5559
rect 21407 5525 21416 5559
rect 21364 5516 21416 5525
rect 24860 5627 24912 5636
rect 24860 5593 24869 5627
rect 24869 5593 24903 5627
rect 24903 5593 24912 5627
rect 24860 5584 24912 5593
rect 25780 5627 25832 5636
rect 25780 5593 25789 5627
rect 25789 5593 25823 5627
rect 25823 5593 25832 5627
rect 25780 5584 25832 5593
rect 27160 5627 27212 5636
rect 27160 5593 27169 5627
rect 27169 5593 27203 5627
rect 27203 5593 27212 5627
rect 27160 5584 27212 5593
rect 35716 5584 35768 5636
rect 25504 5516 25556 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 2964 5312 3016 5364
rect 27160 5312 27212 5364
rect 28816 5287 28868 5296
rect 28816 5253 28825 5287
rect 28825 5253 28859 5287
rect 28859 5253 28868 5287
rect 28816 5244 28868 5253
rect 1308 5176 1360 5228
rect 8392 5176 8444 5228
rect 12440 5176 12492 5228
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 15476 5108 15528 5160
rect 21364 5176 21416 5228
rect 22192 5219 22244 5228
rect 22192 5185 22210 5219
rect 22210 5185 22244 5219
rect 22192 5176 22244 5185
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 29644 5108 29696 5160
rect 31392 5108 31444 5160
rect 1860 4972 1912 5024
rect 17868 4972 17920 5024
rect 20536 4972 20588 5024
rect 22744 4972 22796 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 6828 4768 6880 4820
rect 17408 4768 17460 4820
rect 20260 4811 20312 4820
rect 20260 4777 20269 4811
rect 20269 4777 20303 4811
rect 20303 4777 20312 4811
rect 20260 4768 20312 4777
rect 28816 4768 28868 4820
rect 1308 4632 1360 4684
rect 10048 4632 10100 4684
rect 27528 4632 27580 4684
rect 2872 4564 2924 4616
rect 20260 4564 20312 4616
rect 17684 4428 17736 4480
rect 22744 4496 22796 4548
rect 37464 4496 37516 4548
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1400 4267 1452 4276
rect 1400 4233 1409 4267
rect 1409 4233 1443 4267
rect 1443 4233 1452 4267
rect 1400 4224 1452 4233
rect 1400 4088 1452 4140
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 4160 4088 4212 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 9680 3952 9732 4004
rect 3332 3884 3384 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 10600 3680 10652 3732
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 13452 3612 13504 3664
rect 31944 3612 31996 3664
rect 1308 3544 1360 3596
rect 25780 3544 25832 3596
rect 664 3476 716 3528
rect 2872 3476 2924 3528
rect 4068 3476 4120 3528
rect 12072 3476 12124 3528
rect 35716 3519 35768 3528
rect 35716 3485 35725 3519
rect 35725 3485 35759 3519
rect 35759 3485 35768 3519
rect 35716 3476 35768 3485
rect 32128 3408 32180 3460
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 31760 3340 31812 3392
rect 33600 3340 33652 3392
rect 49424 3408 49476 3460
rect 44088 3340 44140 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 9772 3136 9824 3188
rect 25504 3179 25556 3188
rect 25504 3145 25513 3179
rect 25513 3145 25547 3179
rect 25547 3145 25556 3179
rect 25504 3136 25556 3145
rect 27528 3136 27580 3188
rect 29644 3136 29696 3188
rect 33600 3136 33652 3188
rect 1308 3000 1360 3052
rect 2780 3000 2832 3052
rect 3332 3000 3384 3052
rect 10324 3068 10376 3120
rect 12624 3111 12676 3120
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 15476 3068 15528 3120
rect 17684 3068 17736 3120
rect 31392 3068 31444 3120
rect 7840 3000 7892 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17868 3000 17920 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 26240 3000 26292 3052
rect 28356 3043 28408 3052
rect 28356 3009 28365 3043
rect 28365 3009 28399 3043
rect 28399 3009 28408 3043
rect 28356 3000 28408 3009
rect 31024 3043 31076 3052
rect 31024 3009 31033 3043
rect 31033 3009 31067 3043
rect 31067 3009 31076 3043
rect 31024 3000 31076 3009
rect 33692 3043 33744 3052
rect 33692 3009 33701 3043
rect 33701 3009 33735 3043
rect 33735 3009 33744 3043
rect 33692 3000 33744 3009
rect 37464 3043 37516 3052
rect 37464 3009 37473 3043
rect 37473 3009 37507 3043
rect 37507 3009 37516 3043
rect 37464 3000 37516 3009
rect 5632 2932 5684 2984
rect 17408 2932 17460 2984
rect 35164 2932 35216 2984
rect 8300 2796 8352 2848
rect 12440 2864 12492 2916
rect 30288 2864 30340 2916
rect 46756 2932 46808 2984
rect 41420 2864 41472 2916
rect 17500 2796 17552 2848
rect 20076 2796 20128 2848
rect 21916 2796 21968 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 9588 2592 9640 2644
rect 26240 2635 26292 2644
rect 26240 2601 26249 2635
rect 26249 2601 26283 2635
rect 26283 2601 26292 2635
rect 26240 2592 26292 2601
rect 28356 2592 28408 2644
rect 31024 2592 31076 2644
rect 33692 2592 33744 2644
rect 2780 2524 2832 2576
rect 1216 2456 1268 2508
rect 4068 2456 4120 2508
rect 11612 2524 11664 2576
rect 6736 2456 6788 2508
rect 9404 2456 9456 2508
rect 12072 2456 12124 2508
rect 14740 2456 14792 2508
rect 17408 2456 17460 2508
rect 20168 2456 20220 2508
rect 22744 2456 22796 2508
rect 31576 2456 31628 2508
rect 1308 2320 1360 2372
rect 8300 2388 8352 2440
rect 9772 2388 9824 2440
rect 12440 2388 12492 2440
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 21916 2388 21968 2440
rect 6000 2252 6052 2304
rect 25412 2252 25464 2304
rect 27804 2252 27856 2304
rect 36084 2431 36136 2440
rect 36084 2397 36093 2431
rect 36093 2397 36127 2431
rect 36127 2397 36136 2431
rect 36084 2388 36136 2397
rect 30748 2252 30800 2304
rect 33416 2252 33468 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 2226 26200 2282 27000
rect 2870 26330 2926 27000
rect 2870 26302 3464 26330
rect 2870 26200 2926 26302
rect 572 24336 624 24342
rect 572 24278 624 24284
rect 584 16658 612 24278
rect 1032 24200 1084 24206
rect 1032 24142 1084 24148
rect 664 24132 716 24138
rect 664 24074 716 24080
rect 572 16652 624 16658
rect 572 16594 624 16600
rect 572 15156 624 15162
rect 572 15098 624 15104
rect 480 12708 532 12714
rect 480 12650 532 12656
rect 492 6914 520 12650
rect 584 8634 612 15098
rect 676 10674 704 24074
rect 756 23724 808 23730
rect 756 23666 808 23672
rect 664 10668 716 10674
rect 664 10610 716 10616
rect 572 8628 624 8634
rect 572 8570 624 8576
rect 768 8566 796 23666
rect 848 23588 900 23594
rect 848 23530 900 23536
rect 860 16794 888 23530
rect 940 20392 992 20398
rect 940 20334 992 20340
rect 848 16788 900 16794
rect 848 16730 900 16736
rect 848 16652 900 16658
rect 848 16594 900 16600
rect 756 8560 808 8566
rect 756 8502 808 8508
rect 492 6886 704 6914
rect 676 3534 704 6886
rect 768 6866 796 8502
rect 860 8022 888 16594
rect 848 8016 900 8022
rect 848 7958 900 7964
rect 952 7818 980 20334
rect 1044 9586 1072 24142
rect 1584 23520 1636 23526
rect 1584 23462 1636 23468
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1124 21480 1176 21486
rect 1124 21422 1176 21428
rect 1136 16946 1164 21422
rect 1320 20777 1348 22034
rect 1596 21457 1624 23462
rect 1582 21448 1638 21457
rect 1582 21383 1638 21392
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1780 20466 1808 23462
rect 2240 22234 2268 26200
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2778 24440 2834 24449
rect 2950 24443 3258 24452
rect 2778 24375 2780 24384
rect 2832 24375 2834 24384
rect 2780 24346 2832 24352
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 22250 2820 22986
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 1952 21480 2004 21486
rect 1952 21422 2004 21428
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1766 18864 1822 18873
rect 1400 18828 1452 18834
rect 1766 18799 1822 18808
rect 1400 18770 1452 18776
rect 1412 17921 1440 18770
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 1216 17604 1268 17610
rect 1216 17546 1268 17552
rect 1228 17105 1256 17546
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1136 16918 1256 16946
rect 1124 16788 1176 16794
rect 1124 16730 1176 16736
rect 1136 15162 1164 16730
rect 1124 15156 1176 15162
rect 1124 15098 1176 15104
rect 1122 15056 1178 15065
rect 1122 14991 1178 15000
rect 1136 14958 1164 14991
rect 1124 14952 1176 14958
rect 1124 14894 1176 14900
rect 1122 13424 1178 13433
rect 1122 13359 1178 13368
rect 1136 12782 1164 13359
rect 1124 12776 1176 12782
rect 1124 12718 1176 12724
rect 1122 12200 1178 12209
rect 1122 12135 1178 12144
rect 1136 11762 1164 12135
rect 1124 11756 1176 11762
rect 1124 11698 1176 11704
rect 1032 9580 1084 9586
rect 1032 9522 1084 9528
rect 1228 9042 1256 16918
rect 1320 16697 1348 17070
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1780 14414 1808 18799
rect 1872 17814 1900 20878
rect 1964 19961 1992 21422
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3344 21350 3372 22510
rect 3436 22166 3464 26302
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 3528 24274 3556 26200
rect 3882 25664 3938 25673
rect 3882 25599 3938 25608
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3606 23352 3662 23361
rect 3712 23322 3740 24006
rect 3790 23624 3846 23633
rect 3790 23559 3846 23568
rect 3804 23526 3832 23559
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3606 23287 3608 23296
rect 3660 23287 3662 23296
rect 3700 23316 3752 23322
rect 3608 23258 3660 23264
rect 3700 23258 3752 23264
rect 3514 23216 3570 23225
rect 3514 23151 3570 23160
rect 3424 22160 3476 22166
rect 3424 22102 3476 22108
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 3436 21146 3464 21626
rect 3424 21140 3476 21146
rect 2778 21111 2834 21120
rect 3424 21082 3476 21088
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 1950 19952 2006 19961
rect 1950 19887 2006 19896
rect 2056 19145 2084 20334
rect 2792 19553 2820 20810
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2778 19544 2834 19553
rect 2778 19479 2834 19488
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2042 19136 2098 19145
rect 2042 19071 2098 19080
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 2056 17513 2084 18158
rect 2042 17504 2098 17513
rect 2042 17439 2098 17448
rect 2516 17377 2544 18566
rect 2502 17368 2558 17377
rect 2502 17303 2558 17312
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 1766 13968 1822 13977
rect 1492 13932 1544 13938
rect 1766 13903 1768 13912
rect 1492 13874 1544 13880
rect 1820 13903 1822 13912
rect 1768 13874 1820 13880
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 12918 1348 12951
rect 1308 12912 1360 12918
rect 1308 12854 1360 12860
rect 1308 11824 1360 11830
rect 1306 11792 1308 11801
rect 1360 11792 1362 11801
rect 1306 11727 1362 11736
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 9654 1440 11698
rect 1504 11506 1532 13874
rect 2042 13832 2098 13841
rect 2042 13767 2098 13776
rect 1950 13424 2006 13433
rect 2056 13394 2084 13767
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 1950 13359 2006 13368
rect 2044 13388 2096 13394
rect 1768 13320 1820 13326
rect 1766 13288 1768 13297
rect 1820 13288 1822 13297
rect 1766 13223 1822 13232
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11898 1624 12174
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1504 11478 1624 11506
rect 1490 11384 1546 11393
rect 1596 11354 1624 11478
rect 1490 11319 1546 11328
rect 1584 11348 1636 11354
rect 1400 9648 1452 9654
rect 1400 9590 1452 9596
rect 1216 9036 1268 9042
rect 1216 8978 1268 8984
rect 1306 8120 1362 8129
rect 1306 8055 1362 8064
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 1320 7478 1348 8055
rect 1504 7954 1532 11319
rect 1584 11290 1636 11296
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1308 7472 1360 7478
rect 1308 7414 1360 7420
rect 1596 7410 1624 10911
rect 1688 9654 1716 12718
rect 1780 10810 1808 12854
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1872 8974 1900 12582
rect 1964 11218 1992 13359
rect 2044 13330 2096 13336
rect 2042 13288 2098 13297
rect 2042 13223 2098 13232
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 2056 10742 2084 13223
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 2148 10062 2176 13670
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9722 2176 9998
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 2240 7410 2268 16594
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2332 8974 2360 13942
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 9926 2452 13126
rect 2516 12850 2544 17303
rect 2700 17184 2728 19178
rect 2792 18329 2820 19314
rect 2884 18737 2912 19722
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2870 18728 2926 18737
rect 2870 18663 2926 18672
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2700 17156 2820 17184
rect 2686 17096 2742 17105
rect 2686 17031 2742 17040
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2608 12170 2636 16390
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2516 7886 2544 11630
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2608 10266 2636 11086
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2594 10160 2650 10169
rect 2594 10095 2596 10104
rect 2648 10095 2650 10104
rect 2596 10066 2648 10072
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 1596 7002 1624 7346
rect 2700 7002 2728 17031
rect 2792 12442 2820 17156
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2884 12288 2912 15642
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 3344 13954 3372 20878
rect 3436 20058 3464 21082
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3528 19786 3556 23151
rect 3712 23066 3740 23258
rect 3620 23038 3740 23066
rect 3620 21690 3648 23038
rect 3698 22808 3754 22817
rect 3698 22743 3754 22752
rect 3712 22506 3740 22743
rect 3792 22636 3844 22642
rect 3792 22578 3844 22584
rect 3700 22500 3752 22506
rect 3700 22442 3752 22448
rect 3804 22409 3832 22578
rect 3790 22400 3846 22409
rect 3790 22335 3846 22344
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 18154 3464 19654
rect 3620 19281 3648 21286
rect 3606 19272 3662 19281
rect 3606 19207 3662 19216
rect 3620 18737 3648 19207
rect 3606 18728 3662 18737
rect 3606 18663 3662 18672
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3620 17678 3648 18566
rect 3712 18222 3740 22170
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3804 21593 3832 21966
rect 3790 21584 3846 21593
rect 3790 21519 3846 21528
rect 3896 20482 3924 25599
rect 4066 25256 4122 25265
rect 4066 25191 4122 25200
rect 4080 25090 4108 25191
rect 4068 25084 4120 25090
rect 4068 25026 4120 25032
rect 4066 24848 4122 24857
rect 4066 24783 4068 24792
rect 4120 24783 4122 24792
rect 4068 24754 4120 24760
rect 4066 24032 4122 24041
rect 4066 23967 4122 23976
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 4080 23610 4108 23967
rect 4172 23798 4200 26200
rect 4804 25560 4856 25566
rect 4804 25502 4856 25508
rect 4252 24744 4304 24750
rect 4252 24686 4304 24692
rect 4264 24206 4292 24686
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4816 23730 4844 25502
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 3804 20454 3924 20482
rect 3804 19145 3832 20454
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 19802 3924 20198
rect 3988 20074 4016 23598
rect 4080 23582 4476 23610
rect 4066 23216 4122 23225
rect 4066 23151 4068 23160
rect 4120 23151 4122 23160
rect 4068 23122 4120 23128
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4172 22681 4200 22918
rect 4158 22672 4214 22681
rect 4158 22607 4214 22616
rect 4066 22536 4122 22545
rect 4122 22494 4292 22522
rect 4066 22471 4122 22480
rect 4160 22160 4212 22166
rect 4160 22102 4212 22108
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4080 22001 4108 22034
rect 4066 21992 4122 22001
rect 4066 21927 4122 21936
rect 4172 21486 4200 22102
rect 4264 22094 4292 22494
rect 4264 22066 4384 22094
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4264 21690 4292 21966
rect 4252 21684 4304 21690
rect 4252 21626 4304 21632
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4068 21072 4120 21078
rect 4068 21014 4120 21020
rect 4250 21040 4306 21049
rect 4080 20262 4108 21014
rect 4250 20975 4252 20984
rect 4304 20975 4306 20984
rect 4252 20946 4304 20952
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 3988 20046 4108 20074
rect 3896 19774 4016 19802
rect 3884 19712 3936 19718
rect 3882 19680 3884 19689
rect 3936 19680 3938 19689
rect 3882 19615 3938 19624
rect 3790 19136 3846 19145
rect 3790 19071 3846 19080
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3790 17912 3846 17921
rect 3790 17847 3846 17856
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3804 17542 3832 17847
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3436 17241 3464 17478
rect 3422 17232 3478 17241
rect 3422 17167 3478 17176
rect 3606 16824 3662 16833
rect 3606 16759 3608 16768
rect 3660 16759 3662 16768
rect 3608 16730 3660 16736
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3436 14074 3464 15438
rect 3528 15162 3556 16050
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3344 13926 3464 13954
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2884 12260 3004 12288
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 8498 2820 11494
rect 2884 10538 2912 12106
rect 2976 11898 3004 12260
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3238 10704 3294 10713
rect 3238 10639 3294 10648
rect 3252 10606 3280 10639
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2870 9752 2926 9761
rect 2870 9687 2926 9696
rect 2884 8498 2912 9687
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2778 7304 2834 7313
rect 2884 7274 2912 8434
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7478 3004 7686
rect 3344 7546 3372 13466
rect 3436 11937 3464 13926
rect 3528 13841 3556 14962
rect 3514 13832 3570 13841
rect 3514 13767 3570 13776
rect 3712 13716 3740 15506
rect 3528 13688 3740 13716
rect 3528 13258 3556 13688
rect 3698 13560 3754 13569
rect 3804 13530 3832 17478
rect 3896 16153 3924 17614
rect 3988 16794 4016 19774
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3882 16144 3938 16153
rect 3882 16079 3938 16088
rect 3896 15026 3924 16079
rect 3974 16008 4030 16017
rect 3974 15943 4030 15952
rect 3988 15638 4016 15943
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3896 13938 3924 14554
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3698 13495 3754 13504
rect 3792 13524 3844 13530
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3422 11928 3478 11937
rect 3422 11863 3478 11872
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3436 9178 3464 11698
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3422 9072 3478 9081
rect 3422 9007 3478 9016
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 2778 7239 2834 7248
rect 2872 7268 2924 7274
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 756 6860 808 6866
rect 756 6802 808 6808
rect 1214 6488 1270 6497
rect 1214 6423 1270 6432
rect 1228 5778 1256 6423
rect 2792 6322 2820 7239
rect 2872 7210 2924 7216
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 6338 3188 6734
rect 3344 6458 3372 7346
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3436 6338 3464 9007
rect 3528 8498 3556 13194
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3620 10198 3648 11834
rect 3712 10266 3740 13495
rect 3792 13466 3844 13472
rect 3896 11354 3924 13874
rect 3988 12850 4016 14214
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3988 12442 4016 12786
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3790 10704 3846 10713
rect 3790 10639 3846 10648
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3608 10192 3660 10198
rect 3660 10140 3740 10146
rect 3608 10134 3740 10140
rect 3620 10118 3740 10134
rect 3606 10024 3662 10033
rect 3606 9959 3662 9968
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 6662 3556 8230
rect 3620 7886 3648 9959
rect 3712 9489 3740 10118
rect 3698 9480 3754 9489
rect 3698 9415 3754 9424
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3712 8922 3740 9318
rect 3804 9042 3832 10639
rect 3882 10568 3938 10577
rect 3882 10503 3938 10512
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3712 8894 3832 8922
rect 3698 8392 3754 8401
rect 3698 8327 3700 8336
rect 3752 8327 3754 8336
rect 3700 8298 3752 8304
rect 3712 8090 3740 8298
rect 3804 8294 3832 8894
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3620 7546 3648 7822
rect 3698 7712 3754 7721
rect 3698 7647 3754 7656
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3606 7440 3662 7449
rect 3606 7375 3662 7384
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 2780 6316 2832 6322
rect 3160 6310 3464 6338
rect 2780 6258 2832 6264
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1320 6089 1348 6190
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 2792 5914 2820 6258
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 1216 5772 1268 5778
rect 1216 5714 1268 5720
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 2780 5704 2832 5710
rect 1360 5672 1362 5681
rect 2780 5646 2832 5652
rect 1306 5607 1362 5616
rect 2792 5370 2820 5646
rect 2884 5370 2912 6190
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 3620 5778 3648 7375
rect 3712 6322 3740 7647
rect 3804 6866 3832 7890
rect 3896 6934 3924 10503
rect 3988 9450 4016 12106
rect 4080 10130 4108 20046
rect 4250 19952 4306 19961
rect 4250 19887 4306 19896
rect 4264 19854 4292 19887
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4356 19446 4384 22066
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 4342 19136 4398 19145
rect 4342 19071 4398 19080
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4264 18329 4292 18702
rect 4250 18320 4306 18329
rect 4250 18255 4306 18264
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4172 15026 4200 17614
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4264 16726 4292 17546
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4356 16182 4384 19071
rect 4448 17270 4476 23582
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 4528 23044 4580 23050
rect 4528 22986 4580 22992
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4434 16960 4490 16969
rect 4434 16895 4490 16904
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4448 15570 4476 16895
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12306 4200 13330
rect 4252 13184 4304 13190
rect 4250 13152 4252 13161
rect 4304 13152 4306 13161
rect 4250 13087 4306 13096
rect 4356 12918 4384 15302
rect 4448 13705 4476 15506
rect 4434 13696 4490 13705
rect 4434 13631 4490 13640
rect 4540 13512 4568 22986
rect 4620 22500 4672 22506
rect 4620 22442 4672 22448
rect 4632 20534 4660 22442
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4710 19000 4766 19009
rect 4710 18935 4766 18944
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 17678 4660 18702
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4724 17490 4752 18935
rect 4632 17462 4752 17490
rect 4632 13734 4660 17462
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4724 15162 4752 15982
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4724 14074 4752 14214
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4816 13954 4844 22986
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4908 18034 4936 19314
rect 5000 18698 5028 23122
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26330 8078 27000
rect 7852 26302 8078 26330
rect 5264 24404 5316 24410
rect 5264 24346 5316 24352
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5276 22094 5304 24346
rect 5460 23662 5488 26200
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 6104 23186 6132 26200
rect 6460 24676 6512 24682
rect 6460 24618 6512 24624
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6288 23662 6316 24006
rect 6472 23866 6500 24618
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6564 23497 6592 23666
rect 6550 23488 6606 23497
rect 6550 23423 6606 23432
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 5724 22500 5776 22506
rect 5724 22442 5776 22448
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5184 22066 5304 22094
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 5000 18154 5028 18634
rect 5092 18630 5120 19722
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 4908 18006 5028 18034
rect 4894 17776 4950 17785
rect 4894 17711 4950 17720
rect 4908 14822 4936 17711
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4724 13926 4844 13954
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4448 13484 4568 13512
rect 4618 13560 4674 13569
rect 4618 13495 4674 13504
rect 4448 13308 4476 13484
rect 4448 13280 4568 13308
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4250 12744 4306 12753
rect 4250 12679 4306 12688
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4158 11248 4214 11257
rect 4158 11183 4160 11192
rect 4212 11183 4214 11192
rect 4160 11154 4212 11160
rect 4264 10674 4292 12679
rect 4356 12442 4384 12854
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4356 10554 4384 12174
rect 4264 10526 4384 10554
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4264 10062 4292 10526
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3974 9344 4030 9353
rect 3974 9279 4030 9288
rect 3988 8378 4016 9279
rect 4080 8498 4108 9590
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4264 9178 4292 9454
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4158 8936 4214 8945
rect 4158 8871 4214 8880
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3988 8350 4108 8378
rect 3974 7304 4030 7313
rect 3974 7239 3976 7248
rect 4028 7239 4030 7248
rect 3976 7210 4028 7216
rect 4080 6984 4108 8350
rect 4172 7426 4200 8871
rect 4250 8528 4306 8537
rect 4250 8463 4306 8472
rect 4264 7886 4292 8463
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4172 7410 4292 7426
rect 4172 7404 4304 7410
rect 4172 7398 4252 7404
rect 4252 7346 4304 7352
rect 4080 6956 4200 6984
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 4066 6896 4122 6905
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3896 5914 3924 6870
rect 4066 6831 4122 6840
rect 4080 6798 4108 6831
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3988 6662 4016 6734
rect 3976 6656 4028 6662
rect 4172 6610 4200 6956
rect 4356 6730 4384 10406
rect 4448 7546 4476 12854
rect 4540 9110 4568 13280
rect 4632 11830 4660 13495
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4724 9994 4752 13926
rect 4804 13864 4856 13870
rect 4908 13852 4936 14758
rect 4856 13824 4936 13852
rect 4804 13806 4856 13812
rect 4816 13530 4844 13806
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4816 12782 4844 12854
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4816 12238 4844 12378
rect 5000 12374 5028 18006
rect 5184 16590 5212 22066
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5276 20058 5304 20810
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5276 19786 5304 19994
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5368 18850 5396 22374
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5540 21480 5592 21486
rect 5538 21448 5540 21457
rect 5592 21448 5594 21457
rect 5538 21383 5594 21392
rect 5540 21344 5592 21350
rect 5644 21321 5672 21490
rect 5540 21286 5592 21292
rect 5630 21312 5686 21321
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5460 19922 5488 20878
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5276 18822 5396 18850
rect 5080 16584 5132 16590
rect 5078 16552 5080 16561
rect 5172 16584 5224 16590
rect 5132 16552 5134 16561
rect 5172 16526 5224 16532
rect 5078 16487 5134 16496
rect 5276 15994 5304 18822
rect 5356 18216 5408 18222
rect 5354 18184 5356 18193
rect 5408 18184 5410 18193
rect 5354 18119 5410 18128
rect 5368 17202 5396 18119
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5368 16794 5396 17002
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5184 15966 5304 15994
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5092 14482 5120 14758
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5092 13190 5120 14418
rect 5184 14414 5212 15966
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5276 13938 5304 15846
rect 5368 15638 5396 16730
rect 5356 15632 5408 15638
rect 5356 15574 5408 15580
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5368 14521 5396 15302
rect 5460 15201 5488 19450
rect 5552 15570 5580 21286
rect 5630 21247 5686 21256
rect 5630 20224 5686 20233
rect 5630 20159 5686 20168
rect 5644 18290 5672 20159
rect 5736 19514 5764 22442
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 5816 21616 5868 21622
rect 5816 21558 5868 21564
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5722 19408 5778 19417
rect 5722 19343 5724 19352
rect 5776 19343 5778 19352
rect 5724 19314 5776 19320
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 18057 5672 18226
rect 5736 18222 5764 19110
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5630 18048 5686 18057
rect 5630 17983 5686 17992
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5446 15192 5502 15201
rect 5446 15127 5502 15136
rect 5354 14512 5410 14521
rect 5354 14447 5410 14456
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 14006 5396 14282
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5184 12782 5212 13466
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4988 12368 5040 12374
rect 4894 12336 4950 12345
rect 4988 12310 5040 12316
rect 4894 12271 4950 12280
rect 4908 12238 4936 12271
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 11354 4936 12174
rect 5078 11928 5134 11937
rect 5078 11863 5134 11872
rect 5092 11393 5120 11863
rect 5276 11762 5304 13670
rect 5460 13394 5488 14350
rect 5644 14226 5672 16050
rect 5736 15065 5764 18158
rect 5828 16794 5856 21558
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5920 19310 5948 20742
rect 6104 20466 6132 21830
rect 6276 21616 6328 21622
rect 6276 21558 6328 21564
rect 6184 21412 6236 21418
rect 6184 21354 6236 21360
rect 6196 20874 6224 21354
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5920 18358 5948 19246
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5920 17785 5948 18158
rect 5906 17776 5962 17785
rect 5906 17711 5962 17720
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5906 16688 5962 16697
rect 6012 16658 6040 20402
rect 6196 20330 6224 20810
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6184 20324 6236 20330
rect 6184 20266 6236 20272
rect 6104 17202 6132 20266
rect 6196 18698 6224 20266
rect 6288 20058 6316 21558
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 6196 17610 6224 18634
rect 6380 18222 6408 22578
rect 6748 22166 6776 26200
rect 7392 24274 7420 26200
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 23089 6868 24142
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7196 23112 7248 23118
rect 6826 23080 6882 23089
rect 7196 23054 7248 23060
rect 6826 23015 6882 23024
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6460 21480 6512 21486
rect 6512 21428 6592 21434
rect 6460 21422 6592 21428
rect 6472 21406 6592 21422
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6472 20913 6500 21286
rect 6458 20904 6514 20913
rect 6458 20839 6514 20848
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6472 19417 6500 19450
rect 6458 19408 6514 19417
rect 6458 19343 6514 19352
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6184 17604 6236 17610
rect 6236 17564 6316 17592
rect 6184 17546 6236 17552
rect 6092 17196 6144 17202
rect 6144 17156 6224 17184
rect 6092 17138 6144 17144
rect 5906 16623 5908 16632
rect 5960 16623 5962 16632
rect 6000 16652 6052 16658
rect 5908 16594 5960 16600
rect 6000 16594 6052 16600
rect 6012 16402 6040 16594
rect 6012 16374 6132 16402
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 15570 5856 15846
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5920 15502 5948 15982
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5722 15056 5778 15065
rect 5722 14991 5778 15000
rect 5552 14198 5672 14226
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5460 11898 5488 12582
rect 5552 12170 5580 14198
rect 5828 13988 5856 15302
rect 5920 14929 5948 15438
rect 6012 15366 6040 16050
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5906 14920 5962 14929
rect 5906 14855 5962 14864
rect 5920 14278 5948 14855
rect 6012 14346 6040 15030
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5644 13960 5856 13988
rect 5644 13530 5672 13960
rect 6012 13920 6040 14282
rect 5828 13892 6040 13920
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5828 13326 5856 13892
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5920 13190 5948 13738
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5078 11384 5134 11393
rect 4896 11348 4948 11354
rect 5078 11319 5134 11328
rect 4896 11290 4948 11296
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 10130 4844 11086
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8809 4568 8910
rect 4526 8800 4582 8809
rect 4526 8735 4582 8744
rect 4540 8498 4568 8735
rect 5092 8566 5120 11319
rect 5552 11234 5580 11494
rect 5460 11206 5580 11234
rect 5170 11112 5226 11121
rect 5170 11047 5226 11056
rect 5184 9586 5212 11047
rect 5460 10962 5488 11206
rect 5460 10934 5580 10962
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 5184 8090 5212 9522
rect 5276 8362 5304 10474
rect 5368 8566 5396 10610
rect 5446 9616 5502 9625
rect 5446 9551 5502 9560
rect 5460 8974 5488 9551
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5368 8090 5396 8366
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 5184 7002 5212 8026
rect 5552 7478 5580 10934
rect 5644 10062 5672 12786
rect 5828 12782 5856 13126
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11558 5764 12106
rect 5920 11694 5948 13126
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11354 5764 11494
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5920 11234 5948 11630
rect 5828 11218 5948 11234
rect 5816 11212 5948 11218
rect 5868 11206 5948 11212
rect 5816 11154 5868 11160
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5906 9888 5962 9897
rect 5906 9823 5962 9832
rect 5814 9752 5870 9761
rect 5632 9716 5684 9722
rect 5814 9687 5870 9696
rect 5632 9658 5684 9664
rect 5540 7472 5592 7478
rect 5354 7440 5410 7449
rect 5540 7414 5592 7420
rect 5354 7375 5356 7384
rect 5408 7375 5410 7384
rect 5356 7346 5408 7352
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 3976 6598 4028 6604
rect 4080 6582 4200 6610
rect 4080 6118 4108 6582
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2976 5370 3004 5578
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 1306 5264 1362 5273
rect 1306 5199 1308 5208
rect 1360 5199 1362 5208
rect 1308 5170 1360 5176
rect 1320 4978 1348 5170
rect 1860 5024 1912 5030
rect 1320 4950 1440 4978
rect 1860 4966 1912 4972
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 1320 4690 1348 4791
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1412 4282 1440 4950
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1872 4146 1900 4966
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 664 3528 716 3534
rect 664 3470 716 3476
rect 1320 3233 1348 3538
rect 1306 3224 1362 3233
rect 1306 3159 1362 3168
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1320 2825 1348 2994
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1228 2417 1256 2450
rect 1214 2408 1270 2417
rect 1214 2343 1270 2352
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 2009 1348 2314
rect 1306 2000 1362 2009
rect 1306 1935 1362 1944
rect 1412 800 1440 4082
rect 2884 3641 2912 4558
rect 4158 4448 4214 4457
rect 4158 4383 4214 4392
rect 4172 4146 4200 4383
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2582 2820 2994
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2884 1601 2912 3470
rect 3344 3058 3372 3878
rect 4080 3534 4108 3975
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 5644 2990 5672 9658
rect 5828 9654 5856 9687
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5920 8294 5948 9823
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5724 8016 5776 8022
rect 5722 7984 5724 7993
rect 5776 7984 5778 7993
rect 5722 7919 5778 7928
rect 5736 7818 5764 7919
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 4080 800 4108 2450
rect 6012 2310 6040 13466
rect 6104 12442 6132 16374
rect 6196 15978 6224 17156
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 6288 15094 6316 17564
rect 6472 17202 6500 18634
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6458 17096 6514 17105
rect 6458 17031 6460 17040
rect 6512 17031 6514 17040
rect 6460 17002 6512 17008
rect 6472 16454 6500 17002
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6564 16046 6592 21406
rect 6656 20233 6684 21966
rect 6642 20224 6698 20233
rect 6642 20159 6698 20168
rect 6644 19712 6696 19718
rect 6644 19654 6696 19660
rect 6656 19378 6684 19654
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6656 17814 6684 18090
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6656 15502 6684 15982
rect 6748 15570 6776 18022
rect 6840 17066 6868 22578
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 20777 6960 21966
rect 6918 20768 6974 20777
rect 6918 20703 6974 20712
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6932 19174 6960 20538
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6932 16454 6960 19110
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6196 14482 6224 14962
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6288 14226 6316 14894
rect 6196 14198 6316 14226
rect 6196 13190 6224 14198
rect 6380 14074 6408 15302
rect 6472 14618 6500 15302
rect 6642 15056 6698 15065
rect 6642 14991 6698 15000
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6368 13864 6420 13870
rect 6366 13832 6368 13841
rect 6420 13832 6422 13841
rect 6366 13767 6422 13776
rect 6472 13734 6500 14214
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6196 10962 6224 13126
rect 6288 12850 6316 13262
rect 6472 12918 6500 13670
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6564 12764 6592 13738
rect 6380 12736 6592 12764
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6104 10934 6224 10962
rect 6104 6186 6132 10934
rect 6182 10840 6238 10849
rect 6182 10775 6238 10784
rect 6196 9042 6224 10775
rect 6288 10742 6316 12038
rect 6380 11558 6408 12736
rect 6656 12628 6684 14991
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6748 13870 6776 14554
rect 6840 14550 6868 16390
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6932 14822 6960 15506
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 7024 13512 7052 22646
rect 7116 22094 7144 22918
rect 7208 22681 7236 23054
rect 7194 22672 7250 22681
rect 7194 22607 7250 22616
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7116 22066 7236 22094
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7116 21457 7144 21490
rect 7102 21448 7158 21457
rect 7102 21383 7158 21392
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7116 19446 7144 21286
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7116 17814 7144 18634
rect 7104 17808 7156 17814
rect 7104 17750 7156 17756
rect 7102 17640 7158 17649
rect 7102 17575 7158 17584
rect 7116 15314 7144 17575
rect 7208 16250 7236 22066
rect 7300 21010 7328 22510
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7300 20398 7328 20946
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7300 18086 7328 20198
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7286 17776 7342 17785
rect 7286 17711 7342 17720
rect 7300 17610 7328 17711
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7392 17338 7420 23734
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7470 22672 7526 22681
rect 7470 22607 7526 22616
rect 7484 21146 7512 22607
rect 7576 21622 7604 23598
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7562 21312 7618 21321
rect 7562 21247 7618 21256
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7484 20942 7512 21082
rect 7576 21078 7604 21247
rect 7564 21072 7616 21078
rect 7564 21014 7616 21020
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7576 20466 7604 20742
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7484 19786 7512 20266
rect 7576 20097 7604 20402
rect 7562 20088 7618 20097
rect 7562 20023 7618 20032
rect 7472 19780 7524 19786
rect 7524 19740 7604 19768
rect 7472 19722 7524 19728
rect 7470 18728 7526 18737
rect 7576 18698 7604 19740
rect 7470 18663 7526 18672
rect 7564 18692 7616 18698
rect 7484 17542 7512 18663
rect 7564 18634 7616 18640
rect 7562 18184 7618 18193
rect 7562 18119 7564 18128
rect 7616 18119 7618 18128
rect 7564 18090 7616 18096
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7116 15286 7236 15314
rect 7102 15192 7158 15201
rect 7102 15127 7158 15136
rect 6932 13484 7052 13512
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12850 6868 13126
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6472 12600 6684 12628
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6288 10470 6316 10678
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6288 9722 6316 10406
rect 6380 10062 6408 11494
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6472 9466 6500 12600
rect 6550 12472 6606 12481
rect 6606 12416 6684 12434
rect 6550 12407 6684 12416
rect 6564 12406 6684 12407
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6288 9438 6500 9466
rect 6288 9382 6316 9438
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6564 8378 6592 10406
rect 6656 9602 6684 12406
rect 6748 12238 6776 12786
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6748 11354 6776 12174
rect 6840 11830 6868 12582
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6748 10198 6776 11290
rect 6932 10606 6960 13484
rect 7116 13410 7144 15127
rect 7208 14890 7236 15286
rect 7300 15026 7328 16458
rect 7484 15978 7512 17478
rect 7576 16794 7604 17478
rect 7668 17252 7696 23666
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7760 21010 7788 23258
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26330 10654 27000
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 8484 25084 8536 25090
rect 8484 25026 8536 25032
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7760 18358 7788 19994
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 7852 17814 7880 22578
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7944 21185 7972 21422
rect 7930 21176 7986 21185
rect 7930 21111 7986 21120
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 19938 8248 20198
rect 8312 20058 8340 24754
rect 8390 22128 8446 22137
rect 8390 22063 8446 22072
rect 8404 22030 8432 22063
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8220 19910 8340 19938
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 19242 8340 19910
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8404 18442 8432 20198
rect 8496 19446 8524 25026
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 22094 8616 24142
rect 8680 22574 8708 26200
rect 9324 24342 9352 26200
rect 9680 25628 9732 25634
rect 9680 25570 9732 25576
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9692 24070 9720 25570
rect 9862 24304 9918 24313
rect 9862 24239 9918 24248
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 8760 23248 8812 23254
rect 8760 23190 8812 23196
rect 8772 22574 8800 23190
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8760 22568 8812 22574
rect 8760 22510 8812 22516
rect 8588 22066 8708 22094
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8312 18414 8432 18442
rect 8312 18222 8340 18414
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8496 18272 8524 18770
rect 8588 18737 8616 19654
rect 8574 18728 8630 18737
rect 8574 18663 8630 18672
rect 8576 18284 8628 18290
rect 8496 18244 8576 18272
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 8220 17678 8248 18022
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7746 17368 7802 17377
rect 7950 17371 8258 17380
rect 7802 17312 7972 17320
rect 7746 17303 7972 17312
rect 7760 17292 7972 17303
rect 7668 17224 7788 17252
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7576 15366 7604 16730
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7484 15162 7512 15302
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7378 14920 7434 14929
rect 7196 14884 7248 14890
rect 7378 14855 7434 14864
rect 7196 14826 7248 14832
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14074 7328 14758
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7392 13852 7420 14855
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 13870 7604 14418
rect 7300 13824 7420 13852
rect 7564 13864 7616 13870
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7024 13382 7144 13410
rect 7024 10674 7052 13382
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 12306 7144 13194
rect 7208 12986 7236 13670
rect 7300 13376 7328 13824
rect 7564 13806 7616 13812
rect 7564 13388 7616 13394
rect 7300 13348 7512 13376
rect 7288 13252 7340 13258
rect 7340 13212 7420 13240
rect 7288 13194 7340 13200
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7392 12918 7420 13212
rect 7380 12912 7432 12918
rect 7194 12880 7250 12889
rect 7380 12854 7432 12860
rect 7194 12815 7250 12824
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 10418 6960 10542
rect 6932 10390 7052 10418
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6748 9722 6776 10134
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6656 9574 6960 9602
rect 6932 8566 6960 9574
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7024 8430 7052 10390
rect 7116 9994 7144 11222
rect 7208 11218 7236 12815
rect 7286 12744 7342 12753
rect 7286 12679 7342 12688
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 9382 7144 9930
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7194 9208 7250 9217
rect 7194 9143 7196 9152
rect 7248 9143 7250 9152
rect 7196 9114 7248 9120
rect 7300 8838 7328 12679
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12374 7420 12582
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7392 11762 7420 12310
rect 7484 12238 7512 13348
rect 7564 13330 7616 13336
rect 7576 12714 7604 13330
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7576 12050 7604 12378
rect 7484 12022 7604 12050
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7378 11248 7434 11257
rect 7378 11183 7434 11192
rect 7392 9586 7420 11183
rect 7484 11150 7512 12022
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7012 8424 7064 8430
rect 6564 8350 6684 8378
rect 7012 8366 7064 8372
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6550 8256 6606 8265
rect 6366 8120 6422 8129
rect 6366 8055 6368 8064
rect 6420 8055 6422 8064
rect 6368 8026 6420 8032
rect 6472 7342 6500 8230
rect 6550 8191 6606 8200
rect 6564 8090 6592 8191
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6656 8022 6684 8350
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 7392 7954 7420 9386
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7484 7886 7512 11086
rect 7562 9208 7618 9217
rect 7562 9143 7618 9152
rect 7576 8974 7604 9143
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7576 8090 7604 8910
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6840 4826 6868 7754
rect 7668 7546 7696 16050
rect 7760 12442 7788 17224
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 15638 7880 17138
rect 7944 17134 7972 17292
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 8206 17096 8262 17105
rect 8206 17031 8262 17040
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8128 16697 8156 16730
rect 8114 16688 8170 16697
rect 8114 16623 8116 16632
rect 8168 16623 8170 16632
rect 8116 16594 8168 16600
rect 8220 16454 8248 17031
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 7944 16017 7972 16050
rect 7930 16008 7986 16017
rect 7930 15943 7986 15952
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7944 15348 7972 15846
rect 7852 15320 7972 15348
rect 7852 14482 7880 15320
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7932 14952 7984 14958
rect 7930 14920 7932 14929
rect 7984 14920 7986 14929
rect 7930 14855 7986 14864
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7746 12200 7802 12209
rect 7746 12135 7802 12144
rect 7760 8498 7788 12135
rect 7852 11218 7880 14214
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7944 13190 7972 13806
rect 8312 13394 8340 18022
rect 8404 17882 8432 18226
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8390 17232 8446 17241
rect 8390 17167 8392 17176
rect 8444 17167 8446 17176
rect 8392 17138 8444 17144
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8404 16046 8432 16118
rect 8496 16114 8524 18244
rect 8576 18226 8628 18232
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8588 17610 8616 17818
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8574 17368 8630 17377
rect 8574 17303 8576 17312
rect 8628 17303 8630 17312
rect 8576 17274 8628 17280
rect 8588 16833 8616 17274
rect 8574 16824 8630 16833
rect 8574 16759 8630 16768
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8404 15570 8432 15982
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8496 15337 8524 15370
rect 8482 15328 8538 15337
rect 8482 15263 8538 15272
rect 8390 15192 8446 15201
rect 8496 15162 8524 15263
rect 8390 15127 8446 15136
rect 8484 15156 8536 15162
rect 8404 15094 8432 15127
rect 8484 15098 8536 15104
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8588 15026 8616 16662
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8404 14550 8432 14826
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 12374 8064 12718
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8128 11354 8156 11766
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8312 10826 8340 12038
rect 8404 11694 8432 13398
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8496 11150 8524 14826
rect 8574 14512 8630 14521
rect 8574 14447 8630 14456
rect 8588 14006 8616 14447
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 13462 8616 13738
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8574 11112 8630 11121
rect 8574 11047 8630 11056
rect 8312 10798 8524 10826
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 10130 7880 10406
rect 7840 10124 7892 10130
rect 8036 10112 8064 10678
rect 8128 10662 8340 10690
rect 8128 10606 8156 10662
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8116 10124 8168 10130
rect 8036 10084 8116 10112
rect 7840 10066 7892 10072
rect 8116 10066 8168 10072
rect 7852 9518 7880 10066
rect 8220 9976 8248 10542
rect 8312 10198 8340 10662
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8220 9948 8340 9976
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8312 9704 8340 9948
rect 8220 9676 8340 9704
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 8090 7788 8434
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 7852 3058 7880 9454
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7944 9110 7972 9386
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 8220 8974 8248 9676
rect 8496 9602 8524 10798
rect 8404 9574 8524 9602
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7930 8528 7986 8537
rect 7930 8463 7932 8472
rect 7984 8463 7986 8472
rect 8116 8492 8168 8498
rect 7932 8434 7984 8440
rect 8116 8434 8168 8440
rect 8128 7954 8156 8434
rect 8312 8090 8340 8774
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 8404 5234 8432 9574
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 9110 8524 9454
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8588 8634 8616 11047
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8576 8492 8628 8498
rect 8680 8480 8708 22066
rect 8760 22024 8812 22030
rect 8758 21992 8760 22001
rect 8812 21992 8814 22001
rect 8758 21927 8814 21936
rect 8956 21350 8984 23054
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9048 22166 9076 22918
rect 9036 22160 9088 22166
rect 9036 22102 9088 22108
rect 9048 21554 9076 22102
rect 9508 22094 9536 22986
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9416 22066 9536 22094
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8772 15706 8800 19314
rect 8864 18850 8892 20742
rect 8956 20398 8984 21286
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8956 19922 8984 20334
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 9140 18902 9168 20266
rect 9128 18896 9180 18902
rect 8864 18822 8984 18850
rect 9128 18838 9180 18844
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8864 17134 8892 18634
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8850 16280 8906 16289
rect 8850 16215 8852 16224
rect 8904 16215 8906 16224
rect 8852 16186 8904 16192
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8864 14278 8892 14962
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8772 12646 8800 12854
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8864 12102 8892 14214
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8864 11393 8892 11630
rect 8850 11384 8906 11393
rect 8850 11319 8906 11328
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8864 10674 8892 11222
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8772 9926 8800 10134
rect 8864 10062 8892 10610
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8772 9518 8800 9862
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 9042 8800 9318
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8628 8452 8708 8480
rect 8576 8434 8628 8440
rect 8760 8424 8812 8430
rect 8680 8384 8760 8412
rect 8680 8378 8708 8384
rect 8496 8362 8708 8378
rect 8760 8366 8812 8372
rect 8484 8356 8708 8362
rect 8536 8350 8708 8356
rect 8484 8298 8536 8304
rect 8864 6866 8892 9862
rect 8956 7410 8984 18822
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9140 18057 9168 18090
rect 9126 18048 9182 18057
rect 9126 17983 9182 17992
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 9048 16998 9076 17682
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9048 15094 9076 16458
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 11830 9076 13126
rect 9140 12170 9168 17614
rect 9232 15162 9260 21626
rect 9324 21026 9352 21830
rect 9416 21690 9444 22066
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9324 20998 9444 21026
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 18086 9352 20878
rect 9416 19009 9444 20998
rect 9600 20641 9628 22442
rect 9692 21010 9720 23462
rect 9784 22642 9812 23802
rect 9876 23730 9904 24239
rect 9968 23798 9996 26200
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 10060 24206 10088 25434
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9784 22545 9812 22578
rect 9770 22536 9826 22545
rect 9770 22471 9826 22480
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9586 20632 9642 20641
rect 9496 20596 9548 20602
rect 9586 20567 9642 20576
rect 9496 20538 9548 20544
rect 9508 19394 9536 20538
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9508 19366 9628 19394
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9402 19000 9458 19009
rect 9402 18935 9458 18944
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9416 17882 9444 18566
rect 9508 18154 9536 19178
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9494 18048 9550 18057
rect 9494 17983 9550 17992
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9324 14414 9352 16458
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9416 14278 9444 17546
rect 9508 16726 9536 17983
rect 9600 17626 9628 19366
rect 9692 17746 9720 20198
rect 9770 19544 9826 19553
rect 9770 19479 9826 19488
rect 9784 18970 9812 19479
rect 9968 19281 9996 21830
rect 10060 20058 10088 22034
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10152 20534 10180 21490
rect 10336 20874 10364 21490
rect 10428 21418 10456 21966
rect 10520 21894 10548 21966
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 21593 10548 21830
rect 10506 21584 10562 21593
rect 10506 21519 10562 21528
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10140 20528 10192 20534
rect 10140 20470 10192 20476
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10152 19802 10180 20470
rect 10416 19848 10468 19854
rect 10152 19796 10416 19802
rect 10152 19790 10468 19796
rect 10152 19786 10456 19790
rect 10140 19780 10456 19786
rect 10192 19774 10456 19780
rect 10140 19722 10192 19728
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 9954 19272 10010 19281
rect 9954 19207 10010 19216
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9600 17598 9720 17626
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9600 16538 9628 17274
rect 9508 16510 9628 16538
rect 9508 15366 9536 16510
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 15994 9628 16390
rect 9692 16250 9720 17598
rect 9784 17134 9812 18702
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17202 9904 18022
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 17128 9824 17134
rect 9876 17105 9904 17138
rect 9772 17070 9824 17076
rect 9862 17096 9918 17105
rect 9862 17031 9918 17040
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9784 16590 9812 16662
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9876 16522 9904 16662
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9772 16448 9824 16454
rect 9770 16416 9772 16425
rect 9824 16416 9826 16425
rect 9770 16351 9826 16360
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9784 16153 9812 16351
rect 9770 16144 9826 16153
rect 9770 16079 9826 16088
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9600 15966 9720 15994
rect 9692 15745 9720 15966
rect 9678 15736 9734 15745
rect 9678 15671 9734 15680
rect 9586 15464 9642 15473
rect 9586 15399 9642 15408
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9140 11762 9168 12106
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9034 11656 9090 11665
rect 9034 11591 9090 11600
rect 9048 8430 9076 11591
rect 9140 10266 9168 11698
rect 9232 11218 9260 14010
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9324 12306 9352 13806
rect 9402 13424 9458 13433
rect 9402 13359 9404 13368
rect 9456 13359 9458 13368
rect 9404 13330 9456 13336
rect 9508 12646 9536 13942
rect 9600 12889 9628 15399
rect 9876 15366 9904 16050
rect 9968 15473 9996 18226
rect 10060 17134 10088 18634
rect 10152 17746 10180 18838
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10048 17128 10100 17134
rect 10244 17082 10272 18770
rect 10336 17882 10364 19450
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10414 17912 10470 17921
rect 10324 17876 10376 17882
rect 10414 17847 10470 17856
rect 10324 17818 10376 17824
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10336 17202 10364 17478
rect 10428 17338 10456 17847
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10048 17070 10100 17076
rect 9954 15464 10010 15473
rect 9954 15399 10010 15408
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9692 14482 9720 14826
rect 9784 14482 9812 15030
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 13530 9812 14214
rect 9876 14006 9904 15302
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9586 12880 9642 12889
rect 9586 12815 9642 12824
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9600 12594 9628 12718
rect 9600 12566 9720 12594
rect 9692 12322 9720 12566
rect 9784 12374 9812 13466
rect 9968 12434 9996 15302
rect 10060 14482 10088 17070
rect 10152 17054 10272 17082
rect 10152 16114 10180 17054
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10152 12918 10180 16050
rect 10244 16046 10272 16934
rect 10336 16674 10364 17138
rect 10428 16833 10456 17274
rect 10414 16824 10470 16833
rect 10414 16759 10470 16768
rect 10336 16658 10456 16674
rect 10336 16652 10468 16658
rect 10336 16646 10416 16652
rect 10416 16594 10468 16600
rect 10520 16454 10548 18566
rect 10612 18086 10640 25094
rect 10704 22710 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10796 21894 10824 24822
rect 11150 24712 11206 24721
rect 11150 24647 11206 24656
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10508 16448 10560 16454
rect 10506 16416 10508 16425
rect 10560 16416 10562 16425
rect 10506 16351 10562 16360
rect 10704 16289 10732 21626
rect 10888 21486 10916 22442
rect 10980 21690 11008 22646
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10796 18068 10824 19314
rect 10980 19310 11008 20334
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10980 19174 11008 19246
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10888 18766 10916 19110
rect 11072 18970 11100 22102
rect 11164 21457 11192 24647
rect 11256 22098 11284 26200
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11716 24070 11744 24754
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11532 22982 11560 23462
rect 11808 23225 11836 23666
rect 11900 23610 11928 26200
rect 12072 25424 12124 25430
rect 12072 25366 12124 25372
rect 11900 23582 12020 23610
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 11794 23216 11850 23225
rect 11794 23151 11850 23160
rect 11520 22976 11572 22982
rect 11808 22953 11836 23151
rect 11520 22918 11572 22924
rect 11794 22944 11850 22953
rect 11794 22879 11850 22888
rect 11900 22817 11928 23462
rect 11992 22982 12020 23582
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11886 22808 11942 22817
rect 11886 22743 11942 22752
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11348 22166 11376 22374
rect 11900 22234 11928 22374
rect 11992 22234 12020 22510
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 11336 22160 11388 22166
rect 11336 22102 11388 22108
rect 11244 22092 11296 22098
rect 12084 22094 12112 25366
rect 12348 25356 12400 25362
rect 12348 25298 12400 25304
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 12268 23050 12296 23258
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12360 22930 12388 25298
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12452 23474 12480 24142
rect 12544 23798 12572 26200
rect 12716 25084 12768 25090
rect 12716 25026 12768 25032
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 12530 23488 12586 23497
rect 12452 23446 12530 23474
rect 12530 23423 12586 23432
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12268 22902 12388 22930
rect 12268 22642 12296 22902
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12268 22137 12296 22578
rect 12452 22574 12480 23122
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 11244 22034 11296 22040
rect 11992 22066 12112 22094
rect 12254 22128 12310 22137
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11150 21448 11206 21457
rect 11150 21383 11206 21392
rect 11532 21350 11560 21830
rect 11152 21344 11204 21350
rect 11520 21344 11572 21350
rect 11204 21304 11284 21332
rect 11152 21286 11204 21292
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11164 19718 11192 20198
rect 11256 19854 11284 21304
rect 11520 21286 11572 21292
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11348 20777 11376 20810
rect 11428 20800 11480 20806
rect 11334 20768 11390 20777
rect 11428 20742 11480 20748
rect 11334 20703 11390 20712
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11152 19712 11204 19718
rect 11204 19660 11284 19666
rect 11152 19654 11284 19660
rect 11164 19638 11284 19654
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 11256 18834 11284 19638
rect 11348 18873 11376 20198
rect 11440 19961 11468 20742
rect 11426 19952 11482 19961
rect 11426 19887 11482 19896
rect 11334 18864 11390 18873
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11244 18828 11296 18834
rect 11334 18799 11390 18808
rect 11244 18770 11296 18776
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 11072 18136 11100 18770
rect 11428 18216 11480 18222
rect 11426 18184 11428 18193
rect 11480 18184 11482 18193
rect 11072 18108 11192 18136
rect 11426 18119 11482 18128
rect 10796 18040 11100 18068
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10796 16697 10824 17138
rect 10888 16998 10916 17750
rect 11072 17241 11100 18040
rect 11058 17232 11114 17241
rect 11058 17167 11114 17176
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10874 16824 10930 16833
rect 10874 16759 10930 16768
rect 10888 16726 10916 16759
rect 10876 16720 10928 16726
rect 10782 16688 10838 16697
rect 10876 16662 10928 16668
rect 10782 16623 10838 16632
rect 11164 16561 11192 18108
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 17202 11376 17478
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11150 16552 11206 16561
rect 11150 16487 11206 16496
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 10690 16280 10746 16289
rect 10690 16215 10746 16224
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10244 15094 10272 15982
rect 10324 15632 10376 15638
rect 10324 15574 10376 15580
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 9968 12406 10088 12434
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9600 12294 9720 12322
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9140 9654 9168 9998
rect 9128 9648 9180 9654
rect 9180 9596 9260 9602
rect 9128 9590 9260 9596
rect 9140 9574 9260 9590
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9140 7546 9168 8842
rect 9232 8838 9260 9574
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9232 8430 9260 8774
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9232 8294 9260 8366
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7954 9260 8230
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 9324 5846 9352 12106
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 10674 9444 11494
rect 9508 11150 9536 11766
rect 9600 11626 9628 12294
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11234 9628 11562
rect 9600 11218 9720 11234
rect 9600 11212 9732 11218
rect 9600 11206 9680 11212
rect 9680 11154 9732 11160
rect 9876 11150 9904 11630
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9692 10266 9720 10610
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 9178 9720 9522
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 9042 9812 11018
rect 9876 10470 9904 11086
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9968 9654 9996 10950
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6748 800 6776 2450
rect 8312 2446 8340 2790
rect 9600 2650 9628 5782
rect 9692 4010 9720 8774
rect 9862 8392 9918 8401
rect 9862 8327 9864 8336
rect 9916 8327 9918 8336
rect 9864 8298 9916 8304
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9784 7750 9812 8026
rect 9968 7954 9996 9046
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 10060 4690 10088 12406
rect 10152 9178 10180 12718
rect 10244 12714 10272 14758
rect 10336 14414 10364 15574
rect 10704 15570 10732 16050
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10796 15094 10824 16118
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10416 14816 10468 14822
rect 10508 14816 10560 14822
rect 10416 14758 10468 14764
rect 10506 14784 10508 14793
rect 10560 14784 10562 14793
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10428 12238 10456 14758
rect 10506 14719 10562 14728
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10520 11558 10548 14418
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 12986 10640 14214
rect 10796 13870 10824 14826
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10690 12880 10746 12889
rect 10690 12815 10692 12824
rect 10744 12815 10746 12824
rect 10692 12786 10744 12792
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11830 10640 12038
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10336 8974 10364 10950
rect 10704 10606 10732 12786
rect 10796 11098 10824 13806
rect 10888 13274 10916 16050
rect 10966 16008 11022 16017
rect 10966 15943 10968 15952
rect 11020 15943 11022 15952
rect 10968 15914 11020 15920
rect 11164 15434 11192 16186
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11256 15162 11284 16390
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 10968 15088 11020 15094
rect 11348 15042 11376 17138
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 15337 11468 15846
rect 11426 15328 11482 15337
rect 11426 15263 11482 15272
rect 11426 15192 11482 15201
rect 11426 15127 11482 15136
rect 10968 15030 11020 15036
rect 10980 14618 11008 15030
rect 11256 15014 11376 15042
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10980 14278 11008 14554
rect 11072 14414 11100 14758
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11072 14226 11100 14350
rect 11072 14198 11192 14226
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10888 13246 11008 13274
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12442 10916 13126
rect 10980 12986 11008 13246
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12436 10928 12442
rect 11072 12434 11100 14010
rect 11164 13462 11192 14198
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11256 12442 11284 15014
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11244 12436 11296 12442
rect 11072 12406 11192 12434
rect 10876 12378 10928 12384
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11626 10916 12242
rect 10980 11762 11008 12310
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10796 11070 10916 11098
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10796 10266 10824 10950
rect 10888 10606 10916 11070
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9416 800 9444 2450
rect 9784 2446 9812 3130
rect 10336 3126 10364 8366
rect 10520 6866 10548 8434
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10612 3738 10640 8366
rect 10888 7954 10916 10542
rect 10980 10062 11008 10950
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 11058 10024 11114 10033
rect 11058 9959 11060 9968
rect 11112 9959 11114 9968
rect 11060 9930 11112 9936
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10980 7546 11008 8842
rect 11164 7886 11192 12406
rect 11244 12378 11296 12384
rect 11348 12306 11376 12582
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11256 11762 11284 12242
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10062 11284 10542
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9518 11284 9998
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11348 7410 11376 11290
rect 11440 10742 11468 15127
rect 11532 11121 11560 21286
rect 11808 21078 11836 21286
rect 11796 21072 11848 21078
rect 11796 21014 11848 21020
rect 11992 20942 12020 22066
rect 12254 22063 12310 22072
rect 12162 21448 12218 21457
rect 12162 21383 12218 21392
rect 11704 20936 11756 20942
rect 11980 20936 12032 20942
rect 11704 20878 11756 20884
rect 11794 20904 11850 20913
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11624 17338 11652 19314
rect 11716 19242 11744 20878
rect 11980 20878 12032 20884
rect 11794 20839 11850 20848
rect 11808 20534 11836 20839
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11808 20058 11836 20470
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 11794 19816 11850 19825
rect 11794 19751 11850 19760
rect 11808 19718 11836 19751
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11900 19417 11928 19450
rect 12084 19446 12112 19858
rect 11980 19440 12032 19446
rect 11886 19408 11942 19417
rect 11980 19382 12032 19388
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 11886 19343 11942 19352
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11886 18728 11942 18737
rect 11886 18663 11942 18672
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11716 16998 11744 18566
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11624 16561 11652 16730
rect 11610 16552 11666 16561
rect 11610 16487 11666 16496
rect 11716 16454 11744 16934
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11610 16280 11666 16289
rect 11610 16215 11612 16224
rect 11664 16215 11666 16224
rect 11612 16186 11664 16192
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11624 14006 11652 15302
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11518 11112 11574 11121
rect 11518 11047 11574 11056
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 11440 8566 11468 10678
rect 11624 10112 11652 12378
rect 11716 12102 11744 16390
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11808 11778 11836 18158
rect 11900 18086 11928 18663
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11900 17542 11928 17750
rect 11992 17678 12020 19382
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18290 12112 18566
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12176 17762 12204 21383
rect 12268 18306 12296 22063
rect 12452 21570 12480 22510
rect 12544 22137 12572 23423
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12530 22128 12586 22137
rect 12530 22063 12586 22072
rect 12452 21554 12572 21570
rect 12452 21548 12584 21554
rect 12452 21542 12532 21548
rect 12452 20534 12480 21542
rect 12532 21490 12584 21496
rect 12636 21010 12664 22918
rect 12728 21962 12756 25026
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13280 23633 13308 23666
rect 13266 23624 13322 23633
rect 13266 23559 13322 23568
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22710 12848 22918
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 13280 22574 13308 23122
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13372 22098 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 13636 24676 13688 24682
rect 13636 24618 13688 24624
rect 13648 23050 13676 24618
rect 13832 24138 13860 26200
rect 14372 24268 14424 24274
rect 14476 24256 14504 26200
rect 15016 25016 15068 25022
rect 15016 24958 15068 24964
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14646 24848 14702 24857
rect 14646 24783 14702 24792
rect 14424 24228 14504 24256
rect 14372 24210 14424 24216
rect 14556 24200 14608 24206
rect 14278 24168 14334 24177
rect 13820 24132 13872 24138
rect 14556 24142 14608 24148
rect 14278 24103 14334 24112
rect 13820 24074 13872 24080
rect 14292 24070 14320 24103
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13636 23044 13688 23050
rect 13636 22986 13688 22992
rect 13832 22642 13860 23258
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 13464 21622 13492 22374
rect 13832 21622 13860 22578
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12452 19990 12480 20470
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12268 18278 12388 18306
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12084 17734 12204 17762
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11900 16522 11928 16594
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11992 16114 12020 17614
rect 12084 17184 12112 17734
rect 12268 17610 12296 18090
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12176 17513 12204 17546
rect 12162 17504 12218 17513
rect 12162 17439 12218 17448
rect 12084 17156 12204 17184
rect 12176 16674 12204 17156
rect 12084 16646 12204 16674
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 12084 15722 12112 16646
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11992 15694 12112 15722
rect 11992 15144 12020 15694
rect 12176 15638 12204 16390
rect 12268 16250 12296 17546
rect 12360 16726 12388 18278
rect 12544 17354 12572 20198
rect 12728 19922 12756 21558
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12716 19780 12768 19786
rect 12716 19722 12768 19728
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12452 17326 12572 17354
rect 12348 16720 12400 16726
rect 12348 16662 12400 16668
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12254 15736 12310 15745
rect 12254 15671 12310 15680
rect 12072 15632 12124 15638
rect 12070 15600 12072 15609
rect 12164 15632 12216 15638
rect 12124 15600 12126 15609
rect 12164 15574 12216 15580
rect 12070 15535 12126 15544
rect 12268 15434 12296 15671
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 11900 15116 12020 15144
rect 11900 13938 11928 15116
rect 11978 15056 12034 15065
rect 11978 14991 11980 15000
rect 12032 14991 12034 15000
rect 11980 14962 12032 14968
rect 11980 14408 12032 14414
rect 12360 14385 12388 16458
rect 11980 14350 12032 14356
rect 12346 14376 12402 14385
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 13462 11928 13874
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11900 13161 11928 13398
rect 11992 13394 12020 14350
rect 12346 14311 12402 14320
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11886 13152 11942 13161
rect 11886 13087 11942 13096
rect 12176 12646 12204 13806
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12268 12306 12296 12650
rect 12360 12306 12388 13194
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11716 11750 11836 11778
rect 11716 10266 11744 11750
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 10470 11836 11630
rect 11900 10674 11928 12106
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11532 10084 11652 10112
rect 11532 9178 11560 10084
rect 11610 10024 11666 10033
rect 11808 9994 11836 10406
rect 11992 10248 12020 12038
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12084 10742 12112 11698
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11992 10220 12112 10248
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11610 9959 11666 9968
rect 11796 9988 11848 9994
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11624 8498 11652 9959
rect 11796 9930 11848 9936
rect 11888 9920 11940 9926
rect 11992 9874 12020 10066
rect 11940 9868 12020 9874
rect 11888 9862 12020 9868
rect 11900 9846 12020 9862
rect 11992 9654 12020 9846
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 12084 8090 12112 10220
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11532 7342 11560 7822
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 12084 3738 12112 7414
rect 12176 6390 12204 12242
rect 12268 11558 12296 12242
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12360 11354 12388 12242
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12452 10690 12480 17326
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12544 16794 12572 17138
rect 12636 16946 12664 18226
rect 12728 18086 12756 19722
rect 12820 18850 12848 21286
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13832 21146 13860 21558
rect 14004 21344 14056 21350
rect 13910 21312 13966 21321
rect 14004 21286 14056 21292
rect 13910 21247 13966 21256
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13924 20806 13952 21247
rect 13912 20800 13964 20806
rect 13910 20768 13912 20777
rect 13964 20768 13966 20777
rect 13910 20703 13966 20712
rect 14016 20534 14044 21286
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 13358 20360 13414 20369
rect 13358 20295 13414 20304
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 20058 13400 20295
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13280 19446 13308 19654
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12820 18822 12940 18850
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12820 18358 12848 18634
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12912 18136 12940 18822
rect 13372 18329 13400 19178
rect 13464 19009 13492 20198
rect 13450 19000 13506 19009
rect 13450 18935 13506 18944
rect 13556 18834 13584 20470
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13648 19394 13676 20198
rect 13740 19553 13768 20198
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13726 19544 13782 19553
rect 13726 19479 13782 19488
rect 13648 19366 13768 19394
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13358 18320 13414 18329
rect 13358 18255 13414 18264
rect 12820 18108 12940 18136
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12820 17592 12848 18108
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17678 13400 18022
rect 13648 17814 13676 19246
rect 13740 19145 13768 19366
rect 13832 19242 13860 19654
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13726 19136 13782 19145
rect 13726 19071 13782 19080
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13740 18601 13768 18838
rect 13726 18592 13782 18601
rect 13726 18527 13782 18536
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 12820 17564 13032 17592
rect 13004 17513 13032 17564
rect 12806 17504 12862 17513
rect 12806 17439 12862 17448
rect 12990 17504 13046 17513
rect 12990 17439 13046 17448
rect 12820 16998 12848 17439
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13096 17134 13124 17274
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12808 16992 12860 16998
rect 12636 16918 12756 16946
rect 12808 16934 12860 16940
rect 12622 16824 12678 16833
rect 12532 16788 12584 16794
rect 12622 16759 12624 16768
rect 12532 16730 12584 16736
rect 12676 16759 12678 16768
rect 12624 16730 12676 16736
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12544 16182 12572 16526
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12532 15360 12584 15366
rect 12636 15337 12664 15846
rect 12532 15302 12584 15308
rect 12622 15328 12678 15337
rect 12544 12442 12572 15302
rect 12622 15263 12678 15272
rect 12728 15162 12756 16918
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12820 15706 12848 16458
rect 13372 16114 13400 17614
rect 13648 17338 13676 17750
rect 13740 17338 13768 18362
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 13372 15570 13400 16050
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12912 15026 12940 15506
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12636 14482 12664 14962
rect 13280 14958 13308 15098
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 14482 12756 14758
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14618 13400 14962
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12636 13938 12664 14418
rect 13360 14408 13412 14414
rect 12898 14376 12954 14385
rect 13360 14350 13412 14356
rect 12898 14311 12954 14320
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12912 13870 12940 14311
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 13530 12756 13738
rect 13188 13734 13216 13874
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12716 13524 12768 13530
rect 13372 13512 13400 14350
rect 12716 13466 12768 13472
rect 13188 13484 13400 13512
rect 13188 13240 13216 13484
rect 13268 13388 13320 13394
rect 13320 13348 13400 13376
rect 13268 13330 13320 13336
rect 13268 13252 13320 13258
rect 13188 13212 13268 13240
rect 13188 12918 13216 13212
rect 13268 13194 13320 13200
rect 13372 12918 13400 13348
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 12728 12442 12756 12854
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12900 12640 12952 12646
rect 12820 12600 12900 12628
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12820 11286 12848 12600
rect 13096 12628 13124 12786
rect 12952 12600 13124 12628
rect 12900 12582 12952 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12912 11626 12940 12106
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 13280 11540 13308 12174
rect 13372 11830 13400 12854
rect 13464 12374 13492 17138
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16561 13860 17070
rect 13818 16552 13874 16561
rect 13818 16487 13874 16496
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13556 14958 13584 15982
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13556 14618 13584 14894
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13280 11512 13400 11540
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13372 11354 13400 11512
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 12360 10662 12480 10690
rect 12360 9722 12388 10662
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12452 8634 12480 10542
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12820 9874 12848 9930
rect 12728 9846 12848 9874
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8634 12572 8774
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12438 8528 12494 8537
rect 12728 8498 12756 9846
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12820 9217 12848 9658
rect 13372 9450 13400 11154
rect 13556 10130 13584 13874
rect 13648 13870 13676 15846
rect 13726 15736 13782 15745
rect 13726 15671 13782 15680
rect 13740 15502 13768 15671
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13530 13676 13670
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13740 12986 13768 15302
rect 13818 15192 13874 15201
rect 13818 15127 13874 15136
rect 13832 14822 13860 15127
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13648 12866 13676 12922
rect 13924 12866 13952 19314
rect 14016 19310 14044 20470
rect 14292 20233 14320 23462
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14384 22409 14412 22986
rect 14464 22976 14516 22982
rect 14568 22953 14596 24142
rect 14464 22918 14516 22924
rect 14554 22944 14610 22953
rect 14476 22778 14504 22918
rect 14554 22879 14610 22888
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14370 22400 14426 22409
rect 14370 22335 14426 22344
rect 14568 22234 14596 22879
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 14660 22094 14688 24783
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14568 22066 14688 22094
rect 14568 22030 14596 22066
rect 14556 22024 14608 22030
rect 14554 21992 14556 22001
rect 14608 21992 14610 22001
rect 14554 21927 14610 21936
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14660 21622 14688 21830
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14476 20534 14504 21082
rect 14752 20890 14780 24278
rect 14660 20862 14780 20890
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14278 20224 14334 20233
rect 14278 20159 14334 20168
rect 14292 19990 14320 20159
rect 14476 19990 14504 20470
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 14476 19718 14504 19926
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14568 19514 14596 19790
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14016 18193 14044 19246
rect 14372 19236 14424 19242
rect 14372 19178 14424 19184
rect 14186 18320 14242 18329
rect 14186 18255 14242 18264
rect 14002 18184 14058 18193
rect 14002 18119 14058 18128
rect 14200 15722 14228 18255
rect 14384 17746 14412 19178
rect 14464 18896 14516 18902
rect 14462 18864 14464 18873
rect 14516 18864 14518 18873
rect 14462 18799 14518 18808
rect 14568 18358 14596 19450
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14462 17640 14518 17649
rect 14462 17575 14518 17584
rect 14476 17542 14504 17575
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14370 16552 14426 16561
rect 14370 16487 14426 16496
rect 14384 16454 14412 16487
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14016 15694 14228 15722
rect 14016 12986 14044 15694
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 14618 14136 15506
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14108 14414 14136 14554
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13938 14136 14350
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14200 13190 14228 15302
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14414 14320 14894
rect 14384 14793 14412 14962
rect 14370 14784 14426 14793
rect 14370 14719 14426 14728
rect 14370 14648 14426 14657
rect 14370 14583 14372 14592
rect 14424 14583 14426 14592
rect 14372 14554 14424 14560
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 13326 14320 14350
rect 14384 13920 14412 14554
rect 14476 14074 14504 16594
rect 14568 14482 14596 18022
rect 14660 15366 14688 20862
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 16250 14780 20742
rect 14844 19786 14872 24890
rect 15028 22642 15056 24958
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15120 22098 15148 26200
rect 15474 25256 15530 25265
rect 15384 25220 15436 25226
rect 15474 25191 15530 25200
rect 15384 25162 15436 25168
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14936 21078 14964 21830
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 15028 21010 15056 21286
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15212 20942 15240 21966
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14844 19514 14872 19722
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14844 18834 14872 19450
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 17921 14872 18566
rect 14830 17912 14886 17921
rect 14830 17847 14886 17856
rect 14936 17678 14964 19246
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15028 18970 15056 19110
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 15028 18358 15056 18634
rect 15120 18465 15148 19178
rect 15212 18873 15240 20334
rect 15304 19904 15332 24074
rect 15396 22030 15424 25162
rect 15488 23118 15516 25191
rect 15658 25120 15714 25129
rect 15658 25055 15714 25064
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15566 21448 15622 21457
rect 15566 21383 15568 21392
rect 15620 21383 15622 21392
rect 15568 21354 15620 21360
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15488 19922 15516 20266
rect 15476 19916 15528 19922
rect 15304 19876 15424 19904
rect 15396 18873 15424 19876
rect 15476 19858 15528 19864
rect 15672 19378 15700 25055
rect 15764 23798 15792 26200
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 16026 23488 16082 23497
rect 16026 23423 16082 23432
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15752 20800 15804 20806
rect 15750 20768 15752 20777
rect 15804 20768 15806 20777
rect 15750 20703 15806 20712
rect 15856 19378 15884 23122
rect 16040 21690 16068 23423
rect 16132 22710 16160 26302
rect 16394 26200 16450 26302
rect 17038 26330 17094 27000
rect 17682 26330 17738 27000
rect 17038 26302 17356 26330
rect 17038 26200 17094 26302
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 16500 23769 16528 24346
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16486 23760 16542 23769
rect 16486 23695 16542 23704
rect 16592 23526 16620 24142
rect 17144 24138 17172 24618
rect 17132 24132 17184 24138
rect 17132 24074 17184 24080
rect 17040 24064 17092 24070
rect 17040 24006 17092 24012
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 15948 21593 15976 21626
rect 15934 21584 15990 21593
rect 15934 21519 15936 21528
rect 15988 21519 15990 21528
rect 15936 21490 15988 21496
rect 16224 21010 16252 21626
rect 16408 21010 16436 22170
rect 16684 21418 16712 22646
rect 16868 22574 16896 23054
rect 16960 23050 16988 23666
rect 17052 23594 17080 24006
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 17052 23050 17080 23530
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16672 21412 16724 21418
rect 16672 21354 16724 21360
rect 16578 21176 16634 21185
rect 16578 21111 16580 21120
rect 16632 21111 16634 21120
rect 16580 21082 16632 21088
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16118 20632 16174 20641
rect 16118 20567 16120 20576
rect 16172 20567 16174 20576
rect 16120 20538 16172 20544
rect 16684 20466 16712 21354
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15198 18864 15254 18873
rect 15198 18799 15254 18808
rect 15382 18864 15438 18873
rect 15382 18799 15438 18808
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15106 18456 15162 18465
rect 15106 18391 15162 18400
rect 15016 18352 15068 18358
rect 15016 18294 15068 18300
rect 15108 18216 15160 18222
rect 15014 18184 15070 18193
rect 15108 18158 15160 18164
rect 15014 18119 15016 18128
rect 15068 18119 15070 18128
rect 15016 18090 15068 18096
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 15120 17542 15148 18158
rect 15304 17898 15332 18566
rect 15212 17870 15332 17898
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14752 15502 14780 15846
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14384 13892 14504 13920
rect 14476 13852 14504 13892
rect 14556 13864 14608 13870
rect 14476 13824 14556 13852
rect 14556 13806 14608 13812
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 13648 12838 13952 12866
rect 14200 12442 14228 12922
rect 14292 12918 14320 13262
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 13740 12238 13768 12378
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11150 13768 12174
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10962 13768 11086
rect 13820 11008 13872 11014
rect 13740 10956 13820 10962
rect 13740 10950 13872 10956
rect 13740 10934 13860 10950
rect 13832 10742 13860 10934
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13832 9926 13860 10678
rect 14200 10266 14228 11154
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9654 13860 9862
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12806 9208 12862 9217
rect 12950 9211 13258 9220
rect 12806 9143 12862 9152
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 12438 8463 12494 8472
rect 12716 8492 12768 8498
rect 12452 8090 12480 8463
rect 12716 8434 12768 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12452 7954 12480 8026
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12452 5234 12480 7142
rect 12636 5846 12664 8366
rect 13924 8362 13952 8774
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 14016 8090 14044 9318
rect 14200 9178 14228 10202
rect 14384 9654 14412 13738
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14476 11150 14504 12174
rect 14568 12170 14596 12378
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14660 11354 14688 15302
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14752 14074 14780 15030
rect 14844 14278 14872 16390
rect 14936 16114 14964 17478
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 14936 14618 14964 15030
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14936 13870 14964 14554
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 15028 13530 15056 15506
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14752 12084 14780 12786
rect 14924 12096 14976 12102
rect 14752 12056 14924 12084
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14476 10062 14504 11086
rect 14752 10810 14780 12056
rect 14924 12038 14976 12044
rect 15028 11694 15056 13466
rect 15120 12850 15148 17478
rect 15212 16454 15240 17870
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15304 17202 15332 17750
rect 15396 17678 15424 18799
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15396 16590 15424 17478
rect 15488 17134 15516 18634
rect 15672 18086 15700 19314
rect 16040 18290 16068 19858
rect 16684 19786 16712 20198
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16316 18850 16344 19246
rect 16224 18834 16344 18850
rect 16212 18828 16344 18834
rect 16264 18822 16344 18828
rect 16212 18770 16264 18776
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 14346 15240 15846
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15304 14226 15332 16526
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15488 15162 15516 15302
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15304 14198 15424 14226
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15212 12782 15240 13330
rect 15304 13258 15332 13738
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15304 12374 15332 12718
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15304 11558 15332 11766
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14200 7954 14228 8026
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12084 3534 12112 3674
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 11624 2582 11652 3334
rect 12636 3126 12664 5646
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13464 3670 13492 7822
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13556 7546 13584 7754
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 14292 7410 14320 9386
rect 14384 9042 14412 9590
rect 14476 9518 14504 9998
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14752 8566 14780 9454
rect 14936 8634 14964 10610
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15212 10130 15240 10542
rect 15304 10146 15332 10950
rect 15396 10810 15424 14198
rect 15488 13802 15516 14282
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15488 12374 15516 12650
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15200 10124 15252 10130
rect 15304 10118 15424 10146
rect 15200 10066 15252 10072
rect 15396 9110 15424 10118
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15396 8566 15424 9046
rect 15580 8838 15608 13874
rect 15672 10538 15700 17138
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15764 12209 15792 16934
rect 15856 15706 15884 17070
rect 16132 17066 16160 17818
rect 16316 17746 16344 18822
rect 16408 18630 16436 19654
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16486 18320 16542 18329
rect 16486 18255 16488 18264
rect 16540 18255 16542 18264
rect 16488 18226 16540 18232
rect 16486 17776 16542 17785
rect 16304 17740 16356 17746
rect 16486 17711 16542 17720
rect 16304 17682 16356 17688
rect 16210 17640 16266 17649
rect 16210 17575 16266 17584
rect 16304 17604 16356 17610
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 16224 16794 16252 17575
rect 16304 17546 16356 17552
rect 16316 16794 16344 17546
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 16448 16172 16454
rect 16212 16448 16264 16454
rect 16120 16390 16172 16396
rect 16210 16416 16212 16425
rect 16264 16416 16266 16425
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 16132 15570 16160 16390
rect 16210 16351 16266 16360
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16224 15502 16252 15846
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16316 14822 16344 16594
rect 16408 16114 16436 17478
rect 16500 16833 16528 17711
rect 16486 16824 16542 16833
rect 16486 16759 16542 16768
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 14822 16436 15302
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16316 14482 16344 14758
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12306 15884 13126
rect 16040 12986 16068 13806
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16132 12918 16160 13738
rect 16408 13394 16436 14214
rect 16500 13394 16528 16118
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15750 12200 15806 12209
rect 15750 12135 15806 12144
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15948 9178 15976 11698
rect 16132 11558 16160 12854
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11150 16160 11494
rect 16224 11354 16252 12242
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16132 9382 16160 10542
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9722 16252 10066
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 9194 16160 9318
rect 15936 9172 15988 9178
rect 16132 9166 16252 9194
rect 15936 9114 15988 9120
rect 16224 8906 16252 9166
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 16316 8634 16344 10542
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16500 9178 16528 10474
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 16120 8560 16172 8566
rect 16592 8537 16620 19450
rect 16684 18834 16712 19722
rect 16868 19310 16896 22510
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16960 20602 16988 20742
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16960 19514 16988 20266
rect 17052 19990 17080 20742
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16684 18426 16712 18770
rect 16776 18766 16804 19178
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16672 18420 16724 18426
rect 16724 18380 16804 18408
rect 16672 18362 16724 18368
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16684 16522 16712 18226
rect 16776 17882 16804 18380
rect 16960 18222 16988 18566
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16776 17592 16804 17818
rect 16960 17746 16988 18158
rect 17052 17746 17080 19450
rect 17144 19258 17172 23734
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17236 21078 17264 22918
rect 17328 21486 17356 26302
rect 17420 26302 17738 26330
rect 17420 23186 17448 26302
rect 17682 26200 17738 26302
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26330 21602 27000
rect 21546 26302 22048 26330
rect 21546 26200 21602 26302
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17512 22681 17540 23666
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17590 23216 17646 23225
rect 17590 23151 17646 23160
rect 17604 22953 17632 23151
rect 17590 22944 17646 22953
rect 17590 22879 17646 22888
rect 17498 22672 17554 22681
rect 17498 22607 17554 22616
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 17512 21026 17540 21898
rect 17512 20998 17632 21026
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17224 19984 17276 19990
rect 17222 19952 17224 19961
rect 17276 19952 17278 19961
rect 17222 19887 17278 19896
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17144 19230 17356 19258
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16776 17564 16988 17592
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16776 16794 16804 16934
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 14006 16712 16050
rect 16776 14890 16804 16390
rect 16868 14958 16896 16934
rect 16960 16522 16988 17564
rect 17144 17202 17172 17818
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16948 16176 17000 16182
rect 16946 16144 16948 16153
rect 17000 16144 17002 16153
rect 16946 16079 17002 16088
rect 17052 15502 17080 17002
rect 17236 16658 17264 17138
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17130 16280 17186 16289
rect 17130 16215 17132 16224
rect 17184 16215 17186 16224
rect 17132 16186 17184 16192
rect 17236 16046 17264 16458
rect 17328 16046 17356 19230
rect 17420 18306 17448 19314
rect 17512 18834 17540 20878
rect 17604 20466 17632 20998
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 18902 17632 19654
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17420 18278 17632 18306
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 17052 14498 17080 15438
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 14929 17172 14962
rect 17130 14920 17186 14929
rect 17130 14855 17186 14864
rect 17052 14482 17172 14498
rect 17052 14476 17184 14482
rect 17052 14470 17132 14476
rect 17132 14418 17184 14424
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 17144 13870 17172 14418
rect 17236 14074 17264 14418
rect 17328 14074 17356 15370
rect 17420 15366 17448 17070
rect 17512 16998 17540 18158
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17420 14346 17448 15302
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17512 13870 17540 15914
rect 17604 14822 17632 18278
rect 17696 17814 17724 23462
rect 17788 22817 17816 25230
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23662 18368 26200
rect 18604 24676 18656 24682
rect 18604 24618 18656 24624
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17774 22808 17830 22817
rect 17950 22811 18258 22820
rect 17774 22743 17830 22752
rect 17788 20777 17816 22743
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17866 20904 17922 20913
rect 17866 20839 17868 20848
rect 17920 20839 17922 20848
rect 17868 20810 17920 20816
rect 18328 20800 18380 20806
rect 17774 20768 17830 20777
rect 18328 20742 18380 20748
rect 17774 20703 17830 20712
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17972 20233 18000 20334
rect 17958 20224 18014 20233
rect 17958 20159 18014 20168
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17972 19802 18000 19994
rect 18340 19854 18368 20742
rect 17880 19774 18000 19802
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18432 19802 18460 24142
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18524 23118 18552 24074
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18524 22710 18552 23054
rect 18616 22778 18644 24618
rect 18984 24410 19012 26200
rect 19154 24440 19210 24449
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 19064 24404 19116 24410
rect 19628 24426 19656 26200
rect 19154 24375 19210 24384
rect 19352 24398 19656 24426
rect 19064 24346 19116 24352
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18708 23730 18736 24210
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18708 23526 18736 23666
rect 19076 23662 19104 24346
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 19076 23254 19104 23598
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 19168 23066 19196 24375
rect 19248 23792 19300 23798
rect 19352 23746 19380 24398
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19524 24132 19576 24138
rect 19524 24074 19576 24080
rect 19536 23798 19564 24074
rect 19300 23740 19380 23746
rect 19248 23734 19380 23740
rect 19524 23792 19576 23798
rect 19524 23734 19576 23740
rect 19260 23718 19380 23734
rect 19800 23112 19852 23118
rect 19168 23038 19564 23066
rect 19800 23054 19852 23060
rect 19536 22817 19564 23038
rect 19522 22808 19578 22817
rect 18604 22772 18656 22778
rect 19522 22743 19578 22752
rect 18604 22714 18656 22720
rect 18512 22704 18564 22710
rect 18512 22646 18564 22652
rect 18524 22166 18552 22646
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18512 22160 18564 22166
rect 18512 22102 18564 22108
rect 18524 22030 18552 22102
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18616 21554 18644 22510
rect 19156 22432 19208 22438
rect 19156 22374 19208 22380
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18800 21434 18828 21830
rect 18616 21418 18828 21434
rect 18604 21412 18828 21418
rect 18656 21406 18828 21412
rect 18604 21354 18656 21360
rect 18696 21344 18748 21350
rect 18602 21312 18658 21321
rect 18892 21332 18920 21966
rect 19076 21486 19104 22102
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18748 21304 18920 21332
rect 18696 21286 18748 21292
rect 18602 21247 18658 21256
rect 18616 21010 18644 21247
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18602 20088 18658 20097
rect 18602 20023 18658 20032
rect 18432 19774 18552 19802
rect 17880 19496 17908 19774
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17880 19468 18000 19496
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17880 19174 17908 19314
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17972 18630 18000 19468
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17696 16454 17724 17614
rect 17684 16448 17736 16454
rect 17736 16408 17816 16436
rect 17684 16390 17736 16396
rect 17788 15434 17816 16408
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17788 15094 17816 15370
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13258 17080 13670
rect 17144 13394 17172 13806
rect 17512 13530 17540 13806
rect 17696 13716 17724 13942
rect 17880 13870 17908 18022
rect 18340 17542 18368 18022
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 17270 18368 17478
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18340 16726 18368 17206
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18156 14550 18184 15030
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18156 14362 18184 14486
rect 18340 14482 18368 16526
rect 18432 15162 18460 19654
rect 18524 16454 18552 19774
rect 18616 19689 18644 20023
rect 18602 19680 18658 19689
rect 18602 19615 18658 19624
rect 18800 19174 18828 20946
rect 18892 20942 18920 21304
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18892 20602 18920 20878
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18984 19922 19012 21422
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19076 19514 19104 19790
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18788 19168 18840 19174
rect 18694 19136 18750 19145
rect 18788 19110 18840 19116
rect 18694 19071 18750 19080
rect 18602 19000 18658 19009
rect 18602 18935 18658 18944
rect 18616 18834 18644 18935
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18708 18630 18736 19071
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 17626 18736 18566
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18708 17598 18828 17626
rect 18892 17610 18920 18158
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 16250 18644 16390
rect 18708 16250 18736 17478
rect 18800 17377 18828 17598
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18786 17368 18842 17377
rect 18842 17326 18920 17354
rect 18786 17303 18842 17312
rect 18786 16824 18842 16833
rect 18786 16759 18842 16768
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18510 15192 18566 15201
rect 18420 15156 18472 15162
rect 18510 15127 18566 15136
rect 18420 15098 18472 15104
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18156 14346 18368 14362
rect 18144 14340 18368 14346
rect 18196 14334 18368 14340
rect 18144 14282 18196 14288
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18144 14000 18196 14006
rect 18340 13954 18368 14334
rect 18196 13948 18368 13954
rect 18144 13942 18368 13948
rect 18156 13926 18368 13942
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 18156 13716 18184 13926
rect 17696 13688 18184 13716
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12850 17080 13194
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17512 12714 17540 13330
rect 18156 13258 18184 13688
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18432 12918 18460 15098
rect 18524 14793 18552 15127
rect 18510 14784 18566 14793
rect 18800 14770 18828 16759
rect 18510 14719 18566 14728
rect 18616 14742 18828 14770
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17408 12096 17460 12102
rect 17406 12064 17408 12073
rect 17460 12064 17462 12073
rect 17406 11999 17462 12008
rect 17420 11898 17448 11999
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 9926 16804 10950
rect 16868 10062 16896 11086
rect 16960 10742 16988 11494
rect 17052 10810 17080 11630
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9654 16804 9862
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16868 9518 16896 9998
rect 17052 9994 17080 10746
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 17236 9654 17264 10202
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16776 9178 16804 9454
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16868 9042 16896 9454
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16120 8502 16172 8508
rect 16578 8528 16634 8537
rect 16132 8430 16160 8502
rect 16578 8463 16634 8472
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 14752 7750 14780 8366
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 15028 7478 15056 7822
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 5778 14044 7142
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 15212 4146 15240 7958
rect 16868 5778 16896 8978
rect 17236 8922 17264 9590
rect 17144 8894 17264 8922
rect 17144 8498 17172 8894
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8634 17264 8774
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17328 8566 17356 11018
rect 17420 9178 17448 11630
rect 17512 10674 17540 12650
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17682 12336 17738 12345
rect 17682 12271 17738 12280
rect 17696 11082 17724 12271
rect 17880 11898 17908 12582
rect 17972 12442 18000 12786
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18432 12345 18460 12718
rect 18418 12336 18474 12345
rect 18418 12271 18474 12280
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18432 11694 18460 12038
rect 18524 11898 18552 14719
rect 18616 11898 18644 14742
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18708 13297 18736 14554
rect 18694 13288 18750 13297
rect 18694 13223 18750 13232
rect 18892 13002 18920 17326
rect 18970 17232 19026 17241
rect 18970 17167 19026 17176
rect 18984 14958 19012 17167
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18984 14074 19012 14758
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 18708 12974 18920 13002
rect 18708 12102 18736 12974
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18800 11778 18828 12242
rect 18892 12102 18920 12854
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18800 11750 18920 11778
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18708 11218 18736 11630
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18800 10713 18828 11630
rect 18892 11082 18920 11750
rect 18984 11354 19012 13466
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18786 10704 18842 10713
rect 17500 10668 17552 10674
rect 18892 10674 18920 11018
rect 18786 10639 18842 10648
rect 18880 10668 18932 10674
rect 17500 10610 17552 10616
rect 18880 10610 18932 10616
rect 18892 9994 18920 10610
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18892 9654 18920 9930
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18892 9178 18920 9590
rect 19076 9450 19104 19314
rect 19168 16114 19196 22374
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19168 14385 19196 15302
rect 19154 14376 19210 14385
rect 19154 14311 19210 14320
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19168 13530 19196 13670
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19168 12442 19196 12922
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19260 12186 19288 22578
rect 19444 22098 19472 22578
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19352 19990 19380 21830
rect 19444 21350 19472 22034
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 20942 19472 21286
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20602 19472 20878
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19338 19544 19394 19553
rect 19444 19514 19472 19858
rect 19338 19479 19394 19488
rect 19432 19508 19484 19514
rect 19352 19446 19380 19479
rect 19432 19450 19484 19456
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19536 18714 19564 22743
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 21010 19748 21286
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 19922 19656 20266
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19720 19310 19748 19790
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19720 18834 19748 19246
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19536 18686 19656 18714
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 18290 19380 18566
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 16425 19380 16458
rect 19338 16416 19394 16425
rect 19338 16351 19394 16360
rect 19444 15570 19472 16526
rect 19628 15706 19656 18686
rect 19706 17640 19762 17649
rect 19706 17575 19762 17584
rect 19720 17134 19748 17575
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19720 16114 19748 16730
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19338 14920 19394 14929
rect 19338 14855 19394 14864
rect 19352 14822 19380 14855
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19168 12158 19288 12186
rect 19168 11626 19196 12158
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19260 11150 19288 12038
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 19260 8090 19288 9930
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 12084 800 12112 2450
rect 12452 2446 12480 2858
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14752 800 14780 2450
rect 15028 2446 15056 3878
rect 15488 3126 15516 5102
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 17052 3058 17080 5510
rect 17420 4826 17448 5578
rect 17512 5234 17540 7142
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 19352 6186 19380 14758
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19444 14006 19472 14214
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 11762 19472 12582
rect 19536 12374 19564 14962
rect 19812 14890 19840 23054
rect 19904 20058 19932 24142
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23186 20116 23462
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20088 22710 20116 23122
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 20180 22438 20208 24006
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 20272 21962 20300 26200
rect 20916 24274 20944 26200
rect 21824 25628 21876 25634
rect 21824 25570 21876 25576
rect 21180 25560 21232 25566
rect 21180 25502 21232 25508
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21192 23798 21220 25502
rect 21180 23792 21232 23798
rect 21180 23734 21232 23740
rect 21362 23760 21418 23769
rect 20444 23724 20496 23730
rect 21362 23695 21418 23704
rect 20444 23666 20496 23672
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20364 22778 20392 22986
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20364 22030 20392 22374
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 19984 20868 20036 20874
rect 20088 20856 20116 20946
rect 20036 20828 20116 20856
rect 19984 20810 20036 20816
rect 19982 20496 20038 20505
rect 19982 20431 20038 20440
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19996 19786 20024 20431
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19720 11082 19748 11630
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 10606 19748 11018
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10130 19748 10542
rect 19812 10266 19840 14418
rect 19904 13977 19932 19654
rect 20088 19446 20116 19654
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19982 18456 20038 18465
rect 19982 18391 20038 18400
rect 19996 18290 20024 18391
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 20088 18222 20116 18634
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19996 15586 20024 18090
rect 20074 17912 20130 17921
rect 20074 17847 20130 17856
rect 20088 17814 20116 17847
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 20088 17270 20116 17750
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20180 16522 20208 17138
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 19996 15558 20116 15586
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19996 14929 20024 15370
rect 20088 15337 20116 15558
rect 20168 15496 20220 15502
rect 20272 15484 20300 21354
rect 20456 17898 20484 23666
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20548 22574 20576 23462
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20626 22536 20682 22545
rect 20626 22471 20682 22480
rect 20640 21865 20668 22471
rect 20732 22438 20760 23122
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20626 21856 20682 21865
rect 20626 21791 20682 21800
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20824 21554 20852 21626
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 19922 20576 20742
rect 21008 20534 21036 20810
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20640 19310 20668 20334
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20732 19718 20760 19994
rect 21008 19786 21036 20470
rect 20996 19780 21048 19786
rect 21048 19740 21128 19768
rect 20996 19722 21048 19728
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20220 15456 20300 15484
rect 20364 17870 20484 17898
rect 20168 15438 20220 15444
rect 20074 15328 20130 15337
rect 20074 15263 20130 15272
rect 19982 14920 20038 14929
rect 19982 14855 20038 14864
rect 19890 13968 19946 13977
rect 19890 13903 19946 13912
rect 19996 13326 20024 14855
rect 20364 13870 20392 17870
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20456 16658 20484 17682
rect 20626 17232 20682 17241
rect 20626 17167 20682 17176
rect 20640 17134 20668 17167
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20732 17082 20760 19654
rect 21100 19378 21128 19740
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20996 19236 21048 19242
rect 20996 19178 21048 19184
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20824 18204 20852 18566
rect 21008 18358 21036 19178
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21100 18426 21128 18838
rect 21192 18426 21220 19110
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 20996 18216 21048 18222
rect 20824 18176 20996 18204
rect 20996 18158 21048 18164
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20916 17202 20944 17614
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20732 17054 20944 17082
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20732 16658 20760 16934
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 15026 20668 15506
rect 20732 15094 20760 16390
rect 20824 16250 20852 16934
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20916 14414 20944 17054
rect 21008 15570 21036 18158
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21086 17232 21142 17241
rect 21086 17167 21088 17176
rect 21140 17167 21142 17176
rect 21088 17138 21140 17144
rect 21192 16794 21220 17478
rect 21284 17066 21312 17546
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21270 16688 21326 16697
rect 21270 16623 21326 16632
rect 21284 16250 21312 16623
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21270 16144 21326 16153
rect 21270 16079 21326 16088
rect 21284 16046 21312 16079
rect 21376 16046 21404 23695
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21652 23050 21680 23462
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21640 23044 21692 23050
rect 21640 22986 21692 22992
rect 21652 22710 21680 22986
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 21652 21690 21680 22646
rect 21744 22574 21772 23054
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21744 22166 21772 22510
rect 21836 22166 21864 25570
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 21928 24206 21956 24754
rect 22020 24290 22048 26302
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26330 24822 27000
rect 25410 26330 25466 27000
rect 26054 26330 26110 27000
rect 24504 26302 24822 26330
rect 22020 24274 22140 24290
rect 22020 24268 22152 24274
rect 22020 24262 22100 24268
rect 22100 24210 22152 24216
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 22204 22953 22232 26200
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22558 23624 22614 23633
rect 22296 22982 22324 23598
rect 22558 23559 22614 23568
rect 22284 22976 22336 22982
rect 22190 22944 22246 22953
rect 22284 22918 22336 22924
rect 22190 22879 22246 22888
rect 22466 22536 22522 22545
rect 22466 22471 22522 22480
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 21744 21690 21772 22102
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21652 21078 21680 21626
rect 21640 21072 21692 21078
rect 21640 21014 21692 21020
rect 21652 20874 21680 21014
rect 21640 20868 21692 20874
rect 21640 20810 21692 20816
rect 22204 20618 22232 21830
rect 22296 21146 22324 22102
rect 22480 21554 22508 22471
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22284 20800 22336 20806
rect 22388 20777 22416 20810
rect 22284 20742 22336 20748
rect 22374 20768 22430 20777
rect 21928 20590 22232 20618
rect 21928 20534 21956 20590
rect 21916 20528 21968 20534
rect 21916 20470 21968 20476
rect 21548 19916 21600 19922
rect 21468 19876 21548 19904
rect 21468 18834 21496 19876
rect 21548 19858 21600 19864
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21454 17368 21510 17377
rect 21454 17303 21456 17312
rect 21508 17303 21510 17312
rect 21456 17274 21508 17280
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20168 13728 20220 13734
rect 20088 13688 20168 13716
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20088 12918 20116 13688
rect 20168 13670 20220 13676
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20088 12306 20116 12718
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20364 12170 20392 13126
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19444 5846 19472 9114
rect 20364 8430 20392 12106
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 20456 8362 20484 13874
rect 20548 10470 20576 14214
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20732 12442 20760 13738
rect 20916 12986 20944 14214
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 21008 11354 21036 15506
rect 21468 15366 21496 16458
rect 21560 15745 21588 19314
rect 21744 18698 21772 19382
rect 22112 19174 22140 20590
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22020 18970 22048 19110
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 21744 18290 21772 18634
rect 21732 18284 21784 18290
rect 21732 18226 21784 18232
rect 21744 17678 21772 18226
rect 21836 17814 21864 18770
rect 22112 18630 22140 19110
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21640 17536 21692 17542
rect 21640 17478 21692 17484
rect 21652 17270 21680 17478
rect 21640 17264 21692 17270
rect 21638 17232 21640 17241
rect 21692 17232 21694 17241
rect 21638 17167 21694 17176
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21546 15736 21602 15745
rect 21546 15671 21602 15680
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21652 14278 21680 17070
rect 21836 15994 21864 17750
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21744 15966 21864 15994
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21744 14550 21772 15966
rect 21928 15706 21956 15982
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 14890 21956 15302
rect 22020 15026 22048 17614
rect 22112 15162 22140 18566
rect 22296 17218 22324 20742
rect 22374 20703 22430 20712
rect 22388 19854 22416 20703
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22204 17190 22324 17218
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21928 14346 21956 14826
rect 22020 14482 22048 14962
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 21100 12866 21128 13194
rect 21192 12986 21220 14010
rect 21836 13938 21864 14282
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21652 13462 21680 13874
rect 21836 13734 21864 13874
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 22204 13546 22232 17190
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22296 14929 22324 16662
rect 22282 14920 22338 14929
rect 22282 14855 22338 14864
rect 22388 14618 22416 19654
rect 22468 18896 22520 18902
rect 22466 18864 22468 18873
rect 22520 18864 22522 18873
rect 22466 18799 22522 18808
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22374 14376 22430 14385
rect 22374 14311 22430 14320
rect 22388 13938 22416 14311
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22112 13518 22232 13546
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21284 12866 21312 12922
rect 21100 12838 21312 12866
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21468 11558 21496 12718
rect 21928 12170 21956 12922
rect 22112 12889 22140 13518
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22098 12880 22154 12889
rect 22204 12850 22232 13330
rect 22388 13326 22416 13874
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22480 12918 22508 16390
rect 22572 16114 22600 23559
rect 22664 22094 22692 24754
rect 22848 23633 22876 26200
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22834 23624 22890 23633
rect 22834 23559 22890 23568
rect 23492 23508 23520 26200
rect 24136 24614 24164 26200
rect 24124 24608 24176 24614
rect 24124 24550 24176 24556
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 22848 23480 23520 23508
rect 22742 23352 22798 23361
rect 22848 23338 22876 23480
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22798 23310 22876 23338
rect 23296 23316 23348 23322
rect 22742 23287 22798 23296
rect 23296 23258 23348 23264
rect 23308 23225 23336 23258
rect 23110 23216 23166 23225
rect 23110 23151 23166 23160
rect 23294 23216 23350 23225
rect 23294 23151 23350 23160
rect 23124 22953 23152 23151
rect 23388 22976 23440 22982
rect 23110 22944 23166 22953
rect 23388 22918 23440 22924
rect 23110 22879 23166 22888
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22848 22216 22876 22578
rect 23400 22574 23428 22918
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23400 22234 23428 22510
rect 23584 22438 23612 24142
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23952 23866 23980 24074
rect 23940 23860 23992 23866
rect 23940 23802 23992 23808
rect 23664 23792 23716 23798
rect 23664 23734 23716 23740
rect 23676 23118 23704 23734
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 23254 23796 23462
rect 23848 23316 23900 23322
rect 23848 23258 23900 23264
rect 23756 23248 23808 23254
rect 23756 23190 23808 23196
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23676 22710 23704 23054
rect 23664 22704 23716 22710
rect 23716 22664 23796 22692
rect 23664 22646 23716 22652
rect 23768 22574 23796 22664
rect 23756 22568 23808 22574
rect 23756 22510 23808 22516
rect 23572 22432 23624 22438
rect 23572 22374 23624 22380
rect 23388 22228 23440 22234
rect 22848 22188 22968 22216
rect 22664 22066 22876 22094
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22756 21298 22784 21354
rect 22664 21270 22784 21298
rect 22664 21010 22692 21270
rect 22742 21176 22798 21185
rect 22742 21111 22798 21120
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22664 19446 22692 20742
rect 22756 20262 22784 21111
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22664 18970 22692 19246
rect 22742 19000 22798 19009
rect 22652 18964 22704 18970
rect 22742 18935 22798 18944
rect 22652 18906 22704 18912
rect 22756 18601 22784 18935
rect 22742 18592 22798 18601
rect 22742 18527 22798 18536
rect 22848 18358 22876 22066
rect 22940 21962 22968 22188
rect 23388 22170 23440 22176
rect 23572 22092 23624 22098
rect 23860 22094 23888 23258
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23572 22034 23624 22040
rect 23768 22066 23888 22094
rect 22928 21956 22980 21962
rect 22928 21898 22980 21904
rect 23296 21888 23348 21894
rect 23294 21856 23296 21865
rect 23584 21865 23612 22034
rect 23348 21856 23350 21865
rect 23294 21791 23350 21800
rect 23570 21856 23626 21865
rect 23570 21791 23626 21800
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23400 21554 23428 21626
rect 23572 21616 23624 21622
rect 23768 21604 23796 22066
rect 23952 21622 23980 22374
rect 23624 21576 23796 21604
rect 23940 21616 23992 21622
rect 23572 21558 23624 21564
rect 24044 21604 24072 22510
rect 24136 21706 24164 22918
rect 24308 22160 24360 22166
rect 24308 22102 24360 22108
rect 24136 21678 24256 21706
rect 24124 21616 24176 21622
rect 24044 21576 24124 21604
rect 23940 21558 23992 21564
rect 24124 21558 24176 21564
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23400 21026 23428 21490
rect 23478 21312 23534 21321
rect 23478 21247 23534 21256
rect 23492 21078 23520 21247
rect 23756 21140 23808 21146
rect 23676 21100 23756 21128
rect 23216 20998 23428 21026
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23572 21004 23624 21010
rect 23216 20466 23244 20998
rect 23572 20946 23624 20952
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 23308 20641 23336 20878
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23294 20632 23350 20641
rect 23400 20602 23428 20810
rect 23294 20567 23350 20576
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23584 19786 23612 20946
rect 23676 20806 23704 21100
rect 23756 21082 23808 21088
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23572 19780 23624 19786
rect 23572 19722 23624 19728
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23308 19514 23336 19654
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22848 18222 22876 18294
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22848 17202 22876 18158
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22664 15994 22692 16934
rect 22848 16810 22876 17138
rect 23216 17082 23244 17546
rect 23308 17270 23336 18906
rect 23400 18358 23428 19110
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23296 17264 23348 17270
rect 23296 17206 23348 17212
rect 23400 17082 23428 18294
rect 23216 17054 23428 17082
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22572 15966 22692 15994
rect 22756 16782 22876 16810
rect 22572 15094 22600 15966
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22560 15088 22612 15094
rect 22560 15030 22612 15036
rect 22572 13530 22600 15030
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22468 12912 22520 12918
rect 22468 12854 22520 12860
rect 22098 12815 22154 12824
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22204 12238 22232 12786
rect 22664 12782 22692 15846
rect 22756 14385 22784 16782
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22742 14376 22798 14385
rect 22742 14311 22798 14320
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 21916 12164 21968 12170
rect 21916 12106 21968 12112
rect 21928 11830 21956 12106
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9738 20760 9998
rect 21192 9926 21220 11018
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 10538 21404 10950
rect 21468 10810 21496 11494
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21560 10266 21588 10678
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21560 10062 21588 10202
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21652 9994 21680 11494
rect 21928 11082 21956 11766
rect 22204 11694 22232 12174
rect 22756 11830 22784 14214
rect 22848 13870 22876 16594
rect 23308 16590 23336 16934
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22940 15162 22968 15438
rect 23400 15366 23428 17054
rect 23492 16046 23520 19382
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23584 18766 23612 19110
rect 23676 18834 23704 19654
rect 23768 19378 23796 20742
rect 23860 19922 23888 20946
rect 24228 20913 24256 21678
rect 24214 20904 24270 20913
rect 24214 20839 24270 20848
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23860 19310 23888 19654
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23860 18630 23888 18702
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 23860 18358 23888 18566
rect 24044 18465 24072 18566
rect 24030 18456 24086 18465
rect 24030 18391 24086 18400
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 24044 17649 24072 18391
rect 24030 17640 24086 17649
rect 24030 17575 24086 17584
rect 24044 17270 24072 17575
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 23846 16688 23902 16697
rect 23846 16623 23902 16632
rect 23860 16522 23888 16623
rect 24136 16522 24164 19314
rect 24320 17814 24348 22102
rect 24412 21690 24440 23598
rect 24504 22953 24532 26302
rect 24766 26200 24822 26302
rect 24964 26302 25466 26330
rect 24964 24290 24992 26302
rect 25410 26200 25466 26302
rect 25700 26302 26110 26330
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24780 24262 24992 24290
rect 25056 24274 25084 24686
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25240 24274 25268 24550
rect 25044 24268 25096 24274
rect 24780 24206 24808 24262
rect 25044 24210 25096 24216
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24490 22944 24546 22953
rect 24490 22879 24546 22888
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24412 21078 24440 21626
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 24308 17808 24360 17814
rect 24308 17750 24360 17756
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24412 17338 24440 17478
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24308 17264 24360 17270
rect 24308 17206 24360 17212
rect 24320 16590 24348 17206
rect 24504 17134 24532 17682
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22848 12986 22876 13806
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 13530 23336 15098
rect 23400 15026 23428 15302
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23662 14920 23718 14929
rect 23386 14376 23442 14385
rect 23584 14346 23612 14894
rect 23662 14855 23664 14864
rect 23716 14855 23718 14864
rect 23664 14826 23716 14832
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23386 14311 23442 14320
rect 23572 14340 23624 14346
rect 23400 13938 23428 14311
rect 23572 14282 23624 14288
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23308 13274 23336 13466
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 23032 12850 23060 13262
rect 23308 13258 23428 13274
rect 23308 13252 23440 13258
rect 23308 13246 23388 13252
rect 23388 13194 23440 13200
rect 23112 13184 23164 13190
rect 23492 13138 23520 13330
rect 23164 13132 23520 13138
rect 23112 13126 23520 13132
rect 23124 13110 23520 13126
rect 23492 12986 23520 13110
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21928 10810 21956 11018
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 20640 9710 20760 9738
rect 20640 9586 20668 9710
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 21192 9518 21220 9862
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 22204 7410 22232 11630
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11354 23336 12922
rect 23584 12918 23612 14282
rect 23572 12912 23624 12918
rect 23572 12854 23624 12860
rect 23584 12434 23612 12854
rect 23676 12782 23704 14486
rect 23768 13462 23796 16390
rect 23860 16046 23888 16458
rect 24320 16114 24348 16526
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23860 15706 23888 15982
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23952 15026 23980 15370
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23952 14482 23980 14962
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 24044 13870 24072 15982
rect 24596 15586 24624 24006
rect 24964 23866 24992 24006
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24766 23488 24822 23497
rect 24766 23423 24822 23432
rect 24676 22976 24728 22982
rect 24676 22918 24728 22924
rect 24688 22710 24716 22918
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 24688 22030 24716 22646
rect 24780 22098 24808 23423
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25148 22778 25176 23122
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25318 22536 25374 22545
rect 25318 22471 25374 22480
rect 25332 22438 25360 22471
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 24768 22092 24820 22098
rect 24768 22034 24820 22040
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 24964 21865 24992 21898
rect 24950 21856 25006 21865
rect 24950 21791 25006 21800
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24688 20398 24716 21422
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 24964 19854 24992 20538
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24766 18592 24822 18601
rect 24766 18527 24822 18536
rect 24780 18358 24808 18527
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24688 17746 24716 18022
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 17202 24716 17682
rect 24780 17338 24808 18294
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24872 17218 24900 19246
rect 24676 17196 24728 17202
rect 24872 17190 24992 17218
rect 24728 17156 24808 17184
rect 24676 17138 24728 17144
rect 24780 17116 24808 17156
rect 24780 17088 24900 17116
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24688 16114 24716 16934
rect 24766 16144 24822 16153
rect 24676 16108 24728 16114
rect 24872 16114 24900 17088
rect 24964 16250 24992 17190
rect 25056 16590 25084 19654
rect 25134 19000 25190 19009
rect 25134 18935 25190 18944
rect 25148 16998 25176 18935
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24766 16079 24822 16088
rect 24860 16108 24912 16114
rect 24676 16050 24728 16056
rect 24688 15706 24716 16050
rect 24780 16046 24808 16079
rect 24860 16050 24912 16056
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24504 15558 24624 15586
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23860 13462 23888 13806
rect 23756 13456 23808 13462
rect 23756 13398 23808 13404
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12434 23704 12582
rect 23584 12406 23704 12434
rect 23676 12238 23704 12406
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 23952 11830 23980 12174
rect 24044 12102 24072 13806
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 24044 11694 24072 12038
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 22664 10606 22692 11290
rect 24308 11280 24360 11286
rect 24308 11222 24360 11228
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23400 7750 23428 9454
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21744 5846 21772 6734
rect 22480 5914 22508 7278
rect 22848 6458 22876 7686
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23768 6934 23796 9522
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23952 7002 23980 7482
rect 24320 7478 24348 11222
rect 24504 9722 24532 15558
rect 24964 15162 24992 16186
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 25056 14906 25084 16390
rect 24872 14890 25084 14906
rect 24860 14884 25084 14890
rect 24912 14878 25084 14884
rect 24860 14826 24912 14832
rect 24952 14340 25004 14346
rect 25056 14328 25084 14878
rect 25148 14346 25176 16594
rect 25240 16182 25268 21286
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25332 19446 25360 20946
rect 25516 20602 25544 22578
rect 25700 22438 25728 26302
rect 26054 26200 26110 26302
rect 26698 26330 26754 27000
rect 26698 26302 27016 26330
rect 26698 26200 26754 26302
rect 26424 25356 26476 25362
rect 26424 25298 26476 25304
rect 25964 24676 26016 24682
rect 25964 24618 26016 24624
rect 25976 24138 26004 24618
rect 26146 24168 26202 24177
rect 25964 24132 26016 24138
rect 26202 24126 26280 24154
rect 26436 24138 26464 25298
rect 26988 24410 27016 26302
rect 27342 26200 27398 27000
rect 27986 26200 28042 27000
rect 28630 26200 28686 27000
rect 29274 26330 29330 27000
rect 29274 26302 29592 26330
rect 29274 26200 29330 26302
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 27356 24342 27384 26200
rect 27710 25256 27766 25265
rect 27710 25191 27766 25200
rect 27528 24676 27580 24682
rect 27528 24618 27580 24624
rect 27344 24336 27396 24342
rect 27344 24278 27396 24284
rect 26146 24103 26202 24112
rect 25964 24074 26016 24080
rect 26252 24070 26280 24126
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 25872 24064 25924 24070
rect 25792 24012 25872 24018
rect 25792 24006 25924 24012
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26332 24064 26384 24070
rect 26332 24006 26384 24012
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 25792 23990 25912 24006
rect 25792 22964 25820 23990
rect 26344 23769 26372 24006
rect 26424 23792 26476 23798
rect 26330 23760 26386 23769
rect 26424 23734 26476 23740
rect 26330 23695 26386 23704
rect 25872 23656 25924 23662
rect 25924 23604 26280 23610
rect 25872 23598 26280 23604
rect 25884 23582 26280 23598
rect 25872 22976 25924 22982
rect 25792 22936 25872 22964
rect 25872 22918 25924 22924
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25778 22400 25834 22409
rect 25778 22335 25834 22344
rect 25792 22030 25820 22335
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25700 21350 25728 21830
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25792 21078 25820 21966
rect 25884 21418 25912 22918
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 26068 22234 26096 22442
rect 26252 22234 26280 23582
rect 26332 23588 26384 23594
rect 26332 23530 26384 23536
rect 26344 22778 26372 23530
rect 26436 22778 26464 23734
rect 27160 23656 27212 23662
rect 27212 23616 27292 23644
rect 27160 23598 27212 23604
rect 26608 23520 26660 23526
rect 26606 23488 26608 23497
rect 26660 23488 26662 23497
rect 26606 23423 26662 23432
rect 27264 23186 27292 23616
rect 27252 23180 27304 23186
rect 27252 23122 27304 23128
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 26976 22976 27028 22982
rect 26976 22918 27028 22924
rect 26332 22772 26384 22778
rect 26332 22714 26384 22720
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26056 22228 26108 22234
rect 26056 22170 26108 22176
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 26068 21962 26096 22034
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 26436 21944 26464 22714
rect 26804 22710 26832 22918
rect 26608 22704 26660 22710
rect 26608 22646 26660 22652
rect 26792 22704 26844 22710
rect 26792 22646 26844 22652
rect 26516 21956 26568 21962
rect 26436 21916 26516 21944
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25976 21690 26004 21830
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 26068 21418 26096 21898
rect 25872 21412 25924 21418
rect 25872 21354 25924 21360
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 26056 21140 26108 21146
rect 26108 21100 26372 21128
rect 26056 21082 26108 21088
rect 25780 21072 25832 21078
rect 25780 21014 25832 21020
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 26068 20602 26096 20946
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 25688 20324 25740 20330
rect 25688 20266 25740 20272
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25320 19440 25372 19446
rect 25320 19382 25372 19388
rect 25320 19236 25372 19242
rect 25320 19178 25372 19184
rect 25412 19236 25464 19242
rect 25412 19178 25464 19184
rect 25332 18358 25360 19178
rect 25424 18970 25452 19178
rect 25516 18970 25544 19722
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25700 18698 25728 20266
rect 25962 20088 26018 20097
rect 25962 20023 26018 20032
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25792 19310 25820 19790
rect 25976 19553 26004 20023
rect 25962 19544 26018 19553
rect 25962 19479 26018 19488
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25792 18834 25820 19246
rect 25870 18864 25926 18873
rect 25780 18828 25832 18834
rect 25870 18799 25926 18808
rect 25780 18770 25832 18776
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25410 17912 25466 17921
rect 25410 17847 25466 17856
rect 25424 17610 25452 17847
rect 25792 17746 25820 18770
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25412 17604 25464 17610
rect 25412 17546 25464 17552
rect 25884 16726 25912 18799
rect 25976 16726 26004 19479
rect 26068 18358 26096 20538
rect 26148 19916 26200 19922
rect 26148 19858 26200 19864
rect 26160 19258 26188 19858
rect 26252 19514 26280 20810
rect 26344 20466 26372 21100
rect 26436 20874 26464 21916
rect 26516 21898 26568 21904
rect 26620 21690 26648 22646
rect 26988 22642 27016 22918
rect 27158 22808 27214 22817
rect 27158 22743 27214 22752
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 26988 22545 27016 22578
rect 26974 22536 27030 22545
rect 26974 22471 27030 22480
rect 27172 22273 27200 22743
rect 27264 22574 27292 23122
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27264 22409 27292 22510
rect 27250 22400 27306 22409
rect 27250 22335 27306 22344
rect 27158 22264 27214 22273
rect 27158 22199 27214 22208
rect 27252 22160 27304 22166
rect 27252 22102 27304 22108
rect 27066 21720 27122 21729
rect 26608 21684 26660 21690
rect 27066 21655 27122 21664
rect 26608 21626 26660 21632
rect 26516 21548 26568 21554
rect 26516 21490 26568 21496
rect 26528 21146 26556 21490
rect 26516 21140 26568 21146
rect 26516 21082 26568 21088
rect 27080 21049 27108 21655
rect 27264 21321 27292 22102
rect 27250 21312 27306 21321
rect 27250 21247 27306 21256
rect 27066 21040 27122 21049
rect 27066 20975 27122 20984
rect 26424 20868 26476 20874
rect 26424 20810 26476 20816
rect 26436 20534 26464 20810
rect 27066 20632 27122 20641
rect 27066 20567 27068 20576
rect 27120 20567 27122 20576
rect 27068 20538 27120 20544
rect 26424 20528 26476 20534
rect 26424 20470 26476 20476
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26436 19786 26464 20470
rect 27356 20466 27384 24006
rect 27436 23656 27488 23662
rect 27436 23598 27488 23604
rect 27448 23361 27476 23598
rect 27434 23352 27490 23361
rect 27434 23287 27490 23296
rect 27540 22778 27568 24618
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27528 22500 27580 22506
rect 27528 22442 27580 22448
rect 27540 22234 27568 22442
rect 27528 22228 27580 22234
rect 27528 22170 27580 22176
rect 27526 22128 27582 22137
rect 27526 22063 27582 22072
rect 27540 21321 27568 22063
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27632 21350 27660 21626
rect 27620 21344 27672 21350
rect 27526 21312 27582 21321
rect 27620 21286 27672 21292
rect 27526 21247 27582 21256
rect 27724 21010 27752 25191
rect 28000 24206 28028 26200
rect 28448 25492 28500 25498
rect 28448 25434 28500 25440
rect 28460 24290 28488 25434
rect 28644 24818 28672 26200
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28552 24698 28580 24754
rect 28552 24670 29132 24698
rect 29104 24614 29132 24670
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 28460 24262 28764 24290
rect 27988 24200 28040 24206
rect 27988 24142 28040 24148
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 28368 22710 28396 24006
rect 28460 23866 28488 24142
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28630 23624 28686 23633
rect 28540 23588 28592 23594
rect 28630 23559 28686 23568
rect 28540 23530 28592 23536
rect 28552 23322 28580 23530
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28538 22808 28594 22817
rect 28538 22743 28594 22752
rect 28552 22710 28580 22743
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28540 22704 28592 22710
rect 28540 22646 28592 22652
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28368 22438 28396 22510
rect 28264 22432 28316 22438
rect 28264 22374 28316 22380
rect 28356 22432 28408 22438
rect 28356 22374 28408 22380
rect 28276 22166 28304 22374
rect 28264 22160 28316 22166
rect 28264 22102 28316 22108
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28368 21486 28396 22374
rect 28448 22092 28500 22098
rect 28448 22034 28500 22040
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 27816 21078 27844 21422
rect 27896 21412 27948 21418
rect 27896 21354 27948 21360
rect 27804 21072 27856 21078
rect 27804 21014 27856 21020
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 27158 20224 27214 20233
rect 26528 19922 26556 20198
rect 27158 20159 27214 20168
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26424 19780 26476 19786
rect 26424 19722 26476 19728
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26620 19334 26648 19722
rect 26620 19306 26832 19334
rect 27172 19310 27200 20159
rect 27356 19378 27384 20402
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 27632 19689 27660 19858
rect 27618 19680 27674 19689
rect 27618 19615 27674 19624
rect 27724 19514 27752 20198
rect 27816 20058 27844 21014
rect 27908 20806 27936 21354
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28368 20398 28396 21422
rect 28460 20942 28488 22034
rect 28644 22030 28672 23559
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28644 21865 28672 21966
rect 28736 21894 28764 24262
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28920 23186 28948 23462
rect 29012 23322 29040 24550
rect 29564 24410 29592 26302
rect 29918 26200 29974 27000
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26330 31906 27000
rect 31850 26302 31984 26330
rect 31850 26200 31906 26302
rect 29460 24404 29512 24410
rect 29460 24346 29512 24352
rect 29552 24404 29604 24410
rect 29552 24346 29604 24352
rect 29184 24064 29236 24070
rect 29184 24006 29236 24012
rect 29196 23866 29224 24006
rect 29184 23860 29236 23866
rect 29184 23802 29236 23808
rect 29472 23746 29500 24346
rect 29932 24138 29960 26200
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 30012 25016 30064 25022
rect 30012 24958 30064 24964
rect 29920 24132 29972 24138
rect 29920 24074 29972 24080
rect 29472 23730 29684 23746
rect 29460 23724 29684 23730
rect 29512 23718 29684 23724
rect 29460 23666 29512 23672
rect 29460 23588 29512 23594
rect 29460 23530 29512 23536
rect 29472 23322 29500 23530
rect 29000 23316 29052 23322
rect 29460 23316 29512 23322
rect 29000 23258 29052 23264
rect 29380 23276 29460 23304
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 29380 23118 29408 23276
rect 29460 23258 29512 23264
rect 29368 23112 29420 23118
rect 29368 23054 29420 23060
rect 29380 22710 29408 23054
rect 29368 22704 29420 22710
rect 29368 22646 29420 22652
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 28908 21956 28960 21962
rect 28908 21898 28960 21904
rect 28724 21888 28776 21894
rect 28630 21856 28686 21865
rect 28724 21830 28776 21836
rect 28630 21791 28686 21800
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28356 20256 28408 20262
rect 28356 20198 28408 20204
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27344 19372 27396 19378
rect 27816 19334 27844 19654
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28172 19440 28224 19446
rect 28368 19428 28396 20198
rect 28224 19400 28396 19428
rect 28172 19382 28224 19388
rect 27344 19314 27396 19320
rect 26160 19230 26280 19258
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 26252 18222 26280 19230
rect 26804 19174 26832 19306
rect 26976 19304 27028 19310
rect 26974 19272 26976 19281
rect 27160 19304 27212 19310
rect 27028 19272 27030 19281
rect 27160 19246 27212 19252
rect 27540 19306 27844 19334
rect 26974 19207 27030 19216
rect 27540 19174 27568 19306
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 26700 18896 26752 18902
rect 26700 18838 26752 18844
rect 26712 18426 26740 18838
rect 26804 18766 26832 19110
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 26700 18420 26752 18426
rect 26700 18362 26752 18368
rect 26240 18216 26292 18222
rect 26804 18170 26832 18702
rect 26240 18158 26292 18164
rect 26252 17882 26280 18158
rect 26712 18142 26832 18170
rect 27068 18216 27120 18222
rect 27632 18193 27660 18702
rect 27068 18158 27120 18164
rect 27618 18184 27674 18193
rect 26712 18086 26740 18142
rect 26700 18080 26752 18086
rect 26700 18022 26752 18028
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26712 17610 26740 18022
rect 26700 17604 26752 17610
rect 26700 17546 26752 17552
rect 26712 17270 26740 17546
rect 26700 17264 26752 17270
rect 26700 17206 26752 17212
rect 26712 16998 26740 17206
rect 26700 16992 26752 16998
rect 26700 16934 26752 16940
rect 25872 16720 25924 16726
rect 25872 16662 25924 16668
rect 25964 16720 26016 16726
rect 25964 16662 26016 16668
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25228 16176 25280 16182
rect 25228 16118 25280 16124
rect 25792 15570 25820 16594
rect 25976 16454 26004 16662
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 26146 16416 26202 16425
rect 26146 16351 26202 16360
rect 26160 15978 26188 16351
rect 26712 16114 26740 16934
rect 27080 16658 27108 18158
rect 27618 18119 27674 18128
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27356 17882 27384 18022
rect 27434 17912 27490 17921
rect 27344 17876 27396 17882
rect 27434 17847 27436 17856
rect 27344 17818 27396 17824
rect 27488 17847 27490 17856
rect 27436 17818 27488 17824
rect 27724 17218 27752 18702
rect 28000 18612 28028 19246
rect 28184 19174 28212 19382
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 27816 18584 28028 18612
rect 27816 18290 27844 18584
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 28460 18306 28488 20878
rect 28736 20233 28764 21830
rect 28920 21146 28948 21898
rect 29012 21622 29040 22510
rect 29184 22094 29236 22098
rect 29380 22094 29408 22646
rect 29656 22506 29684 23718
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 29736 23112 29788 23118
rect 29840 23100 29868 23258
rect 29788 23072 29868 23100
rect 29736 23054 29788 23060
rect 29644 22500 29696 22506
rect 29644 22442 29696 22448
rect 29840 22438 29868 23072
rect 29920 23044 29972 23050
rect 29920 22986 29972 22992
rect 29932 22642 29960 22986
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 29828 22432 29880 22438
rect 29828 22374 29880 22380
rect 29840 22234 29868 22374
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 29184 22092 29408 22094
rect 29236 22066 29408 22092
rect 29472 22066 29684 22094
rect 29184 22034 29236 22040
rect 29196 21622 29224 22034
rect 29368 21888 29420 21894
rect 29472 21876 29500 22066
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29420 21848 29500 21876
rect 29564 21865 29592 21966
rect 29656 21962 29684 22066
rect 29644 21956 29696 21962
rect 29644 21898 29696 21904
rect 29550 21856 29606 21865
rect 29368 21830 29420 21836
rect 29550 21791 29606 21800
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 29184 21616 29236 21622
rect 29184 21558 29236 21564
rect 28908 21140 28960 21146
rect 28908 21082 28960 21088
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 28722 20224 28778 20233
rect 28722 20159 28778 20168
rect 29012 19961 29040 20742
rect 29092 20528 29144 20534
rect 29196 20516 29224 21558
rect 29826 21448 29882 21457
rect 29826 21383 29882 21392
rect 29736 21140 29788 21146
rect 29736 21082 29788 21088
rect 29144 20488 29224 20516
rect 29092 20470 29144 20476
rect 28998 19952 29054 19961
rect 28998 19887 29054 19896
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28644 18358 28672 19110
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 28368 18278 28488 18306
rect 28632 18352 28684 18358
rect 28632 18294 28684 18300
rect 27816 17746 27844 18226
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27632 17190 27752 17218
rect 27816 17202 27844 17682
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27804 17196 27856 17202
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27172 16658 27200 16934
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26148 15972 26200 15978
rect 26148 15914 26200 15920
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25004 14300 25084 14328
rect 25136 14340 25188 14346
rect 24952 14282 25004 14288
rect 25136 14282 25188 14288
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24596 14006 24624 14214
rect 25148 14006 25176 14282
rect 24584 14000 24636 14006
rect 25136 14000 25188 14006
rect 24584 13942 24636 13948
rect 25056 13948 25136 13954
rect 25056 13942 25188 13948
rect 25056 13926 25176 13942
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24492 9716 24544 9722
rect 24492 9658 24544 9664
rect 24596 9654 24624 13670
rect 25056 12170 25084 13926
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24688 11830 24716 12038
rect 24676 11824 24728 11830
rect 24676 11766 24728 11772
rect 24688 11558 24716 11766
rect 25148 11694 25176 13806
rect 25240 13190 25268 15302
rect 25608 15201 25636 15438
rect 25594 15192 25650 15201
rect 25594 15127 25650 15136
rect 25792 14550 25820 15506
rect 26252 15026 26280 16050
rect 27172 16046 27200 16594
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 26332 15632 26384 15638
rect 26332 15574 26384 15580
rect 26344 15366 26372 15574
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 25780 14544 25832 14550
rect 25780 14486 25832 14492
rect 26344 14346 26372 15302
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26620 14482 26648 14758
rect 26988 14618 27016 15438
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26988 14414 27016 14554
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25700 14006 25728 14214
rect 25792 14074 25820 14214
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 25228 13184 25280 13190
rect 25228 13126 25280 13132
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24688 11286 24716 11494
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 26896 11218 26924 13194
rect 27632 12434 27660 17190
rect 27804 17138 27856 17144
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27724 16590 27752 17070
rect 27712 16584 27764 16590
rect 28368 16561 28396 18278
rect 29012 17882 29040 19790
rect 29104 19718 29132 20470
rect 29748 20058 29776 21082
rect 29840 20942 29868 21383
rect 30024 21010 30052 24958
rect 30392 23526 30420 25094
rect 30576 25022 30604 26200
rect 30564 25016 30616 25022
rect 30564 24958 30616 24964
rect 30564 24744 30616 24750
rect 30564 24686 30616 24692
rect 30104 23520 30156 23526
rect 30104 23462 30156 23468
rect 30380 23520 30432 23526
rect 30380 23462 30432 23468
rect 30116 23322 30144 23462
rect 30104 23316 30156 23322
rect 30104 23258 30156 23264
rect 30576 22506 30604 24686
rect 31024 24404 31076 24410
rect 31024 24346 31076 24352
rect 30748 24336 30800 24342
rect 30748 24278 30800 24284
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 30668 23798 30696 24006
rect 30760 23798 30788 24278
rect 31036 24206 31064 24346
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 30656 23792 30708 23798
rect 30656 23734 30708 23740
rect 30748 23792 30800 23798
rect 30748 23734 30800 23740
rect 31024 23588 31076 23594
rect 31024 23530 31076 23536
rect 30748 23180 30800 23186
rect 30748 23122 30800 23128
rect 30760 22778 30788 23122
rect 31036 22778 31064 23530
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 31024 22772 31076 22778
rect 31024 22714 31076 22720
rect 30564 22500 30616 22506
rect 30564 22442 30616 22448
rect 30760 22098 30788 22714
rect 30840 22704 30892 22710
rect 30840 22646 30892 22652
rect 30748 22092 30800 22098
rect 30748 22034 30800 22040
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30392 21418 30420 21830
rect 30380 21412 30432 21418
rect 30380 21354 30432 21360
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 29920 21004 29972 21010
rect 29920 20946 29972 20952
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 30104 21004 30156 21010
rect 30104 20946 30156 20952
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29932 20244 29960 20946
rect 30116 20369 30144 20946
rect 30208 20398 30236 21286
rect 30196 20392 30248 20398
rect 30102 20360 30158 20369
rect 30196 20334 30248 20340
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30102 20295 30158 20304
rect 29932 20216 30236 20244
rect 29736 20052 29788 20058
rect 29736 19994 29788 20000
rect 29920 20052 29972 20058
rect 29920 19994 29972 20000
rect 29932 19854 29960 19994
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29828 19780 29880 19786
rect 29828 19722 29880 19728
rect 29092 19712 29144 19718
rect 29840 19689 29868 19722
rect 29092 19654 29144 19660
rect 29826 19680 29882 19689
rect 29104 19446 29132 19654
rect 29826 19615 29882 19624
rect 29092 19440 29144 19446
rect 29092 19382 29144 19388
rect 29104 18698 29132 19382
rect 29828 18828 29880 18834
rect 29828 18770 29880 18776
rect 29092 18692 29144 18698
rect 29092 18634 29144 18640
rect 29104 18358 29132 18634
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29736 18624 29788 18630
rect 29736 18566 29788 18572
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 29104 17882 29132 18294
rect 29656 18290 29684 18566
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29092 17876 29144 17882
rect 29092 17818 29144 17824
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 27712 16526 27764 16532
rect 28354 16552 28410 16561
rect 28460 16522 28488 17750
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 17338 28856 17478
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28816 16652 28868 16658
rect 29012 16640 29040 17818
rect 29104 17338 29132 17818
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 28868 16612 29040 16640
rect 28816 16594 28868 16600
rect 28354 16487 28410 16496
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 29748 15978 29776 18566
rect 29840 18086 29868 18770
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29736 15972 29788 15978
rect 29736 15914 29788 15920
rect 29932 15609 29960 19790
rect 30208 19718 30236 20216
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30116 18426 30144 18566
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30208 18306 30236 19654
rect 30300 19174 30328 20334
rect 30392 19514 30420 21354
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30668 20874 30696 21286
rect 30656 20868 30708 20874
rect 30656 20810 30708 20816
rect 30852 20602 30880 22646
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 31036 22545 31064 22578
rect 31022 22536 31078 22545
rect 31022 22471 31078 22480
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 31036 20330 31064 22471
rect 31220 22166 31248 26200
rect 31300 24676 31352 24682
rect 31300 24618 31352 24624
rect 31312 24410 31340 24618
rect 31300 24404 31352 24410
rect 31300 24346 31352 24352
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31404 22710 31432 24142
rect 31852 23520 31904 23526
rect 31852 23462 31904 23468
rect 31864 23322 31892 23462
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 31496 23050 31800 23066
rect 31484 23044 31800 23050
rect 31536 23038 31800 23044
rect 31484 22986 31536 22992
rect 31392 22704 31444 22710
rect 31392 22646 31444 22652
rect 31772 22642 31800 23038
rect 31760 22636 31812 22642
rect 31760 22578 31812 22584
rect 31864 22506 31892 23258
rect 31956 23186 31984 26302
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26200 33838 27000
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26330 37058 27000
rect 37002 26302 37228 26330
rect 37002 26200 37058 26302
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32036 24132 32088 24138
rect 32036 24074 32088 24080
rect 32048 23798 32076 24074
rect 32036 23792 32088 23798
rect 32036 23734 32088 23740
rect 32324 23730 32352 24754
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32232 23322 32260 23666
rect 32220 23316 32272 23322
rect 32220 23258 32272 23264
rect 31944 23180 31996 23186
rect 31944 23122 31996 23128
rect 32036 22976 32088 22982
rect 32036 22918 32088 22924
rect 32048 22817 32076 22918
rect 32034 22808 32090 22817
rect 31956 22766 32034 22794
rect 31852 22500 31904 22506
rect 31852 22442 31904 22448
rect 31956 22386 31984 22766
rect 32034 22743 32090 22752
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32036 22500 32088 22506
rect 32036 22442 32088 22448
rect 31772 22358 31984 22386
rect 31208 22160 31260 22166
rect 31208 22102 31260 22108
rect 31392 21956 31444 21962
rect 31392 21898 31444 21904
rect 31404 21418 31432 21898
rect 31772 21706 31800 22358
rect 31944 22228 31996 22234
rect 31944 22170 31996 22176
rect 31956 22137 31984 22170
rect 31942 22128 31998 22137
rect 32048 22098 32076 22442
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32140 22273 32168 22374
rect 32126 22264 32182 22273
rect 32126 22199 32182 22208
rect 32128 22160 32180 22166
rect 32128 22102 32180 22108
rect 31942 22063 31998 22072
rect 32036 22092 32088 22098
rect 31680 21678 31800 21706
rect 31392 21412 31444 21418
rect 31392 21354 31444 21360
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31024 20324 31076 20330
rect 31024 20266 31076 20272
rect 30564 20256 30616 20262
rect 30564 20198 30616 20204
rect 30932 20256 30984 20262
rect 30932 20198 30984 20204
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30484 18426 30512 19246
rect 30576 18766 30604 20198
rect 30838 20088 30894 20097
rect 30838 20023 30894 20032
rect 30748 19712 30800 19718
rect 30746 19680 30748 19689
rect 30800 19680 30802 19689
rect 30746 19615 30802 19624
rect 30852 19417 30880 20023
rect 30654 19408 30710 19417
rect 30654 19343 30656 19352
rect 30708 19343 30710 19352
rect 30838 19408 30894 19417
rect 30838 19343 30894 19352
rect 30656 19314 30708 19320
rect 30944 19174 30972 20198
rect 31024 20052 31076 20058
rect 31024 19994 31076 20000
rect 31036 19718 31064 19994
rect 31024 19712 31076 19718
rect 31024 19654 31076 19660
rect 31036 19446 31064 19654
rect 31024 19440 31076 19446
rect 31024 19382 31076 19388
rect 30932 19168 30984 19174
rect 30932 19110 30984 19116
rect 30564 18760 30616 18766
rect 30564 18702 30616 18708
rect 30944 18698 30972 19110
rect 30932 18692 30984 18698
rect 30932 18634 30984 18640
rect 30472 18420 30524 18426
rect 30472 18362 30524 18368
rect 30116 18278 30236 18306
rect 30116 16017 30144 18278
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30392 17814 30420 18090
rect 30380 17808 30432 17814
rect 30380 17750 30432 17756
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 30208 17649 30236 17682
rect 30194 17640 30250 17649
rect 30194 17575 30250 17584
rect 30208 17338 30236 17575
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30392 17134 30420 17750
rect 30748 17604 30800 17610
rect 30748 17546 30800 17552
rect 30760 17270 30788 17546
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30944 16794 30972 17478
rect 31220 17105 31248 20742
rect 31206 17096 31262 17105
rect 31206 17031 31262 17040
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 30102 16008 30158 16017
rect 30102 15943 30158 15952
rect 29918 15600 29974 15609
rect 29918 15535 29974 15544
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 31404 13433 31432 21354
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31588 20262 31616 21286
rect 31680 20602 31708 21678
rect 31760 21616 31812 21622
rect 31760 21558 31812 21564
rect 31852 21616 31904 21622
rect 31852 21558 31904 21564
rect 31772 20602 31800 21558
rect 31864 21146 31892 21558
rect 31852 21140 31904 21146
rect 31852 21082 31904 21088
rect 31668 20596 31720 20602
rect 31668 20538 31720 20544
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 31576 20256 31628 20262
rect 31680 20244 31708 20538
rect 31956 20466 31984 22063
rect 32036 22034 32088 22040
rect 32036 21956 32088 21962
rect 32036 21898 32088 21904
rect 32048 21350 32076 21898
rect 32140 21486 32168 22102
rect 32232 22098 32260 22578
rect 32220 22092 32272 22098
rect 32220 22034 32272 22040
rect 32324 21570 32352 23666
rect 32508 23254 32536 26200
rect 32864 25016 32916 25022
rect 32864 24958 32916 24964
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 32496 23248 32548 23254
rect 32496 23190 32548 23196
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32680 23112 32732 23118
rect 32680 23054 32732 23060
rect 32416 22137 32444 23054
rect 32588 22976 32640 22982
rect 32588 22918 32640 22924
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32402 22128 32458 22137
rect 32402 22063 32458 22072
rect 32232 21542 32352 21570
rect 32404 21548 32456 21554
rect 32128 21480 32180 21486
rect 32128 21422 32180 21428
rect 32036 21344 32088 21350
rect 32036 21286 32088 21292
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 32036 20868 32088 20874
rect 32036 20810 32088 20816
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 31944 20324 31996 20330
rect 31944 20266 31996 20272
rect 31760 20256 31812 20262
rect 31680 20216 31760 20244
rect 31576 20198 31628 20204
rect 31760 20198 31812 20204
rect 31390 13424 31446 13433
rect 31390 13359 31446 13368
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27632 12406 27752 12434
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 27632 7546 27660 11018
rect 27724 10169 27752 12406
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27710 10160 27766 10169
rect 27710 10095 27766 10104
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 31312 9654 31340 11086
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 28172 9580 28224 9586
rect 28224 9540 28304 9568
rect 28172 9522 28224 9528
rect 28276 9500 28304 9540
rect 28276 9472 28396 9500
rect 28368 9382 28396 9472
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23756 6928 23808 6934
rect 23756 6870 23808 6876
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 19432 5840 19484 5846
rect 19432 5782 19484 5788
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17420 2990 17448 4762
rect 17696 4486 17724 5102
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 3126 17724 4422
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17880 3058 17908 4966
rect 20272 4826 20300 5646
rect 23400 5642 23428 6598
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24872 5642 24900 6190
rect 30288 5772 30340 5778
rect 30288 5714 30340 5720
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 25780 5636 25832 5642
rect 25780 5578 25832 5584
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5234 21404 5510
rect 22204 5234 22232 5578
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20272 4622 20300 4762
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 20548 3058 20576 4966
rect 22756 4554 22784 4966
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 25516 3194 25544 5510
rect 25792 3602 25820 5578
rect 27172 5370 27200 5578
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 28816 5296 28868 5302
rect 28816 5238 28868 5244
rect 28828 4826 28856 5238
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 27540 3194 27568 4626
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 29656 3194 29684 5102
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 29644 3188 29696 3194
rect 29644 3130 29696 3136
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 17420 800 17448 2450
rect 17512 2446 17540 2790
rect 20088 2446 20116 2790
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 1170 20208 2450
rect 21928 2446 21956 2790
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 26252 2650 26280 2994
rect 28368 2650 28396 2994
rect 30300 2922 30328 5714
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 31404 3126 31432 5102
rect 31392 3120 31444 3126
rect 31392 3062 31444 3068
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 30288 2916 30340 2922
rect 30288 2858 30340 2864
rect 31036 2650 31064 2994
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 28356 2644 28408 2650
rect 28356 2586 28408 2592
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 31588 2514 31616 9318
rect 31772 3398 31800 20198
rect 31956 17882 31984 20266
rect 31944 17876 31996 17882
rect 31944 17818 31996 17824
rect 31956 17678 31984 17818
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 31956 16658 31984 17614
rect 31944 16652 31996 16658
rect 31944 16594 31996 16600
rect 31956 3670 31984 16594
rect 32048 15473 32076 20810
rect 32140 20777 32168 20878
rect 32126 20768 32182 20777
rect 32126 20703 32182 20712
rect 32232 20602 32260 21542
rect 32404 21490 32456 21496
rect 32416 21434 32444 21490
rect 32324 21418 32444 21434
rect 32312 21412 32444 21418
rect 32364 21406 32444 21412
rect 32312 21354 32364 21360
rect 32128 20596 32180 20602
rect 32128 20538 32180 20544
rect 32220 20596 32272 20602
rect 32220 20538 32272 20544
rect 32140 20262 32168 20538
rect 32128 20256 32180 20262
rect 32128 20198 32180 20204
rect 32034 15464 32090 15473
rect 32034 15399 32090 15408
rect 31944 3664 31996 3670
rect 31944 3606 31996 3612
rect 32140 3466 32168 20198
rect 32324 20097 32352 21354
rect 32404 21344 32456 21350
rect 32404 21286 32456 21292
rect 32310 20088 32366 20097
rect 32310 20023 32366 20032
rect 32416 11898 32444 21286
rect 32508 20262 32536 22578
rect 32600 22166 32628 22918
rect 32692 22166 32720 23054
rect 32588 22160 32640 22166
rect 32588 22102 32640 22108
rect 32680 22160 32732 22166
rect 32680 22102 32732 22108
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32600 21010 32628 21966
rect 32784 21554 32812 23462
rect 32876 23304 32904 24958
rect 33152 24664 33180 26200
rect 33600 25220 33652 25226
rect 33600 25162 33652 25168
rect 33416 25084 33468 25090
rect 33416 25026 33468 25032
rect 33152 24636 33364 24664
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 33336 24206 33364 24636
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32876 23276 33180 23304
rect 33152 23118 33180 23276
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32968 22778 32996 22918
rect 32956 22772 33008 22778
rect 32956 22714 33008 22720
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32678 21448 32734 21457
rect 32678 21383 32734 21392
rect 32692 21185 32720 21383
rect 32772 21344 32824 21350
rect 32770 21312 32772 21321
rect 32824 21312 32826 21321
rect 32770 21247 32826 21256
rect 32678 21176 32734 21185
rect 32678 21111 32734 21120
rect 32588 21004 32640 21010
rect 32588 20946 32640 20952
rect 32876 20777 32904 21966
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 33336 21146 33364 24142
rect 33428 22778 33456 25026
rect 33508 24064 33560 24070
rect 33508 24006 33560 24012
rect 33520 23798 33548 24006
rect 33508 23792 33560 23798
rect 33508 23734 33560 23740
rect 33508 23044 33560 23050
rect 33508 22986 33560 22992
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33428 21554 33456 22578
rect 33416 21548 33468 21554
rect 33416 21490 33468 21496
rect 33428 21457 33456 21490
rect 33414 21448 33470 21457
rect 33414 21383 33470 21392
rect 33324 21140 33376 21146
rect 33324 21082 33376 21088
rect 32862 20768 32918 20777
rect 32862 20703 32918 20712
rect 32496 20256 32548 20262
rect 32496 20198 32548 20204
rect 32404 11892 32456 11898
rect 32404 11834 32456 11840
rect 32508 8634 32536 20198
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 33520 17785 33548 22986
rect 33612 21894 33640 25162
rect 33690 24712 33746 24721
rect 33690 24647 33746 24656
rect 33704 23798 33732 24647
rect 33796 24342 33824 26200
rect 33968 25424 34020 25430
rect 33968 25366 34020 25372
rect 33874 25120 33930 25129
rect 33874 25055 33930 25064
rect 33784 24336 33836 24342
rect 33784 24278 33836 24284
rect 33692 23792 33744 23798
rect 33692 23734 33744 23740
rect 33888 23322 33916 25055
rect 33876 23316 33928 23322
rect 33876 23258 33928 23264
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 33600 21888 33652 21894
rect 33600 21830 33652 21836
rect 33888 21418 33916 23054
rect 33876 21412 33928 21418
rect 33876 21354 33928 21360
rect 33980 21350 34008 25366
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 34058 24848 34114 24857
rect 34058 24783 34114 24792
rect 34072 23526 34100 24783
rect 34152 24064 34204 24070
rect 34152 24006 34204 24012
rect 34060 23520 34112 23526
rect 34060 23462 34112 23468
rect 34164 23118 34192 24006
rect 34242 23216 34298 23225
rect 34242 23151 34298 23160
rect 34152 23112 34204 23118
rect 34152 23054 34204 23060
rect 34256 22642 34284 23151
rect 34244 22636 34296 22642
rect 34244 22578 34296 22584
rect 34348 22094 34376 25230
rect 34440 23746 34468 26200
rect 34796 24404 34848 24410
rect 34796 24346 34848 24352
rect 34808 23866 34836 24346
rect 35084 24206 35112 26200
rect 35532 24744 35584 24750
rect 35532 24686 35584 24692
rect 35544 24274 35572 24686
rect 35624 24336 35676 24342
rect 35624 24278 35676 24284
rect 35532 24268 35584 24274
rect 35532 24210 35584 24216
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 35636 24138 35664 24278
rect 35624 24132 35676 24138
rect 35624 24074 35676 24080
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34440 23730 34560 23746
rect 34440 23724 34572 23730
rect 34440 23718 34520 23724
rect 34520 23666 34572 23672
rect 34532 22778 34560 23666
rect 35440 23520 35492 23526
rect 35440 23462 35492 23468
rect 35452 23118 35480 23462
rect 35728 23118 35756 26200
rect 36174 24984 36230 24993
rect 36174 24919 36230 24928
rect 35992 24064 36044 24070
rect 35992 24006 36044 24012
rect 36004 23798 36032 24006
rect 36188 23798 36216 24919
rect 36372 24206 36400 26200
rect 36544 24880 36596 24886
rect 36544 24822 36596 24828
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 35992 23792 36044 23798
rect 35992 23734 36044 23740
rect 36176 23792 36228 23798
rect 36176 23734 36228 23740
rect 35440 23112 35492 23118
rect 35716 23112 35768 23118
rect 35440 23054 35492 23060
rect 35622 23080 35678 23089
rect 35716 23054 35768 23060
rect 35622 23015 35624 23024
rect 35676 23015 35678 23024
rect 35624 22986 35676 22992
rect 34520 22772 34572 22778
rect 34520 22714 34572 22720
rect 36556 22710 36584 24822
rect 37096 24336 37148 24342
rect 37096 24278 37148 24284
rect 37108 23730 37136 24278
rect 36820 23724 36872 23730
rect 36820 23666 36872 23672
rect 37096 23724 37148 23730
rect 37096 23666 37148 23672
rect 36832 23186 36860 23666
rect 37004 23520 37056 23526
rect 37004 23462 37056 23468
rect 36820 23180 36872 23186
rect 36820 23122 36872 23128
rect 36544 22704 36596 22710
rect 34518 22672 34574 22681
rect 36544 22646 36596 22652
rect 34518 22607 34520 22616
rect 34572 22607 34574 22616
rect 34704 22636 34756 22642
rect 34520 22578 34572 22584
rect 34704 22578 34756 22584
rect 35716 22636 35768 22642
rect 35716 22578 35768 22584
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34164 22066 34376 22094
rect 34060 22024 34112 22030
rect 34060 21966 34112 21972
rect 33968 21344 34020 21350
rect 33968 21286 34020 21292
rect 34072 20806 34100 21966
rect 34164 21010 34192 22066
rect 34532 21049 34560 22374
rect 34518 21040 34574 21049
rect 34152 21004 34204 21010
rect 34518 20975 34574 20984
rect 34152 20946 34204 20952
rect 34060 20800 34112 20806
rect 34060 20742 34112 20748
rect 33506 17776 33562 17785
rect 33506 17711 33562 17720
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 34072 15065 34100 20742
rect 34716 19514 34744 22578
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35452 22030 35480 22170
rect 35164 22024 35216 22030
rect 35070 21992 35126 22001
rect 34980 21956 35032 21962
rect 35164 21966 35216 21972
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 35070 21927 35126 21936
rect 34980 21898 35032 21904
rect 34992 21350 35020 21898
rect 35084 21894 35112 21927
rect 35072 21888 35124 21894
rect 35072 21830 35124 21836
rect 34980 21344 35032 21350
rect 34980 21286 35032 21292
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34058 15056 34114 15065
rect 34058 14991 34114 15000
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 34992 13938 35020 21286
rect 35176 20058 35204 21966
rect 35452 21622 35480 21966
rect 35624 21888 35676 21894
rect 35624 21830 35676 21836
rect 35636 21690 35664 21830
rect 35624 21684 35676 21690
rect 35624 21626 35676 21632
rect 35440 21616 35492 21622
rect 35440 21558 35492 21564
rect 35728 21078 35756 22578
rect 36452 21956 36504 21962
rect 36452 21898 36504 21904
rect 36268 21888 36320 21894
rect 36268 21830 36320 21836
rect 36280 21593 36308 21830
rect 36266 21584 36322 21593
rect 36266 21519 36322 21528
rect 35716 21072 35768 21078
rect 35716 21014 35768 21020
rect 36464 20505 36492 21898
rect 36450 20496 36506 20505
rect 36450 20431 36506 20440
rect 35164 20052 35216 20058
rect 35164 19994 35216 20000
rect 34980 13932 35032 13938
rect 34980 13874 35032 13880
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32128 3460 32180 3466
rect 32128 3402 32180 3408
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33612 3194 33640 3334
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33704 2650 33732 2994
rect 35176 2990 35204 19994
rect 37016 17338 37044 23462
rect 37108 23254 37136 23666
rect 37096 23248 37148 23254
rect 37096 23190 37148 23196
rect 37200 22094 37228 26302
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38290 26302 38516 26330
rect 38290 26200 38346 26302
rect 37372 24064 37424 24070
rect 37372 24006 37424 24012
rect 37200 22066 37320 22094
rect 37292 22030 37320 22066
rect 37280 22024 37332 22030
rect 37280 21966 37332 21972
rect 37384 21486 37412 24006
rect 37464 22976 37516 22982
rect 37464 22918 37516 22924
rect 37476 22778 37504 22918
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37660 22166 37688 26200
rect 38488 24206 38516 26302
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 40866 26200 40922 27000
rect 41510 26200 41566 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26330 43498 27000
rect 43442 26302 43852 26330
rect 43442 26200 43498 26302
rect 38658 24304 38714 24313
rect 38658 24239 38714 24248
rect 38476 24200 38528 24206
rect 38528 24160 38608 24188
rect 38476 24142 38528 24148
rect 38476 24064 38528 24070
rect 38476 24006 38528 24012
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38488 23798 38516 24006
rect 38476 23792 38528 23798
rect 38476 23734 38528 23740
rect 38580 23322 38608 24160
rect 38672 23798 38700 24239
rect 38948 24206 38976 26200
rect 39304 24948 39356 24954
rect 39304 24890 39356 24896
rect 38936 24200 38988 24206
rect 38936 24142 38988 24148
rect 39316 23866 39344 24890
rect 39304 23860 39356 23866
rect 39304 23802 39356 23808
rect 38660 23792 38712 23798
rect 38660 23734 38712 23740
rect 39592 23730 39620 26200
rect 40236 24206 40264 26200
rect 39948 24200 40000 24206
rect 39948 24142 40000 24148
rect 40224 24200 40276 24206
rect 40224 24142 40276 24148
rect 39960 23866 39988 24142
rect 40684 24064 40736 24070
rect 40684 24006 40736 24012
rect 39948 23860 40000 23866
rect 39948 23802 40000 23808
rect 40696 23798 40724 24006
rect 40684 23792 40736 23798
rect 40684 23734 40736 23740
rect 39580 23724 39632 23730
rect 39580 23666 39632 23672
rect 40592 23520 40644 23526
rect 40592 23462 40644 23468
rect 38568 23316 38620 23322
rect 38568 23258 38620 23264
rect 40604 23186 40632 23462
rect 40592 23180 40644 23186
rect 40592 23122 40644 23128
rect 40316 23112 40368 23118
rect 40316 23054 40368 23060
rect 38752 22976 38804 22982
rect 38752 22918 38804 22924
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37648 22160 37700 22166
rect 37648 22102 37700 22108
rect 38764 22098 38792 22918
rect 39580 22432 39632 22438
rect 39580 22374 39632 22380
rect 38752 22092 38804 22098
rect 38752 22034 38804 22040
rect 37464 21888 37516 21894
rect 37464 21830 37516 21836
rect 37556 21888 37608 21894
rect 37556 21830 37608 21836
rect 37372 21480 37424 21486
rect 37372 21422 37424 21428
rect 37476 20534 37504 21830
rect 37464 20528 37516 20534
rect 37464 20470 37516 20476
rect 37568 17610 37596 21830
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 39592 18154 39620 22374
rect 40328 21962 40356 23054
rect 40880 22778 40908 26200
rect 41524 24410 41552 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 41512 24404 41564 24410
rect 41512 24346 41564 24352
rect 42616 24404 42668 24410
rect 42616 24346 42668 24352
rect 41420 24064 41472 24070
rect 41420 24006 41472 24012
rect 40868 22772 40920 22778
rect 40868 22714 40920 22720
rect 41432 22642 41460 24006
rect 42628 23730 42656 24346
rect 43444 24336 43496 24342
rect 43444 24278 43496 24284
rect 43352 24132 43404 24138
rect 43352 24074 43404 24080
rect 42800 24064 42852 24070
rect 42800 24006 42852 24012
rect 42616 23724 42668 23730
rect 42616 23666 42668 23672
rect 42812 22642 42840 24006
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 43260 23112 43312 23118
rect 43260 23054 43312 23060
rect 43272 22778 43300 23054
rect 43260 22772 43312 22778
rect 43260 22714 43312 22720
rect 41420 22636 41472 22642
rect 41420 22578 41472 22584
rect 42800 22636 42852 22642
rect 42800 22578 42852 22584
rect 40684 22432 40736 22438
rect 40684 22374 40736 22380
rect 41328 22432 41380 22438
rect 41328 22374 41380 22380
rect 40316 21956 40368 21962
rect 40316 21898 40368 21904
rect 40696 20913 40724 22374
rect 40682 20904 40738 20913
rect 40682 20839 40738 20848
rect 41340 19854 41368 22374
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42800 22228 42852 22234
rect 42800 22170 42852 22176
rect 41328 19848 41380 19854
rect 41328 19790 41380 19796
rect 39580 18148 39632 18154
rect 39580 18090 39632 18096
rect 37556 17604 37608 17610
rect 37556 17546 37608 17552
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37004 17332 37056 17338
rect 37004 17274 37056 17280
rect 42812 16998 42840 22170
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 43364 18358 43392 24074
rect 43456 19417 43484 24278
rect 43824 23730 43852 26302
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26330 45430 27000
rect 45374 26302 45508 26330
rect 45374 26200 45430 26302
rect 44100 23798 44128 26200
rect 44744 24410 44772 26200
rect 44732 24404 44784 24410
rect 44732 24346 44784 24352
rect 44744 24206 44772 24346
rect 44916 24336 44968 24342
rect 44916 24278 44968 24284
rect 45480 24290 45508 26302
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 44180 24200 44232 24206
rect 44180 24142 44232 24148
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 44088 23792 44140 23798
rect 44088 23734 44140 23740
rect 43812 23724 43864 23730
rect 43812 23666 43864 23672
rect 44192 23322 44220 24142
rect 44640 23724 44692 23730
rect 44640 23666 44692 23672
rect 44364 23520 44416 23526
rect 44364 23462 44416 23468
rect 44180 23316 44232 23322
rect 44180 23258 44232 23264
rect 44376 23118 44404 23462
rect 44652 23322 44680 23666
rect 44928 23594 44956 24278
rect 45480 24262 45600 24290
rect 45572 24206 45600 24262
rect 46032 24206 46060 26200
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 45928 24200 45980 24206
rect 45928 24142 45980 24148
rect 46020 24200 46072 24206
rect 46020 24142 46072 24148
rect 45376 24064 45428 24070
rect 45376 24006 45428 24012
rect 44916 23588 44968 23594
rect 44916 23530 44968 23536
rect 45008 23520 45060 23526
rect 45008 23462 45060 23468
rect 44640 23316 44692 23322
rect 44640 23258 44692 23264
rect 44364 23112 44416 23118
rect 44364 23054 44416 23060
rect 43442 19408 43498 19417
rect 43442 19343 43498 19352
rect 43444 18624 43496 18630
rect 43444 18566 43496 18572
rect 43352 18352 43404 18358
rect 43352 18294 43404 18300
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42800 16992 42852 16998
rect 42800 16934 42852 16940
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 43456 15434 43484 18566
rect 45020 18222 45048 23462
rect 45388 18873 45416 24006
rect 45940 23866 45968 24142
rect 45928 23860 45980 23866
rect 45928 23802 45980 23808
rect 46676 23730 46704 26200
rect 47320 24206 47348 26200
rect 47676 24268 47728 24274
rect 47676 24210 47728 24216
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 47320 23866 47348 24142
rect 47688 23866 47716 24210
rect 47964 24052 47992 26200
rect 48318 24848 48374 24857
rect 48318 24783 48374 24792
rect 47872 24024 47992 24052
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 47676 23860 47728 23866
rect 47676 23802 47728 23808
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 47768 23724 47820 23730
rect 47768 23666 47820 23672
rect 45744 23520 45796 23526
rect 45744 23462 45796 23468
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 45374 18864 45430 18873
rect 45374 18799 45430 18808
rect 45756 18737 45784 23462
rect 46848 22976 46900 22982
rect 46848 22918 46900 22924
rect 46860 22642 46888 22918
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 46204 20800 46256 20806
rect 46204 20742 46256 20748
rect 45742 18728 45798 18737
rect 45742 18663 45798 18672
rect 45008 18216 45060 18222
rect 45008 18158 45060 18164
rect 43444 15428 43496 15434
rect 43444 15370 43496 15376
rect 46216 15366 46244 20742
rect 46952 18970 46980 23462
rect 47492 22976 47544 22982
rect 47492 22918 47544 22924
rect 47504 20806 47532 22918
rect 47780 22778 47808 23666
rect 47872 23118 47900 24024
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 48226 23760 48282 23769
rect 48332 23730 48360 24783
rect 48608 24290 48636 26200
rect 48516 24262 48636 24290
rect 48226 23695 48282 23704
rect 48320 23724 48372 23730
rect 47860 23112 47912 23118
rect 47860 23054 47912 23060
rect 48240 23066 48268 23695
rect 48320 23666 48372 23672
rect 48516 23118 48544 24262
rect 48596 24200 48648 24206
rect 48596 24142 48648 24148
rect 48608 23322 48636 24142
rect 48688 24064 48740 24070
rect 48688 24006 48740 24012
rect 48700 23730 48728 24006
rect 48688 23724 48740 23730
rect 48688 23666 48740 23672
rect 48688 23520 48740 23526
rect 48688 23462 48740 23468
rect 48596 23316 48648 23322
rect 48596 23258 48648 23264
rect 48504 23112 48556 23118
rect 48240 23038 48360 23066
rect 48504 23054 48556 23060
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47768 22772 47820 22778
rect 47768 22714 47820 22720
rect 48332 22642 48360 23038
rect 48412 23044 48464 23050
rect 48412 22986 48464 22992
rect 48320 22636 48372 22642
rect 48320 22578 48372 22584
rect 48424 22166 48452 22986
rect 48504 22432 48556 22438
rect 48504 22374 48556 22380
rect 48412 22160 48464 22166
rect 48412 22102 48464 22108
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47584 21548 47636 21554
rect 47584 21490 47636 21496
rect 47596 21350 47624 21490
rect 47584 21344 47636 21350
rect 47584 21286 47636 21292
rect 47492 20800 47544 20806
rect 47492 20742 47544 20748
rect 46940 18964 46992 18970
rect 46940 18906 46992 18912
rect 46204 15360 46256 15366
rect 46204 15302 46256 15308
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 47596 11150 47624 21286
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 48516 18630 48544 22374
rect 48700 22030 48728 23462
rect 49054 22944 49110 22953
rect 49054 22879 49110 22888
rect 49068 22642 49096 22879
rect 49056 22636 49108 22642
rect 49056 22578 49108 22584
rect 49240 22432 49292 22438
rect 49240 22374 49292 22380
rect 49252 22234 49280 22374
rect 49240 22228 49292 22234
rect 49240 22170 49292 22176
rect 48688 22024 48740 22030
rect 49056 22024 49108 22030
rect 48688 21966 48740 21972
rect 49054 21992 49056 22001
rect 49108 21992 49110 22001
rect 49054 21927 49110 21936
rect 49068 21146 49096 21927
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49056 21140 49108 21146
rect 49056 21082 49108 21088
rect 49160 21049 49188 21422
rect 49146 21040 49202 21049
rect 49146 20975 49202 20984
rect 49252 20058 49280 21830
rect 49240 20052 49292 20058
rect 49240 19994 49292 20000
rect 48504 18624 48556 18630
rect 48504 18566 48556 18572
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47584 11144 47636 11150
rect 47584 11086 47636 11092
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 38752 6180 38804 6186
rect 38752 6122 38804 6128
rect 35716 5636 35768 5642
rect 35716 5578 35768 5584
rect 35728 3534 35756 5578
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37464 4548 37516 4554
rect 37464 4490 37516 4496
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 37476 3058 37504 4490
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 35164 2984 35216 2990
rect 35164 2926 35216 2932
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 31576 2508 31628 2514
rect 31576 2450 31628 2456
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 20088 1142 20208 1170
rect 20088 800 20116 1142
rect 22756 800 22784 2450
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 25412 2304 25464 2310
rect 25412 2246 25464 2252
rect 27804 2304 27856 2310
rect 27804 2246 27856 2252
rect 30748 2304 30800 2310
rect 30748 2246 30800 2252
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 25424 800 25452 2246
rect 1398 0 1454 800
rect 4066 0 4122 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 17406 0 17462 800
rect 20074 0 20130 800
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 27816 762 27844 2246
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28000 870 28120 898
rect 28000 762 28028 870
rect 28092 800 28120 870
rect 30760 800 30788 2246
rect 33428 800 33456 2246
rect 36096 800 36124 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38764 800 38792 6122
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 49424 3460 49476 3466
rect 49424 3402 49476 3408
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 41420 2916 41472 2922
rect 41420 2858 41472 2864
rect 41432 800 41460 2858
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 44100 800 44128 3334
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46768 800 46796 2926
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49436 800 49464 3402
rect 27816 734 28028 762
rect 28078 0 28134 800
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< via2 >>
rect 1582 21392 1638 21448
rect 1306 20712 1362 20768
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2778 24404 2834 24440
rect 2778 24384 2780 24404
rect 2780 24384 2832 24404
rect 2832 24384 2834 24404
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2686 21528 2742 21584
rect 1766 18808 1822 18864
rect 1398 17856 1454 17912
rect 1214 17040 1270 17096
rect 1122 15000 1178 15056
rect 1122 13368 1178 13424
rect 1122 12144 1178 12200
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 1306 15408 1362 15464
rect 1306 14592 1362 14648
rect 2778 21120 2834 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3882 25608 3938 25664
rect 3606 23316 3662 23352
rect 3790 23568 3846 23624
rect 3606 23296 3608 23316
rect 3608 23296 3660 23316
rect 3660 23296 3662 23316
rect 3514 23160 3570 23216
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 1950 19896 2006 19952
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2778 19488 2834 19544
rect 2042 19080 2098 19136
rect 2042 17448 2098 17504
rect 2502 17312 2558 17368
rect 1306 14184 1362 14240
rect 1766 13932 1822 13968
rect 1766 13912 1768 13932
rect 1768 13912 1820 13932
rect 1820 13912 1822 13932
rect 1306 12960 1362 13016
rect 1306 11772 1308 11792
rect 1308 11772 1360 11792
rect 1360 11772 1362 11792
rect 1306 11736 1362 11772
rect 2042 13776 2098 13832
rect 1950 13368 2006 13424
rect 1766 13268 1768 13288
rect 1768 13268 1820 13288
rect 1820 13268 1822 13288
rect 1766 13232 1822 13268
rect 1490 11328 1546 11384
rect 1306 8064 1362 8120
rect 1582 10920 1638 10976
rect 2042 13232 2098 13288
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18672 2926 18728
rect 2778 18264 2834 18320
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2686 17040 2742 17096
rect 2594 10124 2650 10160
rect 2594 10104 2596 10124
rect 2596 10104 2648 10124
rect 2648 10104 2650 10124
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 3698 22752 3754 22808
rect 3790 22344 3846 22400
rect 3606 19216 3662 19272
rect 3606 18672 3662 18728
rect 3790 21528 3846 21584
rect 4066 25200 4122 25256
rect 4066 24812 4122 24848
rect 4066 24792 4068 24812
rect 4068 24792 4120 24812
rect 4120 24792 4122 24812
rect 4066 23976 4122 24032
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 4066 23180 4122 23216
rect 4066 23160 4068 23180
rect 4068 23160 4120 23180
rect 4120 23160 4122 23180
rect 4158 22616 4214 22672
rect 4066 22480 4122 22536
rect 4066 21936 4122 21992
rect 4250 21004 4306 21040
rect 4250 20984 4252 21004
rect 4252 20984 4304 21004
rect 4304 20984 4306 21004
rect 3882 19660 3884 19680
rect 3884 19660 3936 19680
rect 3936 19660 3938 19680
rect 3882 19624 3938 19660
rect 3790 19080 3846 19136
rect 3790 17856 3846 17912
rect 3422 17176 3478 17232
rect 3606 16788 3662 16824
rect 3606 16768 3608 16788
rect 3608 16768 3660 16788
rect 3660 16768 3662 16788
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 3238 10648 3294 10704
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2870 9696 2926 9752
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2778 7248 2834 7304
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3514 13776 3570 13832
rect 3698 13504 3754 13560
rect 3882 16088 3938 16144
rect 3974 15952 4030 16008
rect 3422 11872 3478 11928
rect 3422 9016 3478 9072
rect 1214 6432 1270 6488
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3790 10648 3846 10704
rect 3606 9968 3662 10024
rect 3698 9424 3754 9480
rect 3882 10512 3938 10568
rect 3698 8356 3754 8392
rect 3698 8336 3700 8356
rect 3700 8336 3752 8356
rect 3752 8336 3754 8356
rect 3698 7656 3754 7712
rect 3606 7384 3662 7440
rect 1306 6024 1362 6080
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 4250 19896 4306 19952
rect 4342 19080 4398 19136
rect 4250 18264 4306 18320
rect 4434 16904 4490 16960
rect 4250 13132 4252 13152
rect 4252 13132 4304 13152
rect 4304 13132 4306 13152
rect 4250 13096 4306 13132
rect 4434 13640 4490 13696
rect 4710 18944 4766 19000
rect 6550 23432 6606 23488
rect 4894 17720 4950 17776
rect 4618 13504 4674 13560
rect 4250 12688 4306 12744
rect 4158 11212 4214 11248
rect 4158 11192 4160 11212
rect 4160 11192 4212 11212
rect 4212 11192 4214 11212
rect 3974 9288 4030 9344
rect 4158 8880 4214 8936
rect 3974 7268 4030 7304
rect 3974 7248 3976 7268
rect 3976 7248 4028 7268
rect 4028 7248 4030 7268
rect 4250 8472 4306 8528
rect 4066 6840 4122 6896
rect 5538 21428 5540 21448
rect 5540 21428 5592 21448
rect 5592 21428 5594 21448
rect 5538 21392 5594 21428
rect 5078 16532 5080 16552
rect 5080 16532 5132 16552
rect 5132 16532 5134 16552
rect 5078 16496 5134 16532
rect 5354 18164 5356 18184
rect 5356 18164 5408 18184
rect 5408 18164 5410 18184
rect 5354 18128 5410 18164
rect 5630 21256 5686 21312
rect 5630 20168 5686 20224
rect 5722 19372 5778 19408
rect 5722 19352 5724 19372
rect 5724 19352 5776 19372
rect 5776 19352 5778 19372
rect 5630 17992 5686 18048
rect 5446 15136 5502 15192
rect 5354 14456 5410 14512
rect 4894 12280 4950 12336
rect 5078 11872 5134 11928
rect 5906 17720 5962 17776
rect 5906 16652 5962 16688
rect 6826 23024 6882 23080
rect 6458 20848 6514 20904
rect 6458 19352 6514 19408
rect 5906 16632 5908 16652
rect 5908 16632 5960 16652
rect 5960 16632 5962 16652
rect 5722 15000 5778 15056
rect 5906 14864 5962 14920
rect 5078 11328 5134 11384
rect 4526 8744 4582 8800
rect 5170 11056 5226 11112
rect 5446 9560 5502 9616
rect 5906 9832 5962 9888
rect 5814 9696 5870 9752
rect 5354 7404 5410 7440
rect 5354 7384 5356 7404
rect 5356 7384 5408 7404
rect 5408 7384 5410 7404
rect 1306 5228 1362 5264
rect 1306 5208 1308 5228
rect 1308 5208 1360 5228
rect 1360 5208 1362 5228
rect 1306 4800 1362 4856
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 1306 3168 1362 3224
rect 1306 2760 1362 2816
rect 1214 2352 1270 2408
rect 1306 1944 1362 2000
rect 4158 4392 4214 4448
rect 4066 3984 4122 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2870 3576 2926 3632
rect 5722 7964 5724 7984
rect 5724 7964 5776 7984
rect 5776 7964 5778 7984
rect 5722 7928 5778 7964
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2870 1536 2926 1592
rect 6458 17060 6514 17096
rect 6458 17040 6460 17060
rect 6460 17040 6512 17060
rect 6512 17040 6514 17060
rect 6642 20168 6698 20224
rect 6918 20712 6974 20768
rect 6642 15000 6698 15056
rect 6366 13812 6368 13832
rect 6368 13812 6420 13832
rect 6420 13812 6422 13832
rect 6366 13776 6422 13812
rect 6182 10784 6238 10840
rect 7194 22616 7250 22672
rect 7102 21392 7158 21448
rect 7102 17584 7158 17640
rect 7286 17720 7342 17776
rect 7470 22616 7526 22672
rect 7562 21256 7618 21312
rect 7562 20032 7618 20088
rect 7470 18672 7526 18728
rect 7562 18148 7618 18184
rect 7562 18128 7564 18148
rect 7564 18128 7616 18148
rect 7616 18128 7618 18148
rect 7102 15136 7158 15192
rect 6550 12416 6606 12472
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7930 21120 7986 21176
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 8390 22072 8446 22128
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 9862 24248 9918 24304
rect 8574 18672 8630 18728
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7746 17312 7802 17368
rect 7378 14864 7434 14920
rect 7194 12824 7250 12880
rect 7286 12688 7342 12744
rect 7194 9172 7250 9208
rect 7194 9152 7196 9172
rect 7196 9152 7248 9172
rect 7248 9152 7250 9172
rect 7378 11192 7434 11248
rect 6366 8084 6422 8120
rect 6366 8064 6368 8084
rect 6368 8064 6420 8084
rect 6420 8064 6422 8084
rect 6550 8200 6606 8256
rect 7562 9152 7618 9208
rect 8206 17040 8262 17096
rect 8114 16652 8170 16688
rect 8114 16632 8116 16652
rect 8116 16632 8168 16652
rect 8168 16632 8170 16652
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7930 15952 7986 16008
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7930 14900 7932 14920
rect 7932 14900 7984 14920
rect 7984 14900 7986 14920
rect 7930 14864 7986 14900
rect 7746 12144 7802 12200
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 8390 17196 8446 17232
rect 8390 17176 8392 17196
rect 8392 17176 8444 17196
rect 8444 17176 8446 17196
rect 8574 17332 8630 17368
rect 8574 17312 8576 17332
rect 8576 17312 8628 17332
rect 8628 17312 8630 17332
rect 8574 16768 8630 16824
rect 8482 15272 8538 15328
rect 8390 15136 8446 15192
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 8574 14456 8630 14512
rect 8574 11056 8630 11112
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7930 8492 7986 8528
rect 7930 8472 7932 8492
rect 7932 8472 7984 8492
rect 7984 8472 7986 8492
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 8758 21972 8760 21992
rect 8760 21972 8812 21992
rect 8812 21972 8814 21992
rect 8758 21936 8814 21972
rect 8850 16244 8906 16280
rect 8850 16224 8852 16244
rect 8852 16224 8904 16244
rect 8904 16224 8906 16244
rect 8850 11328 8906 11384
rect 9126 17992 9182 18048
rect 9770 22480 9826 22536
rect 9586 20576 9642 20632
rect 9402 18944 9458 19000
rect 9494 17992 9550 18048
rect 9770 19488 9826 19544
rect 10506 21528 10562 21584
rect 9954 19216 10010 19272
rect 9862 17040 9918 17096
rect 9770 16396 9772 16416
rect 9772 16396 9824 16416
rect 9824 16396 9826 16416
rect 9770 16360 9826 16396
rect 9770 16088 9826 16144
rect 9678 15680 9734 15736
rect 9586 15408 9642 15464
rect 9034 11600 9090 11656
rect 9402 13388 9458 13424
rect 9402 13368 9404 13388
rect 9404 13368 9456 13388
rect 9456 13368 9458 13388
rect 10414 17856 10470 17912
rect 9954 15408 10010 15464
rect 9586 12824 9642 12880
rect 10414 16768 10470 16824
rect 11150 24656 11206 24712
rect 10506 16396 10508 16416
rect 10508 16396 10560 16416
rect 10560 16396 10562 16416
rect 10506 16360 10562 16396
rect 11794 23160 11850 23216
rect 11794 22888 11850 22944
rect 11886 22752 11942 22808
rect 12530 23432 12586 23488
rect 12254 22072 12310 22128
rect 11150 21392 11206 21448
rect 11334 20712 11390 20768
rect 11426 19896 11482 19952
rect 11334 18808 11390 18864
rect 11426 18164 11428 18184
rect 11428 18164 11480 18184
rect 11480 18164 11482 18184
rect 11426 18128 11482 18164
rect 11058 17176 11114 17232
rect 10874 16768 10930 16824
rect 10782 16632 10838 16688
rect 11150 16496 11206 16552
rect 10690 16224 10746 16280
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 9862 8356 9918 8392
rect 9862 8336 9864 8356
rect 9864 8336 9916 8356
rect 9916 8336 9918 8356
rect 10506 14764 10508 14784
rect 10508 14764 10560 14784
rect 10560 14764 10562 14784
rect 10506 14728 10562 14764
rect 10690 12844 10746 12880
rect 10690 12824 10692 12844
rect 10692 12824 10744 12844
rect 10744 12824 10746 12844
rect 10966 15972 11022 16008
rect 10966 15952 10968 15972
rect 10968 15952 11020 15972
rect 11020 15952 11022 15972
rect 11426 15272 11482 15328
rect 11426 15136 11482 15192
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 11058 9988 11114 10024
rect 11058 9968 11060 9988
rect 11060 9968 11112 9988
rect 11112 9968 11114 9988
rect 12162 21392 12218 21448
rect 11794 20848 11850 20904
rect 11794 19760 11850 19816
rect 11886 19352 11942 19408
rect 11886 18672 11942 18728
rect 11610 16496 11666 16552
rect 11610 16244 11666 16280
rect 11610 16224 11612 16244
rect 11612 16224 11664 16244
rect 11664 16224 11666 16244
rect 11518 11056 11574 11112
rect 12530 22072 12586 22128
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 13266 23568 13322 23624
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 14646 24792 14702 24848
rect 14278 24112 14334 24168
rect 12162 17448 12218 17504
rect 12254 15680 12310 15736
rect 12070 15580 12072 15600
rect 12072 15580 12124 15600
rect 12124 15580 12126 15600
rect 12070 15544 12126 15580
rect 11978 15020 12034 15056
rect 11978 15000 11980 15020
rect 11980 15000 12032 15020
rect 12032 15000 12034 15020
rect 12346 14320 12402 14376
rect 11886 13096 11942 13152
rect 11610 9968 11666 10024
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 13910 21256 13966 21312
rect 13910 20748 13912 20768
rect 13912 20748 13964 20768
rect 13964 20748 13966 20768
rect 13910 20712 13966 20748
rect 13358 20304 13414 20360
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13450 18944 13506 19000
rect 13726 19488 13782 19544
rect 13358 18264 13414 18320
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13726 19080 13782 19136
rect 13726 18536 13782 18592
rect 12806 17448 12862 17504
rect 12990 17448 13046 17504
rect 12622 16788 12678 16824
rect 12622 16768 12624 16788
rect 12624 16768 12676 16788
rect 12676 16768 12678 16788
rect 12622 15272 12678 15328
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12898 14320 12954 14376
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13818 16496 13874 16552
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12438 8472 12494 8528
rect 13726 15680 13782 15736
rect 13818 15136 13874 15192
rect 14554 22888 14610 22944
rect 14370 22344 14426 22400
rect 14554 21972 14556 21992
rect 14556 21972 14608 21992
rect 14608 21972 14610 21992
rect 14554 21936 14610 21972
rect 14278 20168 14334 20224
rect 14186 18264 14242 18320
rect 14002 18128 14058 18184
rect 14462 18844 14464 18864
rect 14464 18844 14516 18864
rect 14516 18844 14518 18864
rect 14462 18808 14518 18844
rect 14462 17584 14518 17640
rect 14370 16496 14426 16552
rect 14370 14728 14426 14784
rect 14370 14612 14426 14648
rect 14370 14592 14372 14612
rect 14372 14592 14424 14612
rect 14424 14592 14426 14612
rect 15474 25200 15530 25256
rect 14830 17856 14886 17912
rect 15658 25064 15714 25120
rect 15566 21412 15622 21448
rect 15566 21392 15568 21412
rect 15568 21392 15620 21412
rect 15620 21392 15622 21412
rect 16026 23432 16082 23488
rect 15750 20748 15752 20768
rect 15752 20748 15804 20768
rect 15804 20748 15806 20768
rect 15750 20712 15806 20748
rect 16486 23704 16542 23760
rect 15934 21548 15990 21584
rect 15934 21528 15936 21548
rect 15936 21528 15988 21548
rect 15988 21528 15990 21548
rect 16578 21140 16634 21176
rect 16578 21120 16580 21140
rect 16580 21120 16632 21140
rect 16632 21120 16634 21140
rect 16118 20596 16174 20632
rect 16118 20576 16120 20596
rect 16120 20576 16172 20596
rect 16172 20576 16174 20596
rect 15198 18808 15254 18864
rect 15382 18808 15438 18864
rect 15106 18400 15162 18456
rect 15014 18148 15070 18184
rect 15014 18128 15016 18148
rect 15016 18128 15068 18148
rect 15068 18128 15070 18148
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12806 9152 12862 9208
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 16486 18284 16542 18320
rect 16486 18264 16488 18284
rect 16488 18264 16540 18284
rect 16540 18264 16542 18284
rect 16486 17720 16542 17776
rect 16210 17584 16266 17640
rect 16210 16396 16212 16416
rect 16212 16396 16264 16416
rect 16264 16396 16266 16416
rect 16210 16360 16266 16396
rect 16486 16768 16542 16824
rect 15750 12144 15806 12200
rect 17590 23160 17646 23216
rect 17590 22888 17646 22944
rect 17498 22616 17554 22672
rect 17222 19932 17224 19952
rect 17224 19932 17276 19952
rect 17276 19932 17278 19952
rect 17222 19896 17278 19932
rect 16946 16124 16948 16144
rect 16948 16124 17000 16144
rect 17000 16124 17002 16144
rect 16946 16088 17002 16124
rect 17130 16244 17186 16280
rect 17130 16224 17132 16244
rect 17132 16224 17184 16244
rect 17184 16224 17186 16244
rect 17130 14864 17186 14920
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17774 22752 17830 22808
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17866 20868 17922 20904
rect 17866 20848 17868 20868
rect 17868 20848 17920 20868
rect 17920 20848 17922 20868
rect 17774 20712 17830 20768
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17958 20168 18014 20224
rect 19154 24384 19210 24440
rect 19522 22752 19578 22808
rect 18602 21256 18658 21312
rect 18602 20032 18658 20088
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18602 19624 18658 19680
rect 18694 19080 18750 19136
rect 18602 18944 18658 19000
rect 18786 17312 18842 17368
rect 18786 16768 18842 16824
rect 18510 15136 18566 15192
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18510 14728 18566 14784
rect 17406 12044 17408 12064
rect 17408 12044 17460 12064
rect 17460 12044 17462 12064
rect 17406 12008 17462 12044
rect 16578 8472 16634 8528
rect 17682 12280 17738 12336
rect 18418 12280 18474 12336
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18694 13232 18750 13288
rect 18970 17176 19026 17232
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18786 10648 18842 10704
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 19154 14320 19210 14376
rect 19338 19488 19394 19544
rect 19338 16360 19394 16416
rect 19706 17584 19762 17640
rect 19338 14864 19394 14920
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 21362 23704 21418 23760
rect 19982 20440 20038 20496
rect 19982 18400 20038 18456
rect 20074 17856 20130 17912
rect 20626 22480 20682 22536
rect 20626 21800 20682 21856
rect 20074 15272 20130 15328
rect 19982 14864 20038 14920
rect 19890 13912 19946 13968
rect 20626 17176 20682 17232
rect 21086 17196 21142 17232
rect 21086 17176 21088 17196
rect 21088 17176 21140 17196
rect 21140 17176 21142 17196
rect 21270 16632 21326 16688
rect 21270 16088 21326 16144
rect 22558 23568 22614 23624
rect 22190 22888 22246 22944
rect 22466 22480 22522 22536
rect 21454 17332 21510 17368
rect 21454 17312 21456 17332
rect 21456 17312 21508 17332
rect 21508 17312 21510 17332
rect 21638 17212 21640 17232
rect 21640 17212 21692 17232
rect 21692 17212 21694 17232
rect 21638 17176 21694 17212
rect 21546 15680 21602 15736
rect 22374 20712 22430 20768
rect 22282 14864 22338 14920
rect 22466 18844 22468 18864
rect 22468 18844 22520 18864
rect 22520 18844 22522 18864
rect 22466 18808 22522 18844
rect 22374 14320 22430 14376
rect 22098 12824 22154 12880
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22834 23568 22890 23624
rect 22742 23296 22798 23352
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23110 23160 23166 23216
rect 23294 23160 23350 23216
rect 23110 22888 23166 22944
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22742 21120 22798 21176
rect 22742 18944 22798 19000
rect 22742 18536 22798 18592
rect 23294 21836 23296 21856
rect 23296 21836 23348 21856
rect 23348 21836 23350 21856
rect 23294 21800 23350 21836
rect 23570 21800 23626 21856
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23478 21256 23534 21312
rect 23294 20576 23350 20632
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22742 14320 22798 14376
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 24214 20848 24270 20904
rect 24030 18400 24086 18456
rect 24030 17584 24086 17640
rect 23846 16632 23902 16688
rect 24490 22888 24546 22944
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23386 14320 23442 14376
rect 23662 14884 23718 14920
rect 23662 14864 23664 14884
rect 23664 14864 23716 14884
rect 23716 14864 23718 14884
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 24766 23432 24822 23488
rect 25318 22480 25374 22536
rect 24950 21800 25006 21856
rect 24766 18536 24822 18592
rect 24766 16088 24822 16144
rect 25134 18944 25190 19000
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 26146 24112 26202 24168
rect 27710 25200 27766 25256
rect 26330 23704 26386 23760
rect 25778 22344 25834 22400
rect 26606 23468 26608 23488
rect 26608 23468 26660 23488
rect 26660 23468 26662 23488
rect 26606 23432 26662 23468
rect 25962 20032 26018 20088
rect 25962 19488 26018 19544
rect 25870 18808 25926 18864
rect 25410 17856 25466 17912
rect 27158 22752 27214 22808
rect 26974 22480 27030 22536
rect 27250 22344 27306 22400
rect 27158 22208 27214 22264
rect 27066 21664 27122 21720
rect 27250 21256 27306 21312
rect 27066 20984 27122 21040
rect 27066 20596 27122 20632
rect 27066 20576 27068 20596
rect 27068 20576 27120 20596
rect 27120 20576 27122 20596
rect 27434 23296 27490 23352
rect 27526 22072 27582 22128
rect 27526 21256 27582 21312
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 28630 23568 28686 23624
rect 28538 22752 28594 22808
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27158 20168 27214 20224
rect 27618 19624 27674 19680
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 28630 21800 28686 21856
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 26974 19252 26976 19272
rect 26976 19252 27028 19272
rect 27028 19252 27030 19272
rect 26974 19216 27030 19252
rect 26146 16360 26202 16416
rect 27618 18128 27674 18184
rect 27434 17876 27490 17912
rect 27434 17856 27436 17876
rect 27436 17856 27488 17876
rect 27488 17856 27490 17876
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 29550 21800 29606 21856
rect 28722 20168 28778 20224
rect 29826 21392 29882 21448
rect 28998 19896 29054 19952
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 25594 15136 25650 15192
rect 30102 20304 30158 20360
rect 29826 19624 29882 19680
rect 28354 16496 28410 16552
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 31022 22480 31078 22536
rect 32034 22752 32090 22808
rect 31942 22072 31998 22128
rect 32126 22208 32182 22264
rect 30838 20032 30894 20088
rect 30746 19660 30748 19680
rect 30748 19660 30800 19680
rect 30800 19660 30802 19680
rect 30746 19624 30802 19660
rect 30654 19372 30710 19408
rect 30654 19352 30656 19372
rect 30656 19352 30708 19372
rect 30708 19352 30710 19372
rect 30838 19352 30894 19408
rect 30194 17584 30250 17640
rect 31206 17040 31262 17096
rect 30102 15952 30158 16008
rect 29918 15544 29974 15600
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 32402 22072 32458 22128
rect 31390 13368 31446 13424
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27710 10104 27766 10160
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 32126 20712 32182 20768
rect 32034 15408 32090 15464
rect 32310 20032 32366 20088
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32678 21392 32734 21448
rect 32770 21292 32772 21312
rect 32772 21292 32824 21312
rect 32824 21292 32826 21312
rect 32770 21256 32826 21292
rect 32678 21120 32734 21176
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 33414 21392 33470 21448
rect 32862 20712 32918 20768
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 33690 24656 33746 24712
rect 33874 25064 33930 25120
rect 34058 24792 34114 24848
rect 34242 23160 34298 23216
rect 36174 24928 36230 24984
rect 35622 23044 35678 23080
rect 35622 23024 35624 23044
rect 35624 23024 35676 23044
rect 35676 23024 35678 23044
rect 34518 22636 34574 22672
rect 34518 22616 34520 22636
rect 34520 22616 34572 22636
rect 34572 22616 34574 22636
rect 34518 20984 34574 21040
rect 33506 17720 33562 17776
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 35070 21936 35126 21992
rect 34058 15000 34114 15056
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 36266 21528 36322 21584
rect 36450 20440 36506 20496
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 38658 24248 38714 24304
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 40682 20848 40738 20904
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 43442 19352 43498 19408
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 48318 24792 48374 24848
rect 45374 18808 45430 18864
rect 45742 18672 45798 18728
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 48226 23704 48282 23760
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 49054 22888 49110 22944
rect 49054 21972 49056 21992
rect 49056 21972 49108 21992
rect 49108 21972 49110 21992
rect 49054 21936 49110 21972
rect 49146 20984 49202 21040
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3877 25666 3943 25669
rect 0 25664 3943 25666
rect 0 25608 3882 25664
rect 3938 25608 3943 25664
rect 0 25606 3943 25608
rect 0 25576 800 25606
rect 3877 25603 3943 25606
rect 0 25258 800 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 800 25198
rect 4061 25195 4127 25198
rect 15469 25258 15535 25261
rect 27705 25258 27771 25261
rect 15469 25256 27771 25258
rect 15469 25200 15474 25256
rect 15530 25200 27710 25256
rect 27766 25200 27771 25256
rect 15469 25198 27771 25200
rect 15469 25195 15535 25198
rect 27705 25195 27771 25198
rect 15653 25122 15719 25125
rect 33869 25122 33935 25125
rect 15653 25120 33935 25122
rect 15653 25064 15658 25120
rect 15714 25064 33874 25120
rect 33930 25064 33935 25120
rect 15653 25062 33935 25064
rect 15653 25059 15719 25062
rect 33869 25059 33935 25062
rect 11646 24924 11652 24988
rect 11716 24986 11722 24988
rect 36169 24986 36235 24989
rect 11716 24984 36235 24986
rect 11716 24928 36174 24984
rect 36230 24928 36235 24984
rect 11716 24926 36235 24928
rect 11716 24924 11722 24926
rect 36169 24923 36235 24926
rect 0 24850 800 24880
rect 4061 24850 4127 24853
rect 0 24848 4127 24850
rect 0 24792 4066 24848
rect 4122 24792 4127 24848
rect 0 24790 4127 24792
rect 0 24760 800 24790
rect 4061 24787 4127 24790
rect 14641 24850 14707 24853
rect 34053 24850 34119 24853
rect 14641 24848 34119 24850
rect 14641 24792 14646 24848
rect 14702 24792 34058 24848
rect 34114 24792 34119 24848
rect 14641 24790 34119 24792
rect 14641 24787 14707 24790
rect 34053 24787 34119 24790
rect 48313 24850 48379 24853
rect 50200 24850 51000 24880
rect 48313 24848 51000 24850
rect 48313 24792 48318 24848
rect 48374 24792 51000 24848
rect 48313 24790 51000 24792
rect 48313 24787 48379 24790
rect 50200 24760 51000 24790
rect 11145 24714 11211 24717
rect 33685 24714 33751 24717
rect 11145 24712 33751 24714
rect 11145 24656 11150 24712
rect 11206 24656 33690 24712
rect 33746 24656 33751 24712
rect 11145 24654 33751 24656
rect 11145 24651 11211 24654
rect 33685 24651 33751 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 19149 24442 19215 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 18278 24440 19215 24442
rect 18278 24384 19154 24440
rect 19210 24384 19215 24440
rect 18278 24382 19215 24384
rect 9857 24306 9923 24309
rect 18278 24306 18338 24382
rect 19149 24379 19215 24382
rect 9857 24304 18338 24306
rect 9857 24248 9862 24304
rect 9918 24248 18338 24304
rect 9857 24246 18338 24248
rect 9857 24243 9923 24246
rect 18454 24244 18460 24308
rect 18524 24306 18530 24308
rect 38653 24306 38719 24309
rect 18524 24304 38719 24306
rect 18524 24248 38658 24304
rect 38714 24248 38719 24304
rect 18524 24246 38719 24248
rect 18524 24244 18530 24246
rect 38653 24243 38719 24246
rect 14273 24170 14339 24173
rect 26141 24170 26207 24173
rect 14273 24168 26207 24170
rect 14273 24112 14278 24168
rect 14334 24112 26146 24168
rect 26202 24112 26207 24168
rect 14273 24110 26207 24112
rect 14273 24107 14339 24110
rect 26141 24107 26207 24110
rect 0 24034 800 24064
rect 4061 24034 4127 24037
rect 0 24032 4127 24034
rect 0 23976 4066 24032
rect 4122 23976 4127 24032
rect 0 23974 4127 23976
rect 0 23944 800 23974
rect 4061 23971 4127 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 50200 23898 51000 23928
rect 48454 23838 51000 23898
rect 16481 23762 16547 23765
rect 21357 23762 21423 23765
rect 26325 23762 26391 23765
rect 16481 23760 21423 23762
rect 16481 23704 16486 23760
rect 16542 23704 21362 23760
rect 21418 23704 21423 23760
rect 16481 23702 21423 23704
rect 16481 23699 16547 23702
rect 21357 23699 21423 23702
rect 22694 23760 26391 23762
rect 22694 23704 26330 23760
rect 26386 23704 26391 23760
rect 22694 23702 26391 23704
rect 0 23626 800 23656
rect 3785 23626 3851 23629
rect 0 23624 3851 23626
rect 0 23568 3790 23624
rect 3846 23568 3851 23624
rect 0 23566 3851 23568
rect 0 23536 800 23566
rect 3785 23563 3851 23566
rect 13261 23626 13327 23629
rect 22553 23626 22619 23629
rect 13261 23624 22619 23626
rect 13261 23568 13266 23624
rect 13322 23568 22558 23624
rect 22614 23568 22619 23624
rect 13261 23566 22619 23568
rect 13261 23563 13327 23566
rect 22553 23563 22619 23566
rect 6545 23492 6611 23493
rect 6494 23428 6500 23492
rect 6564 23490 6611 23492
rect 12525 23490 12591 23493
rect 6564 23488 6656 23490
rect 6606 23432 6656 23488
rect 6564 23430 6656 23432
rect 12390 23488 12591 23490
rect 12390 23432 12530 23488
rect 12586 23432 12591 23488
rect 12390 23430 12591 23432
rect 6564 23428 6611 23430
rect 6545 23427 6611 23428
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 3601 23354 3667 23357
rect 12390 23354 12450 23430
rect 12525 23427 12591 23430
rect 16021 23490 16087 23493
rect 22694 23490 22754 23702
rect 26325 23699 26391 23702
rect 48221 23762 48287 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 48221 23760 48514 23762
rect 48221 23704 48226 23760
rect 48282 23704 48514 23760
rect 48221 23702 48514 23704
rect 48221 23699 48287 23702
rect 22829 23626 22895 23629
rect 28625 23626 28691 23629
rect 22829 23624 28691 23626
rect 22829 23568 22834 23624
rect 22890 23568 28630 23624
rect 28686 23568 28691 23624
rect 22829 23566 28691 23568
rect 22829 23563 22895 23566
rect 28625 23563 28691 23566
rect 16021 23488 22754 23490
rect 16021 23432 16026 23488
rect 16082 23432 22754 23488
rect 16021 23430 22754 23432
rect 24761 23490 24827 23493
rect 26601 23490 26667 23493
rect 24761 23488 26986 23490
rect 24761 23432 24766 23488
rect 24822 23432 26606 23488
rect 26662 23432 26986 23488
rect 24761 23430 26986 23432
rect 16021 23427 16087 23430
rect 24761 23427 24827 23430
rect 26601 23427 26667 23430
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 22737 23354 22803 23357
rect 3601 23352 12450 23354
rect 3601 23296 3606 23352
rect 3662 23296 12450 23352
rect 3601 23294 12450 23296
rect 17174 23352 22803 23354
rect 17174 23296 22742 23352
rect 22798 23296 22803 23352
rect 17174 23294 22803 23296
rect 26926 23354 26986 23430
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 27429 23354 27495 23357
rect 26926 23352 27495 23354
rect 26926 23296 27434 23352
rect 27490 23296 27495 23352
rect 26926 23294 27495 23296
rect 3601 23291 3667 23294
rect 0 23218 800 23248
rect 3509 23218 3575 23221
rect 0 23216 3575 23218
rect 0 23160 3514 23216
rect 3570 23160 3575 23216
rect 0 23158 3575 23160
rect 0 23128 800 23158
rect 3509 23155 3575 23158
rect 4061 23218 4127 23221
rect 11789 23218 11855 23221
rect 17174 23218 17234 23294
rect 22737 23291 22803 23294
rect 27429 23291 27495 23294
rect 4061 23216 11855 23218
rect 4061 23160 4066 23216
rect 4122 23160 11794 23216
rect 11850 23160 11855 23216
rect 4061 23158 11855 23160
rect 4061 23155 4127 23158
rect 11789 23155 11855 23158
rect 12206 23158 17234 23218
rect 17585 23218 17651 23221
rect 23105 23218 23171 23221
rect 17585 23216 23171 23218
rect 17585 23160 17590 23216
rect 17646 23160 23110 23216
rect 23166 23160 23171 23216
rect 17585 23158 23171 23160
rect 6310 23020 6316 23084
rect 6380 23082 6386 23084
rect 6821 23082 6887 23085
rect 12206 23082 12266 23158
rect 17585 23155 17651 23158
rect 23105 23155 23171 23158
rect 23289 23218 23355 23221
rect 34237 23218 34303 23221
rect 23289 23216 34303 23218
rect 23289 23160 23294 23216
rect 23350 23160 34242 23216
rect 34298 23160 34303 23216
rect 23289 23158 34303 23160
rect 23289 23155 23355 23158
rect 34237 23155 34303 23158
rect 35617 23082 35683 23085
rect 6380 23080 12266 23082
rect 6380 23024 6826 23080
rect 6882 23024 12266 23080
rect 6380 23022 12266 23024
rect 12390 23080 35683 23082
rect 12390 23024 35622 23080
rect 35678 23024 35683 23080
rect 12390 23022 35683 23024
rect 6380 23020 6386 23022
rect 6821 23019 6887 23022
rect 11789 22946 11855 22949
rect 12390 22946 12450 23022
rect 35617 23019 35683 23022
rect 11789 22944 12450 22946
rect 11789 22888 11794 22944
rect 11850 22888 12450 22944
rect 11789 22886 12450 22888
rect 14549 22946 14615 22949
rect 17585 22946 17651 22949
rect 22185 22948 22251 22949
rect 22134 22946 22140 22948
rect 14549 22944 17651 22946
rect 14549 22888 14554 22944
rect 14610 22888 17590 22944
rect 17646 22888 17651 22944
rect 14549 22886 17651 22888
rect 22094 22886 22140 22946
rect 22204 22944 22251 22948
rect 22246 22888 22251 22944
rect 11789 22883 11855 22886
rect 14549 22883 14615 22886
rect 17585 22883 17651 22886
rect 22134 22884 22140 22886
rect 22204 22884 22251 22888
rect 22185 22883 22251 22884
rect 23105 22946 23171 22949
rect 24485 22946 24551 22949
rect 23105 22944 24551 22946
rect 23105 22888 23110 22944
rect 23166 22888 24490 22944
rect 24546 22888 24551 22944
rect 23105 22886 24551 22888
rect 23105 22883 23171 22886
rect 24485 22883 24551 22886
rect 49049 22946 49115 22949
rect 50200 22946 51000 22976
rect 49049 22944 51000 22946
rect 49049 22888 49054 22944
rect 49110 22888 51000 22944
rect 49049 22886 51000 22888
rect 49049 22883 49115 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 50200 22856 51000 22886
rect 47946 22815 48262 22816
rect 3693 22810 3759 22813
rect 0 22808 3759 22810
rect 0 22752 3698 22808
rect 3754 22752 3759 22808
rect 0 22750 3759 22752
rect 0 22720 800 22750
rect 3693 22747 3759 22750
rect 10174 22748 10180 22812
rect 10244 22810 10250 22812
rect 11881 22810 11947 22813
rect 17769 22810 17835 22813
rect 10244 22808 11947 22810
rect 10244 22752 11886 22808
rect 11942 22752 11947 22808
rect 10244 22750 11947 22752
rect 10244 22748 10250 22750
rect 11881 22747 11947 22750
rect 12390 22808 17835 22810
rect 12390 22752 17774 22808
rect 17830 22752 17835 22808
rect 12390 22750 17835 22752
rect 4153 22674 4219 22677
rect 7189 22676 7255 22677
rect 5390 22674 5396 22676
rect 4153 22672 5396 22674
rect 4153 22616 4158 22672
rect 4214 22616 5396 22672
rect 4153 22614 5396 22616
rect 4153 22611 4219 22614
rect 5390 22612 5396 22614
rect 5460 22612 5466 22676
rect 7189 22672 7236 22676
rect 7300 22674 7306 22676
rect 7465 22674 7531 22677
rect 12390 22674 12450 22750
rect 17769 22747 17835 22750
rect 19517 22810 19583 22813
rect 27153 22810 27219 22813
rect 19517 22808 27219 22810
rect 19517 22752 19522 22808
rect 19578 22752 27158 22808
rect 27214 22752 27219 22808
rect 19517 22750 27219 22752
rect 19517 22747 19583 22750
rect 27153 22747 27219 22750
rect 28533 22810 28599 22813
rect 32029 22810 32095 22813
rect 28533 22808 32095 22810
rect 28533 22752 28538 22808
rect 28594 22752 32034 22808
rect 32090 22752 32095 22808
rect 28533 22750 32095 22752
rect 28533 22747 28599 22750
rect 32029 22747 32095 22750
rect 7189 22616 7194 22672
rect 7189 22612 7236 22616
rect 7300 22614 7346 22674
rect 7465 22672 12450 22674
rect 7465 22616 7470 22672
rect 7526 22616 12450 22672
rect 7465 22614 12450 22616
rect 17493 22674 17559 22677
rect 34513 22674 34579 22677
rect 17493 22672 34579 22674
rect 17493 22616 17498 22672
rect 17554 22616 34518 22672
rect 34574 22616 34579 22672
rect 17493 22614 34579 22616
rect 7300 22612 7306 22614
rect 7189 22611 7255 22612
rect 7465 22611 7531 22614
rect 17493 22611 17559 22614
rect 34513 22611 34579 22614
rect 4061 22538 4127 22541
rect 2270 22536 4127 22538
rect 2270 22480 4066 22536
rect 4122 22480 4127 22536
rect 2270 22478 4127 22480
rect 0 22402 800 22432
rect 2270 22402 2330 22478
rect 4061 22475 4127 22478
rect 9765 22538 9831 22541
rect 20621 22538 20687 22541
rect 9765 22536 20687 22538
rect 9765 22480 9770 22536
rect 9826 22480 20626 22536
rect 20682 22480 20687 22536
rect 9765 22478 20687 22480
rect 9765 22475 9831 22478
rect 20621 22475 20687 22478
rect 22461 22538 22527 22541
rect 25313 22538 25379 22541
rect 22461 22536 25379 22538
rect 22461 22480 22466 22536
rect 22522 22480 25318 22536
rect 25374 22480 25379 22536
rect 22461 22478 25379 22480
rect 22461 22475 22527 22478
rect 25313 22475 25379 22478
rect 26969 22538 27035 22541
rect 31017 22538 31083 22541
rect 26969 22536 31083 22538
rect 26969 22480 26974 22536
rect 27030 22480 31022 22536
rect 31078 22480 31083 22536
rect 26969 22478 31083 22480
rect 26969 22475 27035 22478
rect 31017 22475 31083 22478
rect 0 22342 2330 22402
rect 3785 22402 3851 22405
rect 3918 22402 3924 22404
rect 3785 22400 3924 22402
rect 3785 22344 3790 22400
rect 3846 22344 3924 22400
rect 3785 22342 3924 22344
rect 0 22312 800 22342
rect 3785 22339 3851 22342
rect 3918 22340 3924 22342
rect 3988 22340 3994 22404
rect 14365 22402 14431 22405
rect 25773 22402 25839 22405
rect 27245 22402 27311 22405
rect 14365 22400 22110 22402
rect 14365 22344 14370 22400
rect 14426 22344 22110 22400
rect 14365 22342 22110 22344
rect 14365 22339 14431 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 8385 22130 8451 22133
rect 12249 22130 12315 22133
rect 8385 22128 12315 22130
rect 8385 22072 8390 22128
rect 8446 22072 12254 22128
rect 12310 22072 12315 22128
rect 8385 22070 12315 22072
rect 8385 22067 8451 22070
rect 12249 22067 12315 22070
rect 12525 22130 12591 22133
rect 22050 22130 22110 22342
rect 25773 22400 27311 22402
rect 25773 22344 25778 22400
rect 25834 22344 27250 22400
rect 27306 22344 27311 22400
rect 25773 22342 27311 22344
rect 25773 22339 25839 22342
rect 27245 22339 27311 22342
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 27153 22266 27219 22269
rect 32121 22266 32187 22269
rect 27153 22264 32187 22266
rect 27153 22208 27158 22264
rect 27214 22208 32126 22264
rect 32182 22208 32187 22264
rect 27153 22206 32187 22208
rect 27153 22203 27219 22206
rect 32121 22203 32187 22206
rect 27521 22130 27587 22133
rect 12525 22128 16590 22130
rect 12525 22072 12530 22128
rect 12586 22072 16590 22128
rect 12525 22070 16590 22072
rect 22050 22128 27587 22130
rect 22050 22072 27526 22128
rect 27582 22072 27587 22128
rect 22050 22070 27587 22072
rect 12525 22067 12591 22070
rect 0 21994 800 22024
rect 4061 21994 4127 21997
rect 0 21992 4127 21994
rect 0 21936 4066 21992
rect 4122 21936 4127 21992
rect 0 21934 4127 21936
rect 0 21904 800 21934
rect 4061 21931 4127 21934
rect 8753 21994 8819 21997
rect 14549 21994 14615 21997
rect 8753 21992 14615 21994
rect 8753 21936 8758 21992
rect 8814 21936 14554 21992
rect 14610 21936 14615 21992
rect 8753 21934 14615 21936
rect 16530 21994 16590 22070
rect 27521 22067 27587 22070
rect 31937 22130 32003 22133
rect 32397 22130 32463 22133
rect 31937 22128 32463 22130
rect 31937 22072 31942 22128
rect 31998 22072 32402 22128
rect 32458 22072 32463 22128
rect 31937 22070 32463 22072
rect 31937 22067 32003 22070
rect 32397 22067 32463 22070
rect 35065 21994 35131 21997
rect 16530 21992 35131 21994
rect 16530 21936 35070 21992
rect 35126 21936 35131 21992
rect 16530 21934 35131 21936
rect 8753 21931 8819 21934
rect 14549 21931 14615 21934
rect 35065 21931 35131 21934
rect 49049 21994 49115 21997
rect 50200 21994 51000 22024
rect 49049 21992 51000 21994
rect 49049 21936 49054 21992
rect 49110 21936 51000 21992
rect 49049 21934 51000 21936
rect 49049 21931 49115 21934
rect 50200 21904 51000 21934
rect 20621 21858 20687 21861
rect 20621 21856 22110 21858
rect 20621 21800 20626 21856
rect 20682 21800 22110 21856
rect 20621 21798 22110 21800
rect 20621 21795 20687 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 22050 21722 22110 21798
rect 22686 21796 22692 21860
rect 22756 21858 22762 21860
rect 23289 21858 23355 21861
rect 22756 21856 23355 21858
rect 22756 21800 23294 21856
rect 23350 21800 23355 21856
rect 22756 21798 23355 21800
rect 22756 21796 22762 21798
rect 23289 21795 23355 21798
rect 23565 21858 23631 21861
rect 24945 21858 25011 21861
rect 23565 21856 25011 21858
rect 23565 21800 23570 21856
rect 23626 21800 24950 21856
rect 25006 21800 25011 21856
rect 23565 21798 25011 21800
rect 23565 21795 23631 21798
rect 24945 21795 25011 21798
rect 28625 21858 28691 21861
rect 29545 21858 29611 21861
rect 28625 21856 29611 21858
rect 28625 21800 28630 21856
rect 28686 21800 29550 21856
rect 29606 21800 29611 21856
rect 28625 21798 29611 21800
rect 28625 21795 28691 21798
rect 29545 21795 29611 21798
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 27061 21722 27127 21725
rect 22050 21720 27127 21722
rect 22050 21664 27066 21720
rect 27122 21664 27127 21720
rect 22050 21662 27127 21664
rect 27061 21659 27127 21662
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 3785 21586 3851 21589
rect 10501 21586 10567 21589
rect 3785 21584 10567 21586
rect 3785 21528 3790 21584
rect 3846 21528 10506 21584
rect 10562 21528 10567 21584
rect 3785 21526 10567 21528
rect 3785 21523 3851 21526
rect 10501 21523 10567 21526
rect 15929 21586 15995 21589
rect 36261 21586 36327 21589
rect 15929 21584 36327 21586
rect 15929 21528 15934 21584
rect 15990 21528 36266 21584
rect 36322 21528 36327 21584
rect 15929 21526 36327 21528
rect 15929 21523 15995 21526
rect 36261 21523 36327 21526
rect 1577 21450 1643 21453
rect 4286 21450 4292 21452
rect 1577 21448 4292 21450
rect 1577 21392 1582 21448
rect 1638 21392 4292 21448
rect 1577 21390 4292 21392
rect 1577 21387 1643 21390
rect 4286 21388 4292 21390
rect 4356 21388 4362 21452
rect 5206 21388 5212 21452
rect 5276 21450 5282 21452
rect 5533 21450 5599 21453
rect 5276 21448 5599 21450
rect 5276 21392 5538 21448
rect 5594 21392 5599 21448
rect 5276 21390 5599 21392
rect 5276 21388 5282 21390
rect 5533 21387 5599 21390
rect 7097 21450 7163 21453
rect 11145 21450 11211 21453
rect 12157 21450 12223 21453
rect 7097 21448 12223 21450
rect 7097 21392 7102 21448
rect 7158 21392 11150 21448
rect 11206 21392 12162 21448
rect 12218 21392 12223 21448
rect 7097 21390 12223 21392
rect 7097 21387 7163 21390
rect 11145 21387 11211 21390
rect 12157 21387 12223 21390
rect 15561 21450 15627 21453
rect 29821 21450 29887 21453
rect 15561 21448 29887 21450
rect 15561 21392 15566 21448
rect 15622 21392 29826 21448
rect 29882 21392 29887 21448
rect 15561 21390 29887 21392
rect 15561 21387 15627 21390
rect 29821 21387 29887 21390
rect 32673 21450 32739 21453
rect 33409 21450 33475 21453
rect 32673 21448 33475 21450
rect 32673 21392 32678 21448
rect 32734 21392 33414 21448
rect 33470 21392 33475 21448
rect 32673 21390 33475 21392
rect 32673 21387 32739 21390
rect 33409 21387 33475 21390
rect 5625 21314 5691 21317
rect 5758 21314 5764 21316
rect 5625 21312 5764 21314
rect 5625 21256 5630 21312
rect 5686 21256 5764 21312
rect 5625 21254 5764 21256
rect 5625 21251 5691 21254
rect 5758 21252 5764 21254
rect 5828 21314 5834 21316
rect 7557 21314 7623 21317
rect 5828 21312 7623 21314
rect 5828 21256 7562 21312
rect 7618 21256 7623 21312
rect 5828 21254 7623 21256
rect 5828 21252 5834 21254
rect 7557 21251 7623 21254
rect 13905 21314 13971 21317
rect 18597 21314 18663 21317
rect 13905 21312 18663 21314
rect 13905 21256 13910 21312
rect 13966 21256 18602 21312
rect 18658 21256 18663 21312
rect 13905 21254 18663 21256
rect 13905 21251 13971 21254
rect 18597 21251 18663 21254
rect 23473 21314 23539 21317
rect 27245 21314 27311 21317
rect 23473 21312 27311 21314
rect 23473 21256 23478 21312
rect 23534 21256 27250 21312
rect 27306 21256 27311 21312
rect 23473 21254 27311 21256
rect 23473 21251 23539 21254
rect 27245 21251 27311 21254
rect 27521 21314 27587 21317
rect 32765 21314 32831 21317
rect 27521 21312 32831 21314
rect 27521 21256 27526 21312
rect 27582 21256 32770 21312
rect 32826 21256 32831 21312
rect 27521 21254 32831 21256
rect 27521 21251 27587 21254
rect 32765 21251 32831 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 4286 21116 4292 21180
rect 4356 21178 4362 21180
rect 7925 21178 7991 21181
rect 4356 21176 7991 21178
rect 4356 21120 7930 21176
rect 7986 21120 7991 21176
rect 4356 21118 7991 21120
rect 4356 21116 4362 21118
rect 7925 21115 7991 21118
rect 16573 21178 16639 21181
rect 22737 21178 22803 21181
rect 32673 21178 32739 21181
rect 16573 21176 22803 21178
rect 16573 21120 16578 21176
rect 16634 21120 22742 21176
rect 22798 21120 22803 21176
rect 16573 21118 22803 21120
rect 16573 21115 16639 21118
rect 22737 21115 22803 21118
rect 26926 21176 32739 21178
rect 26926 21120 32678 21176
rect 32734 21120 32739 21176
rect 26926 21118 32739 21120
rect 4245 21042 4311 21045
rect 26926 21042 26986 21118
rect 32673 21115 32739 21118
rect 4245 21040 26986 21042
rect 4245 20984 4250 21040
rect 4306 20984 26986 21040
rect 4245 20982 26986 20984
rect 27061 21042 27127 21045
rect 34513 21042 34579 21045
rect 27061 21040 34579 21042
rect 27061 20984 27066 21040
rect 27122 20984 34518 21040
rect 34574 20984 34579 21040
rect 27061 20982 34579 20984
rect 4245 20979 4311 20982
rect 27061 20979 27127 20982
rect 34513 20979 34579 20982
rect 49141 21042 49207 21045
rect 50200 21042 51000 21072
rect 49141 21040 51000 21042
rect 49141 20984 49146 21040
rect 49202 20984 51000 21040
rect 49141 20982 51000 20984
rect 49141 20979 49207 20982
rect 50200 20952 51000 20982
rect 6453 20906 6519 20909
rect 11789 20906 11855 20909
rect 6453 20904 11855 20906
rect 6453 20848 6458 20904
rect 6514 20848 11794 20904
rect 11850 20848 11855 20904
rect 6453 20846 11855 20848
rect 6453 20843 6519 20846
rect 11789 20843 11855 20846
rect 17861 20906 17927 20909
rect 24209 20906 24275 20909
rect 40677 20906 40743 20909
rect 17861 20904 24275 20906
rect 17861 20848 17866 20904
rect 17922 20848 24214 20904
rect 24270 20848 24275 20904
rect 17861 20846 24275 20848
rect 17861 20843 17927 20846
rect 24209 20843 24275 20846
rect 24350 20904 40743 20906
rect 24350 20848 40682 20904
rect 40738 20848 40743 20904
rect 24350 20846 40743 20848
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 6913 20772 6979 20773
rect 6862 20770 6868 20772
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 6822 20710 6868 20770
rect 6932 20768 6979 20772
rect 6974 20712 6979 20768
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 6862 20708 6868 20710
rect 6932 20708 6979 20712
rect 11094 20708 11100 20772
rect 11164 20770 11170 20772
rect 11329 20770 11395 20773
rect 13905 20772 13971 20773
rect 11164 20768 11395 20770
rect 11164 20712 11334 20768
rect 11390 20712 11395 20768
rect 11164 20710 11395 20712
rect 11164 20708 11170 20710
rect 6913 20707 6979 20708
rect 11329 20707 11395 20710
rect 13854 20708 13860 20772
rect 13924 20770 13971 20772
rect 15745 20770 15811 20773
rect 15878 20770 15884 20772
rect 13924 20768 14016 20770
rect 13966 20712 14016 20768
rect 13924 20710 14016 20712
rect 15745 20768 15884 20770
rect 15745 20712 15750 20768
rect 15806 20712 15884 20768
rect 15745 20710 15884 20712
rect 13924 20708 13971 20710
rect 13905 20707 13971 20708
rect 15745 20707 15811 20710
rect 15878 20708 15884 20710
rect 15948 20708 15954 20772
rect 17166 20708 17172 20772
rect 17236 20770 17242 20772
rect 17769 20770 17835 20773
rect 17236 20768 17835 20770
rect 17236 20712 17774 20768
rect 17830 20712 17835 20768
rect 17236 20710 17835 20712
rect 17236 20708 17242 20710
rect 17769 20707 17835 20710
rect 22369 20770 22435 20773
rect 24350 20770 24410 20846
rect 40677 20843 40743 20846
rect 32121 20772 32187 20773
rect 22369 20768 24410 20770
rect 22369 20712 22374 20768
rect 22430 20712 24410 20768
rect 22369 20710 24410 20712
rect 22369 20707 22435 20710
rect 32070 20708 32076 20772
rect 32140 20770 32187 20772
rect 32140 20768 32232 20770
rect 32182 20712 32232 20768
rect 32140 20710 32232 20712
rect 32140 20708 32187 20710
rect 32622 20708 32628 20772
rect 32692 20770 32698 20772
rect 32857 20770 32923 20773
rect 32692 20768 32923 20770
rect 32692 20712 32862 20768
rect 32918 20712 32923 20768
rect 32692 20710 32923 20712
rect 32692 20708 32698 20710
rect 32121 20707 32187 20708
rect 32857 20707 32923 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 9581 20634 9647 20637
rect 16113 20634 16179 20637
rect 9581 20632 16179 20634
rect 9581 20576 9586 20632
rect 9642 20576 16118 20632
rect 16174 20576 16179 20632
rect 9581 20574 16179 20576
rect 9581 20571 9647 20574
rect 16113 20571 16179 20574
rect 23289 20634 23355 20637
rect 27061 20634 27127 20637
rect 23289 20632 27127 20634
rect 23289 20576 23294 20632
rect 23350 20576 27066 20632
rect 27122 20576 27127 20632
rect 23289 20574 27127 20576
rect 23289 20571 23355 20574
rect 27061 20571 27127 20574
rect 19977 20498 20043 20501
rect 36445 20498 36511 20501
rect 19977 20496 36511 20498
rect 19977 20440 19982 20496
rect 20038 20440 36450 20496
rect 36506 20440 36511 20496
rect 19977 20438 36511 20440
rect 19977 20435 20043 20438
rect 36445 20435 36511 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 13353 20362 13419 20365
rect 30097 20362 30163 20365
rect 13353 20360 30163 20362
rect 13353 20304 13358 20360
rect 13414 20304 30102 20360
rect 30158 20304 30163 20360
rect 13353 20302 30163 20304
rect 13353 20299 13419 20302
rect 30097 20299 30163 20302
rect 5625 20226 5691 20229
rect 6637 20226 6703 20229
rect 14273 20226 14339 20229
rect 17953 20226 18019 20229
rect 5625 20224 12450 20226
rect 5625 20168 5630 20224
rect 5686 20168 6642 20224
rect 6698 20168 12450 20224
rect 5625 20166 12450 20168
rect 5625 20163 5691 20166
rect 6637 20163 6703 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 7557 20092 7623 20093
rect 7557 20090 7604 20092
rect 7512 20088 7604 20090
rect 7512 20032 7562 20088
rect 7512 20030 7604 20032
rect 7557 20028 7604 20030
rect 7668 20028 7674 20092
rect 7557 20027 7623 20028
rect 0 19954 800 19984
rect 1945 19954 2011 19957
rect 0 19952 2011 19954
rect 0 19896 1950 19952
rect 2006 19896 2011 19952
rect 0 19894 2011 19896
rect 0 19864 800 19894
rect 1945 19891 2011 19894
rect 4245 19954 4311 19957
rect 11421 19954 11487 19957
rect 4245 19952 11487 19954
rect 4245 19896 4250 19952
rect 4306 19896 11426 19952
rect 11482 19896 11487 19952
rect 4245 19894 11487 19896
rect 12390 19954 12450 20166
rect 14273 20224 18019 20226
rect 14273 20168 14278 20224
rect 14334 20168 17958 20224
rect 18014 20168 18019 20224
rect 14273 20166 18019 20168
rect 14273 20163 14339 20166
rect 17953 20163 18019 20166
rect 27153 20226 27219 20229
rect 28717 20226 28783 20229
rect 27153 20224 28783 20226
rect 27153 20168 27158 20224
rect 27214 20168 28722 20224
rect 28778 20168 28783 20224
rect 27153 20166 28783 20168
rect 27153 20163 27219 20166
rect 28717 20163 28783 20166
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 18597 20090 18663 20093
rect 16990 20088 18663 20090
rect 16990 20032 18602 20088
rect 18658 20032 18663 20088
rect 16990 20030 18663 20032
rect 16990 19954 17050 20030
rect 18597 20027 18663 20030
rect 25957 20090 26023 20093
rect 30833 20090 30899 20093
rect 32305 20090 32371 20093
rect 25957 20088 30899 20090
rect 25957 20032 25962 20088
rect 26018 20032 30838 20088
rect 30894 20032 30899 20088
rect 25957 20030 30899 20032
rect 25957 20027 26023 20030
rect 30833 20027 30899 20030
rect 31710 20088 32371 20090
rect 31710 20032 32310 20088
rect 32366 20032 32371 20088
rect 31710 20030 32371 20032
rect 12390 19894 17050 19954
rect 17217 19954 17283 19957
rect 28993 19954 29059 19957
rect 17217 19952 29059 19954
rect 17217 19896 17222 19952
rect 17278 19896 28998 19952
rect 29054 19896 29059 19952
rect 17217 19894 29059 19896
rect 4245 19891 4311 19894
rect 11421 19891 11487 19894
rect 17217 19891 17283 19894
rect 28993 19891 29059 19894
rect 11789 19818 11855 19821
rect 31710 19818 31770 20030
rect 32305 20027 32371 20030
rect 11789 19816 31770 19818
rect 11789 19760 11794 19816
rect 11850 19760 31770 19816
rect 11789 19758 31770 19760
rect 11789 19755 11855 19758
rect 3877 19682 3943 19685
rect 7046 19682 7052 19684
rect 3877 19680 7052 19682
rect 3877 19624 3882 19680
rect 3938 19624 7052 19680
rect 3877 19622 7052 19624
rect 3877 19619 3943 19622
rect 7046 19620 7052 19622
rect 7116 19620 7122 19684
rect 18597 19682 18663 19685
rect 27613 19682 27679 19685
rect 18597 19680 27679 19682
rect 18597 19624 18602 19680
rect 18658 19624 27618 19680
rect 27674 19624 27679 19680
rect 18597 19622 27679 19624
rect 18597 19619 18663 19622
rect 27613 19619 27679 19622
rect 29821 19682 29887 19685
rect 30741 19682 30807 19685
rect 29821 19680 30807 19682
rect 29821 19624 29826 19680
rect 29882 19624 30746 19680
rect 30802 19624 30807 19680
rect 29821 19622 30807 19624
rect 29821 19619 29887 19622
rect 30741 19619 30807 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2773 19546 2839 19549
rect 0 19544 2839 19546
rect 0 19488 2778 19544
rect 2834 19488 2839 19544
rect 0 19486 2839 19488
rect 0 19456 800 19486
rect 2773 19483 2839 19486
rect 9765 19546 9831 19549
rect 13721 19546 13787 19549
rect 9765 19544 13787 19546
rect 9765 19488 9770 19544
rect 9826 19488 13726 19544
rect 13782 19488 13787 19544
rect 9765 19486 13787 19488
rect 9765 19483 9831 19486
rect 13721 19483 13787 19486
rect 19333 19546 19399 19549
rect 25957 19546 26023 19549
rect 19333 19544 26023 19546
rect 19333 19488 19338 19544
rect 19394 19488 25962 19544
rect 26018 19488 26023 19544
rect 19333 19486 26023 19488
rect 19333 19483 19399 19486
rect 25957 19483 26023 19486
rect 5717 19410 5783 19413
rect 6453 19410 6519 19413
rect 5717 19408 6519 19410
rect 5717 19352 5722 19408
rect 5778 19352 6458 19408
rect 6514 19352 6519 19408
rect 5717 19350 6519 19352
rect 5717 19347 5783 19350
rect 6453 19347 6519 19350
rect 11881 19410 11947 19413
rect 30649 19410 30715 19413
rect 11881 19408 30715 19410
rect 11881 19352 11886 19408
rect 11942 19352 30654 19408
rect 30710 19352 30715 19408
rect 11881 19350 30715 19352
rect 11881 19347 11947 19350
rect 30649 19347 30715 19350
rect 30833 19410 30899 19413
rect 43437 19410 43503 19413
rect 30833 19408 43503 19410
rect 30833 19352 30838 19408
rect 30894 19352 43442 19408
rect 43498 19352 43503 19408
rect 30833 19350 43503 19352
rect 30833 19347 30899 19350
rect 43437 19347 43503 19350
rect 3601 19274 3667 19277
rect 3601 19272 8218 19274
rect 3601 19216 3606 19272
rect 3662 19216 8218 19272
rect 3601 19214 8218 19216
rect 3601 19211 3667 19214
rect 0 19138 800 19168
rect 2037 19138 2103 19141
rect 0 19136 2103 19138
rect 0 19080 2042 19136
rect 2098 19080 2103 19136
rect 0 19078 2103 19080
rect 0 19048 800 19078
rect 2037 19075 2103 19078
rect 3785 19138 3851 19141
rect 4337 19138 4403 19141
rect 3785 19136 4403 19138
rect 3785 19080 3790 19136
rect 3846 19080 4342 19136
rect 4398 19080 4403 19136
rect 3785 19078 4403 19080
rect 8158 19138 8218 19214
rect 8334 19212 8340 19276
rect 8404 19274 8410 19276
rect 9949 19274 10015 19277
rect 26969 19274 27035 19277
rect 8404 19272 27035 19274
rect 8404 19216 9954 19272
rect 10010 19216 26974 19272
rect 27030 19216 27035 19272
rect 8404 19214 27035 19216
rect 8404 19212 8410 19214
rect 9949 19211 10015 19214
rect 26969 19211 27035 19214
rect 13721 19138 13787 19141
rect 18689 19138 18755 19141
rect 8158 19078 11530 19138
rect 3785 19075 3851 19078
rect 4337 19075 4403 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 4705 19002 4771 19005
rect 9397 19002 9463 19005
rect 4705 19000 9463 19002
rect 4705 18944 4710 19000
rect 4766 18944 9402 19000
rect 9458 18944 9463 19000
rect 4705 18942 9463 18944
rect 4705 18939 4771 18942
rect 9397 18939 9463 18942
rect 1761 18866 1827 18869
rect 11329 18866 11395 18869
rect 1761 18864 11395 18866
rect 1761 18808 1766 18864
rect 1822 18808 11334 18864
rect 11390 18808 11395 18864
rect 1761 18806 11395 18808
rect 1761 18803 1827 18806
rect 11329 18803 11395 18806
rect 0 18730 800 18760
rect 2865 18730 2931 18733
rect 0 18728 2931 18730
rect 0 18672 2870 18728
rect 2926 18672 2931 18728
rect 0 18670 2931 18672
rect 0 18640 800 18670
rect 2865 18667 2931 18670
rect 3601 18730 3667 18733
rect 3734 18730 3740 18732
rect 3601 18728 3740 18730
rect 3601 18672 3606 18728
rect 3662 18672 3740 18728
rect 3601 18670 3740 18672
rect 3601 18667 3667 18670
rect 3734 18668 3740 18670
rect 3804 18668 3810 18732
rect 7465 18730 7531 18733
rect 8569 18730 8635 18733
rect 7465 18728 8635 18730
rect 7465 18672 7470 18728
rect 7526 18672 8574 18728
rect 8630 18672 8635 18728
rect 7465 18670 8635 18672
rect 7465 18667 7531 18670
rect 8569 18667 8635 18670
rect 11470 18594 11530 19078
rect 13721 19136 18755 19138
rect 13721 19080 13726 19136
rect 13782 19080 18694 19136
rect 18750 19080 18755 19136
rect 13721 19078 18755 19080
rect 13721 19075 13787 19078
rect 18689 19075 18755 19078
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 13445 19002 13511 19005
rect 14406 19002 14412 19004
rect 13445 19000 14412 19002
rect 13445 18944 13450 19000
rect 13506 18944 14412 19000
rect 13445 18942 14412 18944
rect 13445 18939 13511 18942
rect 14406 18940 14412 18942
rect 14476 19002 14482 19004
rect 18597 19002 18663 19005
rect 22737 19002 22803 19005
rect 14476 19000 22803 19002
rect 14476 18944 18602 19000
rect 18658 18944 22742 19000
rect 22798 18944 22803 19000
rect 14476 18942 22803 18944
rect 14476 18940 14482 18942
rect 18597 18939 18663 18942
rect 22737 18939 22803 18942
rect 25129 19002 25195 19005
rect 25129 19000 31770 19002
rect 25129 18944 25134 19000
rect 25190 18944 31770 19000
rect 25129 18942 31770 18944
rect 25129 18939 25195 18942
rect 14457 18866 14523 18869
rect 15193 18866 15259 18869
rect 14457 18864 15259 18866
rect 14457 18808 14462 18864
rect 14518 18808 15198 18864
rect 15254 18808 15259 18864
rect 14457 18806 15259 18808
rect 14457 18803 14523 18806
rect 15193 18803 15259 18806
rect 15377 18866 15443 18869
rect 22461 18866 22527 18869
rect 15377 18864 22527 18866
rect 15377 18808 15382 18864
rect 15438 18808 22466 18864
rect 22522 18808 22527 18864
rect 15377 18806 22527 18808
rect 15377 18803 15443 18806
rect 22461 18803 22527 18806
rect 25865 18866 25931 18869
rect 31710 18866 31770 18942
rect 45369 18866 45435 18869
rect 25865 18864 27170 18866
rect 25865 18808 25870 18864
rect 25926 18808 27170 18864
rect 25865 18806 27170 18808
rect 31710 18864 45435 18866
rect 31710 18808 45374 18864
rect 45430 18808 45435 18864
rect 31710 18806 45435 18808
rect 25865 18803 25931 18806
rect 11881 18730 11947 18733
rect 27110 18730 27170 18806
rect 45369 18803 45435 18806
rect 45737 18730 45803 18733
rect 11881 18728 26986 18730
rect 11881 18672 11886 18728
rect 11942 18672 26986 18728
rect 11881 18670 26986 18672
rect 27110 18728 45803 18730
rect 27110 18672 45742 18728
rect 45798 18672 45803 18728
rect 27110 18670 45803 18672
rect 11881 18667 11947 18670
rect 13721 18594 13787 18597
rect 11470 18592 13787 18594
rect 11470 18536 13726 18592
rect 13782 18536 13787 18592
rect 11470 18534 13787 18536
rect 13721 18531 13787 18534
rect 22737 18594 22803 18597
rect 24761 18594 24827 18597
rect 22737 18592 24827 18594
rect 22737 18536 22742 18592
rect 22798 18536 24766 18592
rect 24822 18536 24827 18592
rect 22737 18534 24827 18536
rect 22737 18531 22803 18534
rect 24761 18531 24827 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 15101 18458 15167 18461
rect 19977 18458 20043 18461
rect 24025 18458 24091 18461
rect 12390 18456 15167 18458
rect 12390 18400 15106 18456
rect 15162 18400 15167 18456
rect 12390 18398 15167 18400
rect 0 18322 800 18352
rect 2773 18322 2839 18325
rect 0 18320 2839 18322
rect 0 18264 2778 18320
rect 2834 18264 2839 18320
rect 0 18262 2839 18264
rect 0 18232 800 18262
rect 2773 18259 2839 18262
rect 4245 18322 4311 18325
rect 12390 18322 12450 18398
rect 15101 18395 15167 18398
rect 18462 18456 24091 18458
rect 18462 18400 19982 18456
rect 20038 18400 24030 18456
rect 24086 18400 24091 18456
rect 18462 18398 24091 18400
rect 4245 18320 12450 18322
rect 4245 18264 4250 18320
rect 4306 18264 12450 18320
rect 4245 18262 12450 18264
rect 4245 18259 4311 18262
rect 12750 18260 12756 18324
rect 12820 18322 12826 18324
rect 13353 18322 13419 18325
rect 12820 18320 13419 18322
rect 12820 18264 13358 18320
rect 13414 18264 13419 18320
rect 12820 18262 13419 18264
rect 12820 18260 12826 18262
rect 13353 18259 13419 18262
rect 14181 18322 14247 18325
rect 16481 18322 16547 18325
rect 18462 18322 18522 18398
rect 19977 18395 20043 18398
rect 24025 18395 24091 18398
rect 14181 18320 18522 18322
rect 14181 18264 14186 18320
rect 14242 18264 16486 18320
rect 16542 18264 18522 18320
rect 14181 18262 18522 18264
rect 26926 18322 26986 18670
rect 45737 18667 45803 18670
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 32070 18322 32076 18324
rect 26926 18262 32076 18322
rect 14181 18259 14247 18262
rect 16481 18259 16547 18262
rect 32070 18260 32076 18262
rect 32140 18260 32146 18324
rect 5349 18186 5415 18189
rect 7557 18186 7623 18189
rect 5349 18184 7623 18186
rect 5349 18128 5354 18184
rect 5410 18128 7562 18184
rect 7618 18128 7623 18184
rect 5349 18126 7623 18128
rect 5349 18123 5415 18126
rect 7557 18123 7623 18126
rect 11421 18186 11487 18189
rect 13997 18186 14063 18189
rect 11421 18184 14063 18186
rect 11421 18128 11426 18184
rect 11482 18128 14002 18184
rect 14058 18128 14063 18184
rect 11421 18126 14063 18128
rect 11421 18123 11487 18126
rect 13997 18123 14063 18126
rect 15009 18186 15075 18189
rect 27613 18186 27679 18189
rect 15009 18184 27679 18186
rect 15009 18128 15014 18184
rect 15070 18128 27618 18184
rect 27674 18128 27679 18184
rect 15009 18126 27679 18128
rect 15009 18123 15075 18126
rect 27613 18123 27679 18126
rect 5625 18052 5691 18053
rect 5574 18050 5580 18052
rect 5534 17990 5580 18050
rect 5644 18048 5691 18052
rect 5686 17992 5691 18048
rect 5574 17988 5580 17990
rect 5644 17988 5691 17992
rect 5625 17987 5691 17988
rect 9121 18050 9187 18053
rect 9489 18050 9555 18053
rect 9121 18048 9555 18050
rect 9121 17992 9126 18048
rect 9182 17992 9494 18048
rect 9550 17992 9555 18048
rect 9121 17990 9555 17992
rect 9121 17987 9187 17990
rect 9489 17987 9555 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 3785 17914 3851 17917
rect 10409 17914 10475 17917
rect 3785 17912 10475 17914
rect 3785 17856 3790 17912
rect 3846 17856 10414 17912
rect 10470 17856 10475 17912
rect 3785 17854 10475 17856
rect 3785 17851 3851 17854
rect 10409 17851 10475 17854
rect 14825 17914 14891 17917
rect 20069 17914 20135 17917
rect 14825 17912 20135 17914
rect 14825 17856 14830 17912
rect 14886 17856 20074 17912
rect 20130 17856 20135 17912
rect 14825 17854 20135 17856
rect 14825 17851 14891 17854
rect 20069 17851 20135 17854
rect 25405 17914 25471 17917
rect 27429 17914 27495 17917
rect 25405 17912 27495 17914
rect 25405 17856 25410 17912
rect 25466 17856 27434 17912
rect 27490 17856 27495 17912
rect 25405 17854 27495 17856
rect 25405 17851 25471 17854
rect 27429 17851 27495 17854
rect 4889 17778 4955 17781
rect 5901 17778 5967 17781
rect 4889 17776 5967 17778
rect 4889 17720 4894 17776
rect 4950 17720 5906 17776
rect 5962 17720 5967 17776
rect 4889 17718 5967 17720
rect 4889 17715 4955 17718
rect 5901 17715 5967 17718
rect 7046 17716 7052 17780
rect 7116 17778 7122 17780
rect 7281 17778 7347 17781
rect 11646 17778 11652 17780
rect 7116 17776 11652 17778
rect 7116 17720 7286 17776
rect 7342 17720 11652 17776
rect 7116 17718 11652 17720
rect 7116 17716 7122 17718
rect 7281 17715 7347 17718
rect 11646 17716 11652 17718
rect 11716 17716 11722 17780
rect 12566 17716 12572 17780
rect 12636 17778 12642 17780
rect 16481 17778 16547 17781
rect 33501 17778 33567 17781
rect 12636 17776 16547 17778
rect 12636 17720 16486 17776
rect 16542 17720 16547 17776
rect 12636 17718 16547 17720
rect 12636 17716 12642 17718
rect 16481 17715 16547 17718
rect 16622 17776 33567 17778
rect 16622 17720 33506 17776
rect 33562 17720 33567 17776
rect 16622 17718 33567 17720
rect 7097 17642 7163 17645
rect 14457 17642 14523 17645
rect 7097 17640 14523 17642
rect 7097 17584 7102 17640
rect 7158 17584 14462 17640
rect 14518 17584 14523 17640
rect 7097 17582 14523 17584
rect 7097 17579 7163 17582
rect 14457 17579 14523 17582
rect 16205 17642 16271 17645
rect 16622 17642 16682 17718
rect 33501 17715 33567 17718
rect 19701 17642 19767 17645
rect 16205 17640 16682 17642
rect 16205 17584 16210 17640
rect 16266 17584 16682 17640
rect 16205 17582 16682 17584
rect 17726 17640 19767 17642
rect 17726 17584 19706 17640
rect 19762 17584 19767 17640
rect 17726 17582 19767 17584
rect 16205 17579 16271 17582
rect 0 17506 800 17536
rect 2037 17506 2103 17509
rect 0 17504 2103 17506
rect 0 17448 2042 17504
rect 2098 17448 2103 17504
rect 0 17446 2103 17448
rect 0 17416 800 17446
rect 2037 17443 2103 17446
rect 12157 17506 12223 17509
rect 12801 17506 12867 17509
rect 12157 17504 12867 17506
rect 12157 17448 12162 17504
rect 12218 17448 12806 17504
rect 12862 17448 12867 17504
rect 12157 17446 12867 17448
rect 12157 17443 12223 17446
rect 12801 17443 12867 17446
rect 12985 17506 13051 17509
rect 17726 17506 17786 17582
rect 19701 17579 19767 17582
rect 24025 17642 24091 17645
rect 30189 17642 30255 17645
rect 24025 17640 30255 17642
rect 24025 17584 24030 17640
rect 24086 17584 30194 17640
rect 30250 17584 30255 17640
rect 24025 17582 30255 17584
rect 24025 17579 24091 17582
rect 30189 17579 30255 17582
rect 12985 17504 17786 17506
rect 12985 17448 12990 17504
rect 13046 17448 17786 17504
rect 12985 17446 17786 17448
rect 12985 17443 13051 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 2497 17370 2563 17373
rect 7741 17370 7807 17373
rect 2497 17368 7807 17370
rect 2497 17312 2502 17368
rect 2558 17312 7746 17368
rect 7802 17312 7807 17368
rect 2497 17310 7807 17312
rect 2497 17307 2563 17310
rect 7741 17307 7807 17310
rect 8569 17370 8635 17373
rect 12382 17370 12388 17372
rect 8569 17368 12388 17370
rect 8569 17312 8574 17368
rect 8630 17312 12388 17368
rect 8569 17310 12388 17312
rect 8569 17307 8635 17310
rect 12382 17308 12388 17310
rect 12452 17308 12458 17372
rect 18781 17370 18847 17373
rect 21449 17370 21515 17373
rect 12574 17310 17786 17370
rect 3417 17234 3483 17237
rect 8385 17234 8451 17237
rect 11053 17234 11119 17237
rect 12574 17234 12634 17310
rect 2730 17232 8451 17234
rect 2730 17176 3422 17232
rect 3478 17176 8390 17232
rect 8446 17176 8451 17232
rect 2730 17174 8451 17176
rect 0 17098 800 17128
rect 2730 17101 2790 17174
rect 3417 17171 3483 17174
rect 8385 17171 8451 17174
rect 9630 17174 10242 17234
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 2681 17096 2790 17101
rect 2681 17040 2686 17096
rect 2742 17040 2790 17096
rect 2681 17038 2790 17040
rect 6453 17098 6519 17101
rect 8201 17098 8267 17101
rect 9630 17098 9690 17174
rect 9857 17100 9923 17101
rect 6453 17096 9690 17098
rect 6453 17040 6458 17096
rect 6514 17040 8206 17096
rect 8262 17040 9690 17096
rect 6453 17038 9690 17040
rect 2681 17035 2747 17038
rect 6453 17035 6519 17038
rect 8201 17035 8267 17038
rect 9806 17036 9812 17100
rect 9876 17098 9923 17100
rect 10182 17098 10242 17174
rect 11053 17232 12634 17234
rect 11053 17176 11058 17232
rect 11114 17176 12634 17232
rect 11053 17174 12634 17176
rect 17726 17234 17786 17310
rect 18781 17368 21515 17370
rect 18781 17312 18786 17368
rect 18842 17312 21454 17368
rect 21510 17312 21515 17368
rect 18781 17310 21515 17312
rect 18781 17307 18847 17310
rect 21449 17307 21515 17310
rect 18965 17234 19031 17237
rect 17726 17232 19031 17234
rect 17726 17176 18970 17232
rect 19026 17176 19031 17232
rect 17726 17174 19031 17176
rect 11053 17171 11119 17174
rect 18965 17171 19031 17174
rect 20621 17234 20687 17237
rect 21081 17234 21147 17237
rect 21633 17234 21699 17237
rect 20621 17232 21699 17234
rect 20621 17176 20626 17232
rect 20682 17176 21086 17232
rect 21142 17176 21638 17232
rect 21694 17176 21699 17232
rect 20621 17174 21699 17176
rect 20621 17171 20687 17174
rect 21081 17171 21147 17174
rect 21633 17171 21699 17174
rect 31201 17098 31267 17101
rect 9876 17096 9968 17098
rect 9918 17040 9968 17096
rect 9876 17038 9968 17040
rect 10182 17096 31267 17098
rect 10182 17040 31206 17096
rect 31262 17040 31267 17096
rect 10182 17038 31267 17040
rect 9876 17036 9923 17038
rect 9857 17035 9923 17036
rect 31201 17035 31267 17038
rect 4429 16962 4495 16965
rect 4429 16960 12450 16962
rect 4429 16904 4434 16960
rect 4490 16904 12450 16960
rect 4429 16902 12450 16904
rect 4429 16899 4495 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 3601 16826 3667 16829
rect 8569 16826 8635 16829
rect 3601 16824 8635 16826
rect 3601 16768 3606 16824
rect 3662 16768 8574 16824
rect 8630 16768 8635 16824
rect 3601 16766 8635 16768
rect 3601 16763 3667 16766
rect 8569 16763 8635 16766
rect 10409 16826 10475 16829
rect 10869 16826 10935 16829
rect 10409 16824 10935 16826
rect 10409 16768 10414 16824
rect 10470 16768 10874 16824
rect 10930 16768 10935 16824
rect 10409 16766 10935 16768
rect 12390 16826 12450 16902
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 12617 16826 12683 16829
rect 12390 16824 12683 16826
rect 12390 16768 12622 16824
rect 12678 16768 12683 16824
rect 12390 16766 12683 16768
rect 10409 16763 10475 16766
rect 10869 16763 10935 16766
rect 12617 16763 12683 16766
rect 16481 16826 16547 16829
rect 18781 16826 18847 16829
rect 16481 16824 22110 16826
rect 16481 16768 16486 16824
rect 16542 16768 18786 16824
rect 18842 16768 22110 16824
rect 16481 16766 22110 16768
rect 16481 16763 16547 16766
rect 18781 16763 18847 16766
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 5901 16690 5967 16693
rect 8109 16690 8175 16693
rect 5901 16688 8175 16690
rect 5901 16632 5906 16688
rect 5962 16632 8114 16688
rect 8170 16632 8175 16688
rect 5901 16630 8175 16632
rect 5901 16627 5967 16630
rect 8109 16627 8175 16630
rect 10777 16690 10843 16693
rect 21265 16690 21331 16693
rect 10777 16688 21331 16690
rect 10777 16632 10782 16688
rect 10838 16632 21270 16688
rect 21326 16632 21331 16688
rect 10777 16630 21331 16632
rect 22050 16690 22110 16766
rect 23841 16690 23907 16693
rect 22050 16688 23907 16690
rect 22050 16632 23846 16688
rect 23902 16632 23907 16688
rect 22050 16630 23907 16632
rect 10777 16627 10843 16630
rect 21265 16627 21331 16630
rect 23841 16627 23907 16630
rect 5073 16554 5139 16557
rect 11145 16554 11211 16557
rect 5073 16552 11211 16554
rect 5073 16496 5078 16552
rect 5134 16496 11150 16552
rect 11206 16496 11211 16552
rect 5073 16494 11211 16496
rect 5073 16491 5139 16494
rect 11145 16491 11211 16494
rect 11605 16554 11671 16557
rect 13813 16554 13879 16557
rect 11605 16552 13879 16554
rect 11605 16496 11610 16552
rect 11666 16496 13818 16552
rect 13874 16496 13879 16552
rect 11605 16494 13879 16496
rect 11605 16491 11671 16494
rect 13813 16491 13879 16494
rect 14365 16554 14431 16557
rect 28349 16554 28415 16557
rect 14365 16552 28415 16554
rect 14365 16496 14370 16552
rect 14426 16496 28354 16552
rect 28410 16496 28415 16552
rect 14365 16494 28415 16496
rect 14365 16491 14431 16494
rect 28349 16491 28415 16494
rect 9765 16418 9831 16421
rect 10501 16418 10567 16421
rect 16205 16418 16271 16421
rect 9765 16416 10567 16418
rect 9765 16360 9770 16416
rect 9826 16360 10506 16416
rect 10562 16360 10567 16416
rect 9765 16358 10567 16360
rect 9765 16355 9831 16358
rect 10501 16355 10567 16358
rect 11424 16416 16271 16418
rect 11424 16360 16210 16416
rect 16266 16360 16271 16416
rect 11424 16358 16271 16360
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 8845 16282 8911 16285
rect 10685 16282 10751 16285
rect 11424 16282 11484 16358
rect 16205 16355 16271 16358
rect 19333 16418 19399 16421
rect 26141 16418 26207 16421
rect 19333 16416 26207 16418
rect 19333 16360 19338 16416
rect 19394 16360 26146 16416
rect 26202 16360 26207 16416
rect 19333 16358 26207 16360
rect 19333 16355 19399 16358
rect 26141 16355 26207 16358
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 11605 16284 11671 16285
rect 17125 16284 17191 16285
rect 11605 16282 11652 16284
rect 8845 16280 11484 16282
rect 8845 16224 8850 16280
rect 8906 16224 10690 16280
rect 10746 16224 11484 16280
rect 8845 16222 11484 16224
rect 11560 16280 11652 16282
rect 11560 16224 11610 16280
rect 11560 16222 11652 16224
rect 8845 16219 8911 16222
rect 10685 16219 10751 16222
rect 11605 16220 11652 16222
rect 11716 16220 11722 16284
rect 17125 16282 17172 16284
rect 17080 16280 17172 16282
rect 17080 16224 17130 16280
rect 17080 16222 17172 16224
rect 17125 16220 17172 16222
rect 17236 16220 17242 16284
rect 11605 16219 11671 16220
rect 17125 16219 17191 16220
rect 3877 16146 3943 16149
rect 9765 16146 9831 16149
rect 3877 16144 9831 16146
rect 3877 16088 3882 16144
rect 3938 16088 9770 16144
rect 9826 16088 9831 16144
rect 3877 16086 9831 16088
rect 3877 16083 3943 16086
rect 9765 16083 9831 16086
rect 16941 16146 17007 16149
rect 18454 16146 18460 16148
rect 16941 16144 18460 16146
rect 16941 16088 16946 16144
rect 17002 16088 18460 16144
rect 16941 16086 18460 16088
rect 16941 16083 17007 16086
rect 18454 16084 18460 16086
rect 18524 16084 18530 16148
rect 21265 16146 21331 16149
rect 24761 16146 24827 16149
rect 21265 16144 24827 16146
rect 21265 16088 21270 16144
rect 21326 16088 24766 16144
rect 24822 16088 24827 16144
rect 21265 16086 24827 16088
rect 21265 16083 21331 16086
rect 24761 16083 24827 16086
rect 3969 16010 4035 16013
rect 7925 16010 7991 16013
rect 8518 16010 8524 16012
rect 3969 16008 8524 16010
rect 3969 15952 3974 16008
rect 4030 15952 7930 16008
rect 7986 15952 8524 16008
rect 3969 15950 8524 15952
rect 3969 15947 4035 15950
rect 7925 15947 7991 15950
rect 8518 15948 8524 15950
rect 8588 15948 8594 16012
rect 10961 16010 11027 16013
rect 30097 16010 30163 16013
rect 10961 16008 30163 16010
rect 10961 15952 10966 16008
rect 11022 15952 30102 16008
rect 30158 15952 30163 16008
rect 10961 15950 30163 15952
rect 10961 15947 11027 15950
rect 30097 15947 30163 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 9673 15738 9739 15741
rect 12249 15738 12315 15741
rect 9673 15736 12315 15738
rect 9673 15680 9678 15736
rect 9734 15680 12254 15736
rect 12310 15680 12315 15736
rect 9673 15678 12315 15680
rect 9673 15675 9739 15678
rect 12249 15675 12315 15678
rect 13721 15738 13787 15741
rect 21541 15738 21607 15741
rect 13721 15736 21607 15738
rect 13721 15680 13726 15736
rect 13782 15680 21546 15736
rect 21602 15680 21607 15736
rect 13721 15678 21607 15680
rect 13721 15675 13787 15678
rect 21541 15675 21607 15678
rect 12065 15602 12131 15605
rect 29913 15602 29979 15605
rect 12065 15600 29979 15602
rect 12065 15544 12070 15600
rect 12126 15544 29918 15600
rect 29974 15544 29979 15600
rect 12065 15542 29979 15544
rect 12065 15539 12131 15542
rect 29913 15539 29979 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 9581 15466 9647 15469
rect 9949 15466 10015 15469
rect 32029 15466 32095 15469
rect 9581 15464 10015 15466
rect 9581 15408 9586 15464
rect 9642 15408 9954 15464
rect 10010 15408 10015 15464
rect 9581 15406 10015 15408
rect 9581 15403 9647 15406
rect 9949 15403 10015 15406
rect 10182 15464 32095 15466
rect 10182 15408 32034 15464
rect 32090 15408 32095 15464
rect 10182 15406 32095 15408
rect 8477 15330 8543 15333
rect 10182 15330 10242 15406
rect 32029 15403 32095 15406
rect 8477 15328 10242 15330
rect 8477 15272 8482 15328
rect 8538 15272 10242 15328
rect 8477 15270 10242 15272
rect 11421 15330 11487 15333
rect 12617 15330 12683 15333
rect 11421 15328 12683 15330
rect 11421 15272 11426 15328
rect 11482 15272 12622 15328
rect 12678 15272 12683 15328
rect 11421 15270 12683 15272
rect 8477 15267 8543 15270
rect 11421 15267 11487 15270
rect 12617 15267 12683 15270
rect 20069 15330 20135 15333
rect 20069 15328 20178 15330
rect 20069 15272 20074 15328
rect 20130 15272 20178 15328
rect 20069 15267 20178 15272
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 5441 15194 5507 15197
rect 7097 15194 7163 15197
rect 5441 15192 7163 15194
rect 5441 15136 5446 15192
rect 5502 15136 7102 15192
rect 7158 15136 7163 15192
rect 5441 15134 7163 15136
rect 5441 15131 5507 15134
rect 7097 15131 7163 15134
rect 8385 15194 8451 15197
rect 11421 15194 11487 15197
rect 13813 15194 13879 15197
rect 8385 15192 13879 15194
rect 8385 15136 8390 15192
rect 8446 15136 11426 15192
rect 11482 15136 13818 15192
rect 13874 15136 13879 15192
rect 8385 15134 13879 15136
rect 8385 15131 8451 15134
rect 11421 15131 11487 15134
rect 13813 15131 13879 15134
rect 18505 15194 18571 15197
rect 20118 15194 20178 15267
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 25589 15194 25655 15197
rect 18505 15192 25655 15194
rect 18505 15136 18510 15192
rect 18566 15136 25594 15192
rect 25650 15136 25655 15192
rect 18505 15134 25655 15136
rect 18505 15131 18571 15134
rect 25589 15131 25655 15134
rect 0 15058 800 15088
rect 1117 15058 1183 15061
rect 0 15056 1183 15058
rect 0 15000 1122 15056
rect 1178 15000 1183 15056
rect 0 14998 1183 15000
rect 0 14968 800 14998
rect 1117 14995 1183 14998
rect 5717 15058 5783 15061
rect 6637 15058 6703 15061
rect 5717 15056 6703 15058
rect 5717 15000 5722 15056
rect 5778 15000 6642 15056
rect 6698 15000 6703 15056
rect 5717 14998 6703 15000
rect 5717 14995 5783 14998
rect 6637 14995 6703 14998
rect 11973 15058 12039 15061
rect 34053 15058 34119 15061
rect 11973 15056 34119 15058
rect 11973 15000 11978 15056
rect 12034 15000 34058 15056
rect 34114 15000 34119 15056
rect 11973 14998 34119 15000
rect 11973 14995 12039 14998
rect 34053 14995 34119 14998
rect 5901 14922 5967 14925
rect 7373 14922 7439 14925
rect 7925 14922 7991 14925
rect 17125 14922 17191 14925
rect 19333 14922 19399 14925
rect 5901 14920 9690 14922
rect 5901 14864 5906 14920
rect 5962 14864 7378 14920
rect 7434 14864 7930 14920
rect 7986 14864 9690 14920
rect 5901 14862 9690 14864
rect 5901 14859 5967 14862
rect 7373 14859 7439 14862
rect 7925 14859 7991 14862
rect 9630 14786 9690 14862
rect 17125 14920 19399 14922
rect 17125 14864 17130 14920
rect 17186 14864 19338 14920
rect 19394 14864 19399 14920
rect 17125 14862 19399 14864
rect 17125 14859 17191 14862
rect 19333 14859 19399 14862
rect 19977 14922 20043 14925
rect 22277 14922 22343 14925
rect 23657 14922 23723 14925
rect 19977 14920 23723 14922
rect 19977 14864 19982 14920
rect 20038 14864 22282 14920
rect 22338 14864 23662 14920
rect 23718 14864 23723 14920
rect 19977 14862 23723 14864
rect 19977 14859 20043 14862
rect 22277 14859 22343 14862
rect 23657 14859 23723 14862
rect 10501 14786 10567 14789
rect 9630 14784 10567 14786
rect 9630 14728 10506 14784
rect 10562 14728 10567 14784
rect 9630 14726 10567 14728
rect 10501 14723 10567 14726
rect 14365 14786 14431 14789
rect 18505 14786 18571 14789
rect 14365 14784 18571 14786
rect 14365 14728 14370 14784
rect 14426 14728 18510 14784
rect 18566 14728 18571 14784
rect 14365 14726 18571 14728
rect 14365 14723 14431 14726
rect 18505 14723 18571 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 14365 14652 14431 14653
rect 14365 14650 14412 14652
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 14320 14648 14412 14650
rect 14320 14592 14370 14648
rect 14320 14590 14412 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 14365 14588 14412 14590
rect 14476 14588 14482 14652
rect 14365 14587 14431 14588
rect 5349 14514 5415 14517
rect 8569 14514 8635 14517
rect 5349 14512 8635 14514
rect 5349 14456 5354 14512
rect 5410 14456 8574 14512
rect 8630 14456 8635 14512
rect 5349 14454 8635 14456
rect 5349 14451 5415 14454
rect 8569 14451 8635 14454
rect 12341 14378 12407 14381
rect 12893 14378 12959 14381
rect 19149 14378 19215 14381
rect 12341 14376 19215 14378
rect 12341 14320 12346 14376
rect 12402 14320 12898 14376
rect 12954 14320 19154 14376
rect 19210 14320 19215 14376
rect 12341 14318 19215 14320
rect 12341 14315 12407 14318
rect 12893 14315 12959 14318
rect 19149 14315 19215 14318
rect 22369 14378 22435 14381
rect 22737 14378 22803 14381
rect 23381 14378 23447 14381
rect 22369 14376 23447 14378
rect 22369 14320 22374 14376
rect 22430 14320 22742 14376
rect 22798 14320 23386 14376
rect 23442 14320 23447 14376
rect 22369 14318 23447 14320
rect 22369 14315 22435 14318
rect 22737 14315 22803 14318
rect 23381 14315 23447 14318
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 1761 13970 1827 13973
rect 19885 13970 19951 13973
rect 1761 13968 19951 13970
rect 1761 13912 1766 13968
rect 1822 13912 19890 13968
rect 19946 13912 19951 13968
rect 1761 13910 19951 13912
rect 1761 13907 1827 13910
rect 19885 13907 19951 13910
rect 0 13834 800 13864
rect 2037 13834 2103 13837
rect 0 13832 2103 13834
rect 0 13776 2042 13832
rect 2098 13776 2103 13832
rect 0 13774 2103 13776
rect 0 13744 800 13774
rect 2037 13771 2103 13774
rect 3509 13834 3575 13837
rect 3509 13832 3618 13834
rect 3509 13776 3514 13832
rect 3570 13776 3618 13832
rect 3509 13771 3618 13776
rect 5022 13772 5028 13836
rect 5092 13834 5098 13836
rect 6361 13834 6427 13837
rect 5092 13832 6427 13834
rect 5092 13776 6366 13832
rect 6422 13776 6427 13832
rect 5092 13774 6427 13776
rect 5092 13772 5098 13774
rect 6361 13771 6427 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 3558 13562 3618 13771
rect 4429 13696 4495 13701
rect 4429 13640 4434 13696
rect 4490 13640 4495 13696
rect 4429 13635 4495 13640
rect 7414 13636 7420 13700
rect 7484 13698 7490 13700
rect 11094 13698 11100 13700
rect 7484 13638 11100 13698
rect 7484 13636 7490 13638
rect 11094 13636 11100 13638
rect 11164 13636 11170 13700
rect 3693 13562 3759 13565
rect 3558 13560 3759 13562
rect 3558 13504 3698 13560
rect 3754 13504 3759 13560
rect 3558 13502 3759 13504
rect 4432 13562 4492 13635
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 4613 13562 4679 13565
rect 4432 13560 4679 13562
rect 4432 13504 4618 13560
rect 4674 13504 4679 13560
rect 4432 13502 4679 13504
rect 3693 13499 3759 13502
rect 4613 13499 4679 13502
rect 0 13426 800 13456
rect 1117 13426 1183 13429
rect 0 13424 1183 13426
rect 0 13368 1122 13424
rect 1178 13368 1183 13424
rect 0 13366 1183 13368
rect 0 13336 800 13366
rect 1117 13363 1183 13366
rect 1945 13426 2011 13429
rect 8334 13426 8340 13428
rect 1945 13424 8340 13426
rect 1945 13368 1950 13424
rect 2006 13368 8340 13424
rect 1945 13366 8340 13368
rect 1945 13363 2011 13366
rect 8334 13364 8340 13366
rect 8404 13364 8410 13428
rect 9397 13426 9463 13429
rect 31385 13426 31451 13429
rect 9397 13424 31451 13426
rect 9397 13368 9402 13424
rect 9458 13368 31390 13424
rect 31446 13368 31451 13424
rect 9397 13366 31451 13368
rect 9397 13363 9463 13366
rect 31385 13363 31451 13366
rect 1761 13290 1827 13293
rect 2037 13290 2103 13293
rect 18689 13290 18755 13293
rect 1761 13288 18755 13290
rect 1761 13232 1766 13288
rect 1822 13232 2042 13288
rect 2098 13232 18694 13288
rect 18750 13232 18755 13288
rect 1761 13230 18755 13232
rect 1761 13227 1827 13230
rect 2037 13227 2103 13230
rect 18689 13227 18755 13230
rect 4245 13154 4311 13157
rect 5574 13154 5580 13156
rect 4245 13152 5580 13154
rect 4245 13096 4250 13152
rect 4306 13096 5580 13152
rect 4245 13094 5580 13096
rect 4245 13091 4311 13094
rect 5574 13092 5580 13094
rect 5644 13092 5650 13156
rect 11278 13092 11284 13156
rect 11348 13154 11354 13156
rect 11881 13154 11947 13157
rect 11348 13152 11947 13154
rect 11348 13096 11886 13152
rect 11942 13096 11947 13152
rect 11348 13094 11947 13096
rect 11348 13092 11354 13094
rect 11881 13091 11947 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 7189 12882 7255 12885
rect 9581 12882 9647 12885
rect 7189 12880 9647 12882
rect 7189 12824 7194 12880
rect 7250 12824 9586 12880
rect 9642 12824 9647 12880
rect 7189 12822 9647 12824
rect 7189 12819 7255 12822
rect 9581 12819 9647 12822
rect 10685 12882 10751 12885
rect 22093 12882 22159 12885
rect 10685 12880 22159 12882
rect 10685 12824 10690 12880
rect 10746 12824 22098 12880
rect 22154 12824 22159 12880
rect 10685 12822 22159 12824
rect 10685 12819 10751 12822
rect 22093 12819 22159 12822
rect 4245 12746 4311 12749
rect 2730 12744 4311 12746
rect 2730 12688 4250 12744
rect 4306 12688 4311 12744
rect 2730 12686 4311 12688
rect 0 12610 800 12640
rect 2730 12610 2790 12686
rect 4245 12683 4311 12686
rect 7281 12746 7347 12749
rect 7598 12746 7604 12748
rect 7281 12744 7604 12746
rect 7281 12688 7286 12744
rect 7342 12688 7604 12744
rect 7281 12686 7604 12688
rect 7281 12683 7347 12686
rect 7598 12684 7604 12686
rect 7668 12684 7674 12748
rect 0 12550 2790 12610
rect 0 12520 800 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 6545 12474 6611 12477
rect 6862 12474 6868 12476
rect 6545 12472 6868 12474
rect 6545 12416 6550 12472
rect 6606 12416 6868 12472
rect 6545 12414 6868 12416
rect 6545 12411 6611 12414
rect 6862 12412 6868 12414
rect 6932 12412 6938 12476
rect 4889 12338 4955 12341
rect 10174 12338 10180 12340
rect 4889 12336 10180 12338
rect 4889 12280 4894 12336
rect 4950 12280 10180 12336
rect 4889 12278 10180 12280
rect 4889 12275 4955 12278
rect 10174 12276 10180 12278
rect 10244 12276 10250 12340
rect 17677 12338 17743 12341
rect 18413 12338 18479 12341
rect 17677 12336 18479 12338
rect 17677 12280 17682 12336
rect 17738 12280 18418 12336
rect 18474 12280 18479 12336
rect 17677 12278 18479 12280
rect 17677 12275 17743 12278
rect 18413 12275 18479 12278
rect 0 12202 800 12232
rect 1117 12202 1183 12205
rect 0 12200 1183 12202
rect 0 12144 1122 12200
rect 1178 12144 1183 12200
rect 0 12142 1183 12144
rect 0 12112 800 12142
rect 1117 12139 1183 12142
rect 7741 12202 7807 12205
rect 15745 12202 15811 12205
rect 7741 12200 15811 12202
rect 7741 12144 7746 12200
rect 7802 12144 15750 12200
rect 15806 12144 15811 12200
rect 7741 12142 15811 12144
rect 7741 12139 7807 12142
rect 15745 12139 15811 12142
rect 8518 12004 8524 12068
rect 8588 12066 8594 12068
rect 17401 12066 17467 12069
rect 8588 12064 17467 12066
rect 8588 12008 17406 12064
rect 17462 12008 17467 12064
rect 8588 12006 17467 12008
rect 8588 12004 8594 12006
rect 17401 12003 17467 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 3417 11930 3483 11933
rect 5073 11930 5139 11933
rect 3417 11928 5139 11930
rect 3417 11872 3422 11928
rect 3478 11872 5078 11928
rect 5134 11872 5139 11928
rect 3417 11870 5139 11872
rect 3417 11867 3483 11870
rect 5073 11867 5139 11870
rect 0 11794 800 11824
rect 1301 11794 1367 11797
rect 0 11792 1367 11794
rect 0 11736 1306 11792
rect 1362 11736 1367 11792
rect 0 11734 1367 11736
rect 0 11704 800 11734
rect 1301 11731 1367 11734
rect 9029 11658 9095 11661
rect 22686 11658 22692 11660
rect 9029 11656 22692 11658
rect 9029 11600 9034 11656
rect 9090 11600 22692 11656
rect 9029 11598 22692 11600
rect 9029 11595 9095 11598
rect 22686 11596 22692 11598
rect 22756 11596 22762 11660
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 5073 11386 5139 11389
rect 8845 11386 8911 11389
rect 5073 11384 8911 11386
rect 5073 11328 5078 11384
rect 5134 11328 8850 11384
rect 8906 11328 8911 11384
rect 5073 11326 8911 11328
rect 5073 11323 5139 11326
rect 8845 11323 8911 11326
rect 4153 11250 4219 11253
rect 4286 11250 4292 11252
rect 4153 11248 4292 11250
rect 4153 11192 4158 11248
rect 4214 11192 4292 11248
rect 4153 11190 4292 11192
rect 4153 11187 4219 11190
rect 4286 11188 4292 11190
rect 4356 11188 4362 11252
rect 7373 11250 7439 11253
rect 15878 11250 15884 11252
rect 7373 11248 15884 11250
rect 7373 11192 7378 11248
rect 7434 11192 15884 11248
rect 7373 11190 15884 11192
rect 7373 11187 7439 11190
rect 15878 11188 15884 11190
rect 15948 11188 15954 11252
rect 5165 11116 5231 11117
rect 5165 11114 5212 11116
rect 5120 11112 5212 11114
rect 5120 11056 5170 11112
rect 5120 11054 5212 11056
rect 5165 11052 5212 11054
rect 5276 11052 5282 11116
rect 8569 11114 8635 11117
rect 11513 11114 11579 11117
rect 8569 11112 11579 11114
rect 8569 11056 8574 11112
rect 8630 11056 11518 11112
rect 11574 11056 11579 11112
rect 8569 11054 11579 11056
rect 5165 11051 5231 11052
rect 8569 11051 8635 11054
rect 11513 11051 11579 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 6177 10842 6243 10845
rect 7230 10842 7236 10844
rect 6177 10840 7236 10842
rect 6177 10784 6182 10840
rect 6238 10784 7236 10840
rect 6177 10782 7236 10784
rect 6177 10779 6243 10782
rect 7230 10780 7236 10782
rect 7300 10780 7306 10844
rect 3233 10706 3299 10709
rect 3785 10706 3851 10709
rect 18781 10706 18847 10709
rect 3233 10704 18847 10706
rect 3233 10648 3238 10704
rect 3294 10648 3790 10704
rect 3846 10648 18786 10704
rect 18842 10648 18847 10704
rect 3233 10646 18847 10648
rect 3233 10643 3299 10646
rect 3785 10643 3851 10646
rect 18781 10643 18847 10646
rect 0 10570 800 10600
rect 3877 10570 3943 10573
rect 0 10568 3943 10570
rect 0 10512 3882 10568
rect 3938 10512 3943 10568
rect 0 10510 3943 10512
rect 0 10480 800 10510
rect 3877 10507 3943 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 2589 10162 2655 10165
rect 27705 10162 27771 10165
rect 0 10102 2284 10162
rect 0 10072 800 10102
rect 2224 10026 2284 10102
rect 2589 10160 27771 10162
rect 2589 10104 2594 10160
rect 2650 10104 27710 10160
rect 27766 10104 27771 10160
rect 2589 10102 27771 10104
rect 2589 10099 2655 10102
rect 27705 10099 27771 10102
rect 3601 10026 3667 10029
rect 2224 10024 3667 10026
rect 2224 9968 3606 10024
rect 3662 9968 3667 10024
rect 2224 9966 3667 9968
rect 3601 9963 3667 9966
rect 11053 10026 11119 10029
rect 11605 10026 11671 10029
rect 12750 10026 12756 10028
rect 11053 10024 12756 10026
rect 11053 9968 11058 10024
rect 11114 9968 11610 10024
rect 11666 9968 12756 10024
rect 11053 9966 12756 9968
rect 11053 9963 11119 9966
rect 11605 9963 11671 9966
rect 12750 9964 12756 9966
rect 12820 9964 12826 10028
rect 5758 9828 5764 9892
rect 5828 9890 5834 9892
rect 5901 9890 5967 9893
rect 5828 9888 5967 9890
rect 5828 9832 5906 9888
rect 5962 9832 5967 9888
rect 5828 9830 5967 9832
rect 5828 9828 5834 9830
rect 5901 9827 5967 9830
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 2865 9754 2931 9757
rect 0 9752 2931 9754
rect 0 9696 2870 9752
rect 2926 9696 2931 9752
rect 0 9694 2931 9696
rect 0 9664 800 9694
rect 2865 9691 2931 9694
rect 5809 9754 5875 9757
rect 6494 9754 6500 9756
rect 5809 9752 6500 9754
rect 5809 9696 5814 9752
rect 5870 9696 6500 9752
rect 5809 9694 6500 9696
rect 5809 9691 5875 9694
rect 6494 9692 6500 9694
rect 6564 9692 6570 9756
rect 5441 9620 5507 9621
rect 5390 9618 5396 9620
rect 5350 9558 5396 9618
rect 5460 9616 5507 9620
rect 5502 9560 5507 9616
rect 5390 9556 5396 9558
rect 5460 9556 5507 9560
rect 5441 9555 5507 9556
rect 3693 9482 3759 9485
rect 3693 9480 3986 9482
rect 3693 9424 3698 9480
rect 3754 9424 3986 9480
rect 3693 9422 3986 9424
rect 3693 9419 3759 9422
rect 0 9346 800 9376
rect 3926 9349 3986 9422
rect 0 9286 1594 9346
rect 3926 9344 4035 9349
rect 3926 9288 3974 9344
rect 4030 9288 4035 9344
rect 3926 9286 4035 9288
rect 0 9256 800 9286
rect 1534 9074 1594 9286
rect 3969 9283 4035 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 7189 9210 7255 9213
rect 7414 9210 7420 9212
rect 7189 9208 7420 9210
rect 7189 9152 7194 9208
rect 7250 9152 7420 9208
rect 7189 9150 7420 9152
rect 7189 9147 7255 9150
rect 7414 9148 7420 9150
rect 7484 9148 7490 9212
rect 7557 9210 7623 9213
rect 12801 9210 12867 9213
rect 7557 9208 12867 9210
rect 7557 9152 7562 9208
rect 7618 9152 12806 9208
rect 12862 9152 12867 9208
rect 7557 9150 12867 9152
rect 7557 9147 7623 9150
rect 12801 9147 12867 9150
rect 3417 9074 3483 9077
rect 1534 9072 3483 9074
rect 1534 9016 3422 9072
rect 3478 9016 3483 9072
rect 1534 9014 3483 9016
rect 3417 9011 3483 9014
rect 0 8938 800 8968
rect 4153 8938 4219 8941
rect 0 8936 4219 8938
rect 0 8880 4158 8936
rect 4214 8880 4219 8936
rect 0 8878 4219 8880
rect 0 8848 800 8878
rect 4153 8875 4219 8878
rect 3918 8740 3924 8804
rect 3988 8802 3994 8804
rect 4521 8802 4587 8805
rect 3988 8800 4587 8802
rect 3988 8744 4526 8800
rect 4582 8744 4587 8800
rect 3988 8742 4587 8744
rect 3988 8740 3994 8742
rect 4521 8739 4587 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 4245 8530 4311 8533
rect 0 8528 4311 8530
rect 0 8472 4250 8528
rect 4306 8472 4311 8528
rect 0 8470 4311 8472
rect 0 8440 800 8470
rect 4245 8467 4311 8470
rect 7925 8530 7991 8533
rect 11278 8530 11284 8532
rect 7925 8528 11284 8530
rect 7925 8472 7930 8528
rect 7986 8472 11284 8528
rect 7925 8470 11284 8472
rect 7925 8467 7991 8470
rect 11278 8468 11284 8470
rect 11348 8468 11354 8532
rect 12433 8530 12499 8533
rect 16573 8530 16639 8533
rect 12433 8528 16639 8530
rect 12433 8472 12438 8528
rect 12494 8472 16578 8528
rect 16634 8472 16639 8528
rect 12433 8470 16639 8472
rect 12433 8467 12499 8470
rect 16573 8467 16639 8470
rect 3693 8396 3759 8397
rect 3693 8394 3740 8396
rect 3648 8392 3740 8394
rect 3648 8336 3698 8392
rect 3648 8334 3740 8336
rect 3693 8332 3740 8334
rect 3804 8332 3810 8396
rect 9857 8394 9923 8397
rect 32622 8394 32628 8396
rect 9857 8392 32628 8394
rect 9857 8336 9862 8392
rect 9918 8336 32628 8392
rect 9857 8334 32628 8336
rect 3693 8331 3759 8332
rect 9857 8331 9923 8334
rect 32622 8332 32628 8334
rect 32692 8332 32698 8396
rect 6310 8196 6316 8260
rect 6380 8258 6386 8260
rect 6545 8258 6611 8261
rect 6380 8256 6611 8258
rect 6380 8200 6550 8256
rect 6606 8200 6611 8256
rect 6380 8198 6611 8200
rect 6380 8196 6386 8198
rect 6545 8195 6611 8198
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1301 8122 1367 8125
rect 0 8120 1367 8122
rect 0 8064 1306 8120
rect 1362 8064 1367 8120
rect 0 8062 1367 8064
rect 0 8032 800 8062
rect 1301 8059 1367 8062
rect 5574 8060 5580 8124
rect 5644 8122 5650 8124
rect 6361 8122 6427 8125
rect 5644 8120 6427 8122
rect 5644 8064 6366 8120
rect 6422 8064 6427 8120
rect 5644 8062 6427 8064
rect 5644 8060 5650 8062
rect 6361 8059 6427 8062
rect 5717 7986 5783 7989
rect 9806 7986 9812 7988
rect 5717 7984 9812 7986
rect 5717 7928 5722 7984
rect 5778 7928 9812 7984
rect 5717 7926 9812 7928
rect 5717 7923 5783 7926
rect 9806 7924 9812 7926
rect 9876 7924 9882 7988
rect 0 7714 800 7744
rect 3693 7714 3759 7717
rect 0 7712 3759 7714
rect 0 7656 3698 7712
rect 3754 7656 3759 7712
rect 0 7654 3759 7656
rect 0 7624 800 7654
rect 3693 7651 3759 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 3601 7442 3667 7445
rect 5022 7442 5028 7444
rect 3601 7440 5028 7442
rect 3601 7384 3606 7440
rect 3662 7384 5028 7440
rect 3601 7382 5028 7384
rect 3601 7379 3667 7382
rect 5022 7380 5028 7382
rect 5092 7380 5098 7444
rect 5349 7442 5415 7445
rect 22134 7442 22140 7444
rect 5349 7440 22140 7442
rect 5349 7384 5354 7440
rect 5410 7384 22140 7440
rect 5349 7382 22140 7384
rect 5349 7379 5415 7382
rect 22134 7380 22140 7382
rect 22204 7380 22210 7444
rect 0 7306 800 7336
rect 2773 7306 2839 7309
rect 0 7304 2839 7306
rect 0 7248 2778 7304
rect 2834 7248 2839 7304
rect 0 7246 2839 7248
rect 0 7216 800 7246
rect 2773 7243 2839 7246
rect 3969 7306 4035 7309
rect 13854 7306 13860 7308
rect 3969 7304 13860 7306
rect 3969 7248 3974 7304
rect 4030 7248 13860 7304
rect 3969 7246 13860 7248
rect 3969 7243 4035 7246
rect 13854 7244 13860 7246
rect 13924 7244 13930 7308
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6808 800 6838
rect 4061 6835 4127 6838
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1209 6490 1275 6493
rect 0 6488 1275 6490
rect 0 6432 1214 6488
rect 1270 6432 1275 6488
rect 0 6430 1275 6432
rect 0 6400 800 6430
rect 1209 6427 1275 6430
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 0 4450 800 4480
rect 4153 4450 4219 4453
rect 0 4448 4219 4450
rect 0 4392 4158 4448
rect 4214 4392 4219 4448
rect 0 4390 4219 4392
rect 0 4360 800 4390
rect 4153 4387 4219 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4042 800 4072
rect 4061 4042 4127 4045
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 0 3952 800 3982
rect 4061 3979 4127 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 2865 3634 2931 3637
rect 0 3632 2931 3634
rect 0 3576 2870 3632
rect 2926 3576 2931 3632
rect 0 3574 2931 3576
rect 0 3544 800 3574
rect 2865 3571 2931 3574
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 0 2410 800 2440
rect 1209 2410 1275 2413
rect 0 2408 1275 2410
rect 0 2352 1214 2408
rect 1270 2352 1275 2408
rect 0 2350 1275 2352
rect 0 2320 800 2350
rect 1209 2347 1275 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1301 2002 1367 2005
rect 0 2000 1367 2002
rect 0 1944 1306 2000
rect 1362 1944 1367 2000
rect 0 1942 1367 1944
rect 0 1912 800 1942
rect 1301 1939 1367 1942
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
<< via3 >>
rect 11652 24924 11716 24988
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 18460 24244 18524 24308
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 6500 23488 6564 23492
rect 6500 23432 6550 23488
rect 6550 23432 6564 23488
rect 6500 23428 6564 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 6316 23020 6380 23084
rect 22140 22944 22204 22948
rect 22140 22888 22190 22944
rect 22190 22888 22204 22944
rect 22140 22884 22204 22888
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 10180 22748 10244 22812
rect 5396 22612 5460 22676
rect 7236 22672 7300 22676
rect 7236 22616 7250 22672
rect 7250 22616 7300 22672
rect 7236 22612 7300 22616
rect 3924 22340 3988 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 22692 21796 22756 21860
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 4292 21388 4356 21452
rect 5212 21388 5276 21452
rect 5764 21252 5828 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 4292 21116 4356 21180
rect 6868 20768 6932 20772
rect 6868 20712 6918 20768
rect 6918 20712 6932 20768
rect 6868 20708 6932 20712
rect 11100 20708 11164 20772
rect 13860 20768 13924 20772
rect 13860 20712 13910 20768
rect 13910 20712 13924 20768
rect 13860 20708 13924 20712
rect 15884 20708 15948 20772
rect 17172 20708 17236 20772
rect 32076 20768 32140 20772
rect 32076 20712 32126 20768
rect 32126 20712 32140 20768
rect 32076 20708 32140 20712
rect 32628 20708 32692 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 7604 20088 7668 20092
rect 7604 20032 7618 20088
rect 7618 20032 7668 20088
rect 7604 20028 7668 20032
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7052 19620 7116 19684
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 8340 19212 8404 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 3740 18668 3804 18732
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 14412 18940 14476 19004
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 12756 18260 12820 18324
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 32076 18260 32140 18324
rect 5580 18048 5644 18052
rect 5580 17992 5630 18048
rect 5630 17992 5644 18048
rect 5580 17988 5644 17992
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7052 17716 7116 17780
rect 11652 17716 11716 17780
rect 12572 17716 12636 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 12388 17308 12452 17372
rect 9812 17096 9876 17100
rect 9812 17040 9862 17096
rect 9862 17040 9876 17096
rect 9812 17036 9876 17040
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 11652 16280 11716 16284
rect 11652 16224 11666 16280
rect 11666 16224 11716 16280
rect 11652 16220 11716 16224
rect 17172 16280 17236 16284
rect 17172 16224 17186 16280
rect 17186 16224 17236 16280
rect 17172 16220 17236 16224
rect 18460 16084 18524 16148
rect 8524 15948 8588 16012
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 14412 14648 14476 14652
rect 14412 14592 14426 14648
rect 14426 14592 14476 14648
rect 14412 14588 14476 14592
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 5028 13772 5092 13836
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 7420 13636 7484 13700
rect 11100 13636 11164 13700
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 8340 13364 8404 13428
rect 5580 13092 5644 13156
rect 11284 13092 11348 13156
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 7604 12684 7668 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 6868 12412 6932 12476
rect 10180 12276 10244 12340
rect 8524 12004 8588 12068
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 22692 11596 22756 11660
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 4292 11188 4356 11252
rect 15884 11188 15948 11252
rect 5212 11112 5276 11116
rect 5212 11056 5226 11112
rect 5226 11056 5276 11112
rect 5212 11052 5276 11056
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 7236 10780 7300 10844
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 12756 9964 12820 10028
rect 5764 9828 5828 9892
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 6500 9692 6564 9756
rect 5396 9616 5460 9620
rect 5396 9560 5446 9616
rect 5446 9560 5460 9616
rect 5396 9556 5460 9560
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7420 9148 7484 9212
rect 3924 8740 3988 8804
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 11284 8468 11348 8532
rect 3740 8392 3804 8396
rect 3740 8336 3754 8392
rect 3754 8336 3804 8392
rect 3740 8332 3804 8336
rect 32628 8332 32692 8396
rect 6316 8196 6380 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 5580 8060 5644 8124
rect 9812 7924 9876 7988
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 5028 7380 5092 7444
rect 22140 7380 22204 7444
rect 13860 7244 13924 7308
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 11651 24988 11717 24989
rect 11651 24924 11652 24988
rect 11716 24924 11717 24988
rect 11651 24923 11717 24924
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 6499 23492 6565 23493
rect 6499 23428 6500 23492
rect 6564 23428 6565 23492
rect 6499 23427 6565 23428
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 6315 23084 6381 23085
rect 6315 23020 6316 23084
rect 6380 23020 6381 23084
rect 6315 23019 6381 23020
rect 5395 22676 5461 22677
rect 5395 22612 5396 22676
rect 5460 22612 5461 22676
rect 5395 22611 5461 22612
rect 3923 22404 3989 22405
rect 3923 22340 3924 22404
rect 3988 22340 3989 22404
rect 3923 22339 3989 22340
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 3739 18732 3805 18733
rect 3739 18668 3740 18732
rect 3804 18668 3805 18732
rect 3739 18667 3805 18668
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 3742 8397 3802 18667
rect 3926 8805 3986 22339
rect 4291 21452 4357 21453
rect 4291 21388 4292 21452
rect 4356 21388 4357 21452
rect 4291 21387 4357 21388
rect 5211 21452 5277 21453
rect 5211 21388 5212 21452
rect 5276 21388 5277 21452
rect 5211 21387 5277 21388
rect 4294 21181 4354 21387
rect 4291 21180 4357 21181
rect 4291 21116 4292 21180
rect 4356 21116 4357 21180
rect 4291 21115 4357 21116
rect 4294 11253 4354 21115
rect 5027 13836 5093 13837
rect 5027 13772 5028 13836
rect 5092 13772 5093 13836
rect 5027 13771 5093 13772
rect 4291 11252 4357 11253
rect 4291 11188 4292 11252
rect 4356 11188 4357 11252
rect 4291 11187 4357 11188
rect 3923 8804 3989 8805
rect 3923 8740 3924 8804
rect 3988 8740 3989 8804
rect 3923 8739 3989 8740
rect 3739 8396 3805 8397
rect 3739 8332 3740 8396
rect 3804 8332 3805 8396
rect 3739 8331 3805 8332
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 5030 7445 5090 13771
rect 5214 11117 5274 21387
rect 5211 11116 5277 11117
rect 5211 11052 5212 11116
rect 5276 11052 5277 11116
rect 5211 11051 5277 11052
rect 5398 9621 5458 22611
rect 5763 21316 5829 21317
rect 5763 21252 5764 21316
rect 5828 21252 5829 21316
rect 5763 21251 5829 21252
rect 5579 18052 5645 18053
rect 5579 17988 5580 18052
rect 5644 17988 5645 18052
rect 5579 17987 5645 17988
rect 5582 13157 5642 17987
rect 5579 13156 5645 13157
rect 5579 13092 5580 13156
rect 5644 13092 5645 13156
rect 5579 13091 5645 13092
rect 5395 9620 5461 9621
rect 5395 9556 5396 9620
rect 5460 9556 5461 9620
rect 5395 9555 5461 9556
rect 5582 8125 5642 13091
rect 5766 9893 5826 21251
rect 5763 9892 5829 9893
rect 5763 9828 5764 9892
rect 5828 9828 5829 9892
rect 5763 9827 5829 9828
rect 6318 8261 6378 23019
rect 6502 9757 6562 23427
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7235 22676 7301 22677
rect 7235 22612 7236 22676
rect 7300 22612 7301 22676
rect 7235 22611 7301 22612
rect 6867 20772 6933 20773
rect 6867 20708 6868 20772
rect 6932 20708 6933 20772
rect 6867 20707 6933 20708
rect 6870 12477 6930 20707
rect 7051 19684 7117 19685
rect 7051 19620 7052 19684
rect 7116 19620 7117 19684
rect 7051 19619 7117 19620
rect 7054 17781 7114 19619
rect 7051 17780 7117 17781
rect 7051 17716 7052 17780
rect 7116 17716 7117 17780
rect 7051 17715 7117 17716
rect 6867 12476 6933 12477
rect 6867 12412 6868 12476
rect 6932 12412 6933 12476
rect 6867 12411 6933 12412
rect 7238 10845 7298 22611
rect 7944 21792 8264 22816
rect 10179 22812 10245 22813
rect 10179 22748 10180 22812
rect 10244 22748 10245 22812
rect 10179 22747 10245 22748
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7603 20092 7669 20093
rect 7603 20028 7604 20092
rect 7668 20028 7669 20092
rect 7603 20027 7669 20028
rect 7419 13700 7485 13701
rect 7419 13636 7420 13700
rect 7484 13636 7485 13700
rect 7419 13635 7485 13636
rect 7235 10844 7301 10845
rect 7235 10780 7236 10844
rect 7300 10780 7301 10844
rect 7235 10779 7301 10780
rect 6499 9756 6565 9757
rect 6499 9692 6500 9756
rect 6564 9692 6565 9756
rect 6499 9691 6565 9692
rect 7422 9213 7482 13635
rect 7606 12749 7666 20027
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 8339 19276 8405 19277
rect 8339 19212 8340 19276
rect 8404 19212 8405 19276
rect 8339 19211 8405 19212
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 8342 13429 8402 19211
rect 9811 17100 9877 17101
rect 9811 17036 9812 17100
rect 9876 17036 9877 17100
rect 9811 17035 9877 17036
rect 8523 16012 8589 16013
rect 8523 15948 8524 16012
rect 8588 15948 8589 16012
rect 8523 15947 8589 15948
rect 8339 13428 8405 13429
rect 8339 13364 8340 13428
rect 8404 13364 8405 13428
rect 8339 13363 8405 13364
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7603 12748 7669 12749
rect 7603 12684 7604 12748
rect 7668 12684 7669 12748
rect 7603 12683 7669 12684
rect 7944 12000 8264 13024
rect 8526 12069 8586 15947
rect 8523 12068 8589 12069
rect 8523 12004 8524 12068
rect 8588 12004 8589 12068
rect 8523 12003 8589 12004
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7419 9212 7485 9213
rect 7419 9148 7420 9212
rect 7484 9148 7485 9212
rect 7419 9147 7485 9148
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 6315 8260 6381 8261
rect 6315 8196 6316 8260
rect 6380 8196 6381 8260
rect 6315 8195 6381 8196
rect 5579 8124 5645 8125
rect 5579 8060 5580 8124
rect 5644 8060 5645 8124
rect 5579 8059 5645 8060
rect 7944 7648 8264 8672
rect 9814 7989 9874 17035
rect 10182 12341 10242 22747
rect 11099 20772 11165 20773
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 11102 13701 11162 20707
rect 11654 17781 11714 24923
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 17944 23968 18264 24528
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 18459 24308 18525 24309
rect 18459 24244 18460 24308
rect 18524 24244 18525 24308
rect 18459 24243 18525 24244
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 13859 20772 13925 20773
rect 13859 20708 13860 20772
rect 13924 20708 13925 20772
rect 13859 20707 13925 20708
rect 15883 20772 15949 20773
rect 15883 20708 15884 20772
rect 15948 20708 15949 20772
rect 15883 20707 15949 20708
rect 17171 20772 17237 20773
rect 17171 20708 17172 20772
rect 17236 20708 17237 20772
rect 17171 20707 17237 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12755 18324 12821 18325
rect 12755 18260 12756 18324
rect 12820 18260 12821 18324
rect 12755 18259 12821 18260
rect 11651 17780 11717 17781
rect 11651 17716 11652 17780
rect 11716 17716 11717 17780
rect 11651 17715 11717 17716
rect 12571 17780 12637 17781
rect 12571 17716 12572 17780
rect 12636 17716 12637 17780
rect 12571 17715 12637 17716
rect 11654 16285 11714 17715
rect 12387 17372 12453 17373
rect 12387 17308 12388 17372
rect 12452 17370 12453 17372
rect 12574 17370 12634 17715
rect 12452 17310 12634 17370
rect 12452 17308 12453 17310
rect 12387 17307 12453 17308
rect 11651 16284 11717 16285
rect 11651 16220 11652 16284
rect 11716 16220 11717 16284
rect 11651 16219 11717 16220
rect 11099 13700 11165 13701
rect 11099 13636 11100 13700
rect 11164 13636 11165 13700
rect 11099 13635 11165 13636
rect 11283 13156 11349 13157
rect 11283 13092 11284 13156
rect 11348 13092 11349 13156
rect 11283 13091 11349 13092
rect 10179 12340 10245 12341
rect 10179 12276 10180 12340
rect 10244 12276 10245 12340
rect 10179 12275 10245 12276
rect 11286 8533 11346 13091
rect 12758 10029 12818 18259
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12755 10028 12821 10029
rect 12755 9964 12756 10028
rect 12820 9964 12821 10028
rect 12755 9963 12821 9964
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 11283 8532 11349 8533
rect 11283 8468 11284 8532
rect 11348 8468 11349 8532
rect 11283 8467 11349 8468
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 9811 7988 9877 7989
rect 9811 7924 9812 7988
rect 9876 7924 9877 7988
rect 9811 7923 9877 7924
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 5027 7444 5093 7445
rect 5027 7380 5028 7444
rect 5092 7380 5093 7444
rect 5027 7379 5093 7380
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 7104 13264 8128
rect 13862 7309 13922 20707
rect 14411 19004 14477 19005
rect 14411 18940 14412 19004
rect 14476 18940 14477 19004
rect 14411 18939 14477 18940
rect 14414 14653 14474 18939
rect 14411 14652 14477 14653
rect 14411 14588 14412 14652
rect 14476 14588 14477 14652
rect 14411 14587 14477 14588
rect 15886 11253 15946 20707
rect 17174 16285 17234 20707
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17171 16284 17237 16285
rect 17171 16220 17172 16284
rect 17236 16220 17237 16284
rect 17171 16219 17237 16220
rect 17944 15264 18264 16288
rect 18462 16149 18522 24243
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22139 22948 22205 22949
rect 22139 22884 22140 22948
rect 22204 22884 22205 22948
rect 22139 22883 22205 22884
rect 18459 16148 18525 16149
rect 18459 16084 18460 16148
rect 18524 16084 18525 16148
rect 18459 16083 18525 16084
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 15883 11252 15949 11253
rect 15883 11188 15884 11252
rect 15948 11188 15949 11252
rect 15883 11187 15949 11188
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 13859 7308 13925 7309
rect 13859 7244 13860 7308
rect 13924 7244 13925 7308
rect 13859 7243 13925 7244
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 6560 18264 7584
rect 22142 7445 22202 22883
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22691 21860 22757 21861
rect 22691 21796 22692 21860
rect 22756 21796 22757 21860
rect 22691 21795 22757 21796
rect 22694 11661 22754 21795
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22691 11660 22757 11661
rect 22691 11596 22692 11660
rect 22756 11596 22757 11660
rect 22691 11595 22757 11596
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22139 7444 22205 7445
rect 22139 7380 22140 7444
rect 22204 7380 22205 7444
rect 22139 7379 22205 7380
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32075 20772 32141 20773
rect 32075 20708 32076 20772
rect 32140 20708 32141 20772
rect 32075 20707 32141 20708
rect 32627 20772 32693 20773
rect 32627 20708 32628 20772
rect 32692 20708 32693 20772
rect 32627 20707 32693 20708
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 32078 18325 32138 20707
rect 32075 18324 32141 18325
rect 32075 18260 32076 18324
rect 32140 18260 32141 18324
rect 32075 18259 32141 18260
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 32630 8397 32690 20707
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32627 8396 32693 8397
rect 32627 8332 32628 8396
rect 32692 8332 32693 8396
rect 32627 8331 32693 8332
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22448 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1679235063
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1679235063
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1679235063
transform 1 0 10672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1679235063
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1679235063
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1679235063
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 4140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1679235063
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1679235063
transform 1 0 3956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1679235063
transform 1 0 6072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1679235063
transform 1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2208 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1679235063
transform 1 0 2116 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1679235063
transform 1 0 4232 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1679235063
transform 1 0 20884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1679235063
transform 1 0 2576 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _132_
timestamp 1679235063
transform 1 0 8372 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1679235063
transform 1 0 2116 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _134_
timestamp 1679235063
transform 1 0 5888 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _135_
timestamp 1679235063
transform 1 0 3404 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1679235063
transform 1 0 4232 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _137_
timestamp 1679235063
transform 1 0 2576 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 35512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 36248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 33856 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 32292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 33028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 31280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 34868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 33856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _147_
timestamp 1679235063
transform 1 0 29716 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _149_
timestamp 1679235063
transform 1 0 28244 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1679235063
transform 1 0 18584 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _151_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1679235063
transform 1 0 34224 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1679235063
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1679235063
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1679235063
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1679235063
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1679235063
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 4416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 3956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 6532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 33396 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 13616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 13800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1679235063
transform 1 0 15180 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1679235063
transform 1 0 15364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1679235063
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1679235063
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1679235063
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1679235063
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1679235063
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1679235063
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1679235063
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1679235063
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1679235063
transform 1 0 3864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1679235063
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1679235063
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1679235063
transform 1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 5612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1679235063
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1679235063
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1679235063
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1679235063
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1679235063
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1679235063
transform 1 0 1564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1679235063
transform 1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1679235063
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1679235063
transform 1 0 32476 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 34408 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 34776 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1679235063
transform 1 0 34040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 22448 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform 1 0 30360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1679235063
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1679235063
transform 1 0 16376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 11132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 9016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 9016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 6440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 21620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 23644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
timestamp 1679235063
transform 1 0 22816 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1679235063
transform 1 0 28520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 28336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
timestamp 1679235063
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 32016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 19320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 14996 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 19320 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 26496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold7_A
timestamp 1679235063
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1679235063
transform 1 0 27876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold14_A
timestamp 1679235063
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold16_A
timestamp 1679235063
transform 1 0 25208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold18_A
timestamp 1679235063
transform 1 0 30544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold20_A
timestamp 1679235063
transform 1 0 33580 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold21_A
timestamp 1679235063
transform 1 0 32844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold22_A
timestamp 1679235063
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold23_A
timestamp 1679235063
transform 1 0 38088 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold24_A
timestamp 1679235063
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold25_A
timestamp 1679235063
transform 1 0 34224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold26_A
timestamp 1679235063
transform 1 0 36800 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold27_A
timestamp 1679235063
transform 1 0 42044 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold28_A
timestamp 1679235063
transform 1 0 37904 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold29_A
timestamp 1679235063
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold30_A
timestamp 1679235063
transform 1 0 40848 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold31_A
timestamp 1679235063
transform 1 0 41032 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold32_A
timestamp 1679235063
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold33_A
timestamp 1679235063
transform 1 0 33764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold34_A
timestamp 1679235063
transform 1 0 36892 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold35_A
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold36_A
timestamp 1679235063
transform 1 0 47380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold39_A
timestamp 1679235063
transform 1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 4416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 4140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 5428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 5060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 3312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 4416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 5244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 34592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 35420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 37904 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 39376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 31832 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 39192 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 37904 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 41768 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 6532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 32660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 33580 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 34316 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 46276 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 47564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 44620 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 46092 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1679235063
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1679235063
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform 1 0 47932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform 1 0 47748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1679235063
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1679235063
transform 1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1679235063
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1679235063
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1679235063
transform 1 0 1656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1679235063
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1679235063
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1679235063
transform 1 0 19872 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1679235063
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1679235063
transform 1 0 27416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1679235063
transform 1 0 10856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 1679235063
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output142_A
timestamp 1679235063
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20884 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14904 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 21896 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 27232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 27876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 29992 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 30176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 31740 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 33396 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 29808 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 32016 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 36064 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 31556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 32200 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 29716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 30912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 37444 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 21620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20056 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 4140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31740 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 28796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 12328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22264 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23920 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 32384 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 32568 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28152 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_19.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 32292 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_49.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 31464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 30728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 30544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 25576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 26128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 25668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 25944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21528 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22724 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 30176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 32936 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 31096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14996 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 1472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 33488 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 33120 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22448 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8096 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 4140 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4140 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 5336 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 5428 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 7360 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8004 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8464 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10028 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 11224 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 11960 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9200 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9568 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 4232 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 6808 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191
timestamp 1679235063
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 4048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10580 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 3956 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14260 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 8096 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 9384 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10856 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14352 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193
timestamp 1679235063
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 6716 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 28612 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8740 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 26956 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 20884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 25760 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 22908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22172 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 24656 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27508 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29716 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17112 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9568 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 14720 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 14904 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 8464 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 13616 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 12788 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 19504 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 18952 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 23092 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 19596 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 24932 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 25300 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22
timestamp 1679235063
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1679235063
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1679235063
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1679235063
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1679235063
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1679235063
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1679235063
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1679235063
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1679235063
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1679235063
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1679235063
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_264
timestamp 1679235063
transform 1 0 25392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1679235063
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1679235063
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_289
timestamp 1679235063
transform 1 0 27692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_293
timestamp 1679235063
transform 1 0 28060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_303
timestamp 1679235063
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1679235063
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_309
timestamp 1679235063
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_317
timestamp 1679235063
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_322
timestamp 1679235063
transform 1 0 30728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1679235063
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1679235063
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1679235063
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1679235063
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1679235063
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1679235063
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_395
timestamp 1679235063
transform 1 0 37444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_407
timestamp 1679235063
transform 1 0 38548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1679235063
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1679235063
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1679235063
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1679235063
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1679235063
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1679235063
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1679235063
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1679235063
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1679235063
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1679235063
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1679235063
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1679235063
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1679235063
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1679235063
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1679235063
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1679235063
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_67
timestamp 1679235063
transform 1 0 7268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1679235063
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1679235063
transform 1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1679235063
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1679235063
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1679235063
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1679235063
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1679235063
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_142
timestamp 1679235063
transform 1 0 14168 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1679235063
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1679235063
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1679235063
transform 1 0 17112 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp 1679235063
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_188
timestamp 1679235063
transform 1 0 18400 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1679235063
transform 1 0 19504 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1679235063
transform 1 0 20240 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1679235063
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1679235063
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1679235063
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_261
timestamp 1679235063
transform 1 0 25116 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_268
timestamp 1679235063
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1679235063
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_293
timestamp 1679235063
transform 1 0 28060 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_297
timestamp 1679235063
transform 1 0 28428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_309
timestamp 1679235063
transform 1 0 29532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_321
timestamp 1679235063
transform 1 0 30636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1679235063
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1679235063
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1679235063
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_349
timestamp 1679235063
transform 1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_355
timestamp 1679235063
transform 1 0 33764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1679235063
transform 1 0 34868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1679235063
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1679235063
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1679235063
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_411
timestamp 1679235063
transform 1 0 38916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_423
timestamp 1679235063
transform 1 0 40020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_435
timestamp 1679235063
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1679235063
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1679235063
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1679235063
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1679235063
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1679235063
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1679235063
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1679235063
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1679235063
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1679235063
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1679235063
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1679235063
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1679235063
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_34
timestamp 1679235063
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_40
timestamp 1679235063
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_52
timestamp 1679235063
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1679235063
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1679235063
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1679235063
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_120
timestamp 1679235063
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1679235063
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1679235063
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1679235063
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1679235063
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1679235063
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1679235063
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1679235063
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1679235063
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1679235063
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1679235063
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1679235063
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1679235063
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1679235063
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1679235063
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1679235063
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1679235063
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1679235063
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1679235063
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1679235063
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1679235063
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_365
timestamp 1679235063
transform 1 0 34684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_373
timestamp 1679235063
transform 1 0 35420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_392
timestamp 1679235063
transform 1 0 37168 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_398
timestamp 1679235063
transform 1 0 37720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1679235063
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1679235063
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1679235063
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1679235063
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1679235063
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1679235063
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1679235063
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1679235063
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1679235063
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1679235063
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1679235063
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1679235063
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1679235063
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_5
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1679235063
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1679235063
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1679235063
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1679235063
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1679235063
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1679235063
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1679235063
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1679235063
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1679235063
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1679235063
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1679235063
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1679235063
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1679235063
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1679235063
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1679235063
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1679235063
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1679235063
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1679235063
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1679235063
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1679235063
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1679235063
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1679235063
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1679235063
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1679235063
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1679235063
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1679235063
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1679235063
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1679235063
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1679235063
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1679235063
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1679235063
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1679235063
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1679235063
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1679235063
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1679235063
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1679235063
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1679235063
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1679235063
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1679235063
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1679235063
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1679235063
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1679235063
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1679235063
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1679235063
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1679235063
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1679235063
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1679235063
transform 1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1679235063
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1679235063
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1679235063
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1679235063
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1679235063
transform 1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1679235063
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1679235063
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1679235063
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1679235063
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1679235063
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1679235063
transform 1 0 24840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1679235063
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_281
timestamp 1679235063
transform 1 0 26956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_293
timestamp 1679235063
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1679235063
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1679235063
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1679235063
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1679235063
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1679235063
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1679235063
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1679235063
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1679235063
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1679235063
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1679235063
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1679235063
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1679235063
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1679235063
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1679235063
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1679235063
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1679235063
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1679235063
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1679235063
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1679235063
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1679235063
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1679235063
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1679235063
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1679235063
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1679235063
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_25
timestamp 1679235063
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_37
timestamp 1679235063
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1679235063
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1679235063
transform 1 0 15548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1679235063
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp 1679235063
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1679235063
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1679235063
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1679235063
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1679235063
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_238
timestamp 1679235063
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1679235063
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1679235063
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1679235063
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1679235063
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1679235063
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_312
timestamp 1679235063
transform 1 0 29808 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_324
timestamp 1679235063
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1679235063
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1679235063
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1679235063
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1679235063
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1679235063
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1679235063
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1679235063
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1679235063
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1679235063
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1679235063
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1679235063
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1679235063
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1679235063
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1679235063
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1679235063
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1679235063
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1679235063
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1679235063
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1679235063
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1679235063
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1679235063
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_22
timestamp 1679235063
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1679235063
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_199
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_211
timestamp 1679235063
transform 1 0 20516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1679235063
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_225
timestamp 1679235063
transform 1 0 21804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_237
timestamp 1679235063
transform 1 0 22908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1679235063
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_269
timestamp 1679235063
transform 1 0 25852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1679235063
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1679235063
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1679235063
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1679235063
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1679235063
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1679235063
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1679235063
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1679235063
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1679235063
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1679235063
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1679235063
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1679235063
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1679235063
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1679235063
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1679235063
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1679235063
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1679235063
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1679235063
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1679235063
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1679235063
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1679235063
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1679235063
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1679235063
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1679235063
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1679235063
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_22
timestamp 1679235063
transform 1 0 3128 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_29
timestamp 1679235063
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1679235063
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1679235063
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1679235063
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1679235063
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1679235063
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1679235063
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp 1679235063
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_238
timestamp 1679235063
transform 1 0 23000 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_250
timestamp 1679235063
transform 1 0 24104 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_262
timestamp 1679235063
transform 1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1679235063
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1679235063
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1679235063
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1679235063
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1679235063
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1679235063
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1679235063
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1679235063
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1679235063
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1679235063
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1679235063
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1679235063
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1679235063
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1679235063
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1679235063
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1679235063
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1679235063
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1679235063
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1679235063
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1679235063
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1679235063
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1679235063
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1679235063
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1679235063
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1679235063
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1679235063
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1679235063
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1679235063
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1679235063
transform 1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1679235063
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1679235063
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1679235063
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_34
timestamp 1679235063
transform 1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_42
timestamp 1679235063
transform 1 0 4968 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_54
timestamp 1679235063
transform 1 0 6072 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_66
timestamp 1679235063
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1679235063
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_106
timestamp 1679235063
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1679235063
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1679235063
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1679235063
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1679235063
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1679235063
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1679235063
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1679235063
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_243
timestamp 1679235063
transform 1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1679235063
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1679235063
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1679235063
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1679235063
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1679235063
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1679235063
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1679235063
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1679235063
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1679235063
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1679235063
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1679235063
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1679235063
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1679235063
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1679235063
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1679235063
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1679235063
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1679235063
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1679235063
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1679235063
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1679235063
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1679235063
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1679235063
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1679235063
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1679235063
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1679235063
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1679235063
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1679235063
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1679235063
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1679235063
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1679235063
transform 1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_28
timestamp 1679235063
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_34
timestamp 1679235063
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_41
timestamp 1679235063
transform 1 0 4876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1679235063
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1679235063
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1679235063
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1679235063
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_120
timestamp 1679235063
transform 1 0 12144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_127
timestamp 1679235063
transform 1 0 12788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_133
timestamp 1679235063
transform 1 0 13340 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_144
timestamp 1679235063
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 1679235063
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1679235063
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1679235063
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1679235063
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1679235063
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1679235063
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1679235063
transform 1 0 24012 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1679235063
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1679235063
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1679235063
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1679235063
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1679235063
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1679235063
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1679235063
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1679235063
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1679235063
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1679235063
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1679235063
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1679235063
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1679235063
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1679235063
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1679235063
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1679235063
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1679235063
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1679235063
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1679235063
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1679235063
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1679235063
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1679235063
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1679235063
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1679235063
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1679235063
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1679235063
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1679235063
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1679235063
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1679235063
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1679235063
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1679235063
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1679235063
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_51
timestamp 1679235063
transform 1 0 5796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_61
timestamp 1679235063
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_66
timestamp 1679235063
transform 1 0 7176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_75
timestamp 1679235063
transform 1 0 8004 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_81
timestamp 1679235063
transform 1 0 8556 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1679235063
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_101
timestamp 1679235063
transform 1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_120
timestamp 1679235063
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1679235063
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_128
timestamp 1679235063
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1679235063
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_143
timestamp 1679235063
transform 1 0 14260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1679235063
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_161
timestamp 1679235063
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_173
timestamp 1679235063
transform 1 0 17020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1679235063
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1679235063
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1679235063
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1679235063
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1679235063
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1679235063
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1679235063
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1679235063
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1679235063
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1679235063
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1679235063
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1679235063
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1679235063
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1679235063
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1679235063
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1679235063
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1679235063
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1679235063
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1679235063
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1679235063
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1679235063
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1679235063
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1679235063
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1679235063
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1679235063
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1679235063
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1679235063
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1679235063
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1679235063
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1679235063
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1679235063
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1679235063
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1679235063
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1679235063
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1679235063
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1679235063
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_33
timestamp 1679235063
transform 1 0 4140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1679235063
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1679235063
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_45
timestamp 1679235063
transform 1 0 5244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_48
timestamp 1679235063
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1679235063
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_59
timestamp 1679235063
transform 1 0 6532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1679235063
transform 1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1679235063
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1679235063
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1679235063
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_107
timestamp 1679235063
transform 1 0 10948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1679235063
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1679235063
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_129
timestamp 1679235063
transform 1 0 12972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1679235063
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1679235063
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1679235063
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1679235063
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1679235063
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1679235063
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1679235063
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1679235063
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1679235063
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1679235063
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1679235063
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1679235063
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1679235063
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1679235063
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1679235063
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1679235063
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1679235063
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1679235063
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1679235063
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1679235063
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1679235063
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1679235063
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1679235063
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1679235063
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1679235063
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1679235063
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1679235063
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1679235063
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1679235063
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1679235063
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1679235063
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1679235063
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1679235063
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1679235063
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1679235063
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1679235063
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1679235063
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1679235063
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1679235063
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1679235063
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1679235063
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_8
timestamp 1679235063
transform 1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1679235063
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_34
timestamp 1679235063
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1679235063
transform 1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1679235063
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1679235063
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1679235063
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1679235063
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1679235063
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1679235063
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1679235063
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1679235063
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1679235063
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_152
timestamp 1679235063
transform 1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1679235063
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1679235063
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1679235063
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1679235063
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1679235063
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_193
timestamp 1679235063
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1679235063
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1679235063
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1679235063
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1679235063
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1679235063
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1679235063
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1679235063
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1679235063
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1679235063
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1679235063
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1679235063
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1679235063
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1679235063
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1679235063
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1679235063
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1679235063
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1679235063
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1679235063
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1679235063
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1679235063
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1679235063
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1679235063
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1679235063
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1679235063
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1679235063
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1679235063
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1679235063
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1679235063
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1679235063
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1679235063
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1679235063
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1679235063
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1679235063
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_21
timestamp 1679235063
transform 1 0 3036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1679235063
transform 1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1679235063
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_44
timestamp 1679235063
transform 1 0 5152 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1679235063
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1679235063
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_59
timestamp 1679235063
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1679235063
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1679235063
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1679235063
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1679235063
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1679235063
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1679235063
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1679235063
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1679235063
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1679235063
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1679235063
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1679235063
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1679235063
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1679235063
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1679235063
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1679235063
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1679235063
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_294
timestamp 1679235063
transform 1 0 28152 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_300
timestamp 1679235063
transform 1 0 28704 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_312
timestamp 1679235063
transform 1 0 29808 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_324
timestamp 1679235063
transform 1 0 30912 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1679235063
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1679235063
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1679235063
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1679235063
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1679235063
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1679235063
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1679235063
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1679235063
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1679235063
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1679235063
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1679235063
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1679235063
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1679235063
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1679235063
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1679235063
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1679235063
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1679235063
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1679235063
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1679235063
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1679235063
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1679235063
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1679235063
transform 1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1679235063
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1679235063
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_31
timestamp 1679235063
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1679235063
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_48
timestamp 1679235063
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_54
timestamp 1679235063
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1679235063
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1679235063
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1679235063
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1679235063
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1679235063
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1679235063
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1679235063
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_143
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1679235063
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1679235063
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_219
timestamp 1679235063
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_225
timestamp 1679235063
transform 1 0 21804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_237
timestamp 1679235063
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1679235063
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1679235063
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1679235063
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1679235063
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1679235063
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1679235063
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1679235063
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1679235063
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1679235063
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1679235063
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1679235063
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1679235063
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1679235063
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1679235063
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1679235063
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1679235063
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1679235063
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1679235063
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1679235063
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1679235063
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1679235063
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1679235063
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1679235063
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1679235063
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1679235063
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1679235063
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1679235063
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1679235063
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1679235063
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1679235063
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_35
timestamp 1679235063
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1679235063
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1679235063
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1679235063
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1679235063
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1679235063
transform 1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1679235063
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1679235063
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_116
timestamp 1679235063
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1679235063
transform 1 0 13892 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1679235063
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1679235063
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1679235063
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_229
timestamp 1679235063
transform 1 0 22172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_241
timestamp 1679235063
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_253
timestamp 1679235063
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_265
timestamp 1679235063
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1679235063
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1679235063
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1679235063
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1679235063
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1679235063
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1679235063
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1679235063
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1679235063
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1679235063
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1679235063
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1679235063
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1679235063
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1679235063
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1679235063
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1679235063
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1679235063
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1679235063
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1679235063
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1679235063
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1679235063
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1679235063
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1679235063
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1679235063
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1679235063
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1679235063
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1679235063
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1679235063
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1679235063
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1679235063
transform 1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1679235063
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1679235063
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_31
timestamp 1679235063
transform 1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_36
timestamp 1679235063
transform 1 0 4416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1679235063
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1679235063
transform 1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1679235063
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1679235063
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1679235063
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1679235063
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1679235063
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_145
timestamp 1679235063
transform 1 0 14444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1679235063
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_172
timestamp 1679235063
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1679235063
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_235
timestamp 1679235063
transform 1 0 22724 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_239
timestamp 1679235063
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1679235063
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1679235063
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1679235063
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1679235063
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1679235063
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1679235063
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1679235063
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_334
timestamp 1679235063
transform 1 0 31832 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1679235063
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1679235063
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1679235063
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1679235063
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1679235063
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1679235063
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1679235063
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1679235063
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1679235063
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1679235063
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1679235063
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1679235063
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1679235063
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1679235063
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1679235063
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1679235063
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1679235063
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1679235063
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1679235063
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1679235063
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1679235063
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_25
timestamp 1679235063
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1679235063
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1679235063
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1679235063
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1679235063
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1679235063
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1679235063
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1679235063
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1679235063
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1679235063
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1679235063
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1679235063
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1679235063
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1679235063
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_228
timestamp 1679235063
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_251
timestamp 1679235063
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_255
timestamp 1679235063
transform 1 0 24564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_267
timestamp 1679235063
transform 1 0 25668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1679235063
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1679235063
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1679235063
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1679235063
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1679235063
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1679235063
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1679235063
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1679235063
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1679235063
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1679235063
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1679235063
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1679235063
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1679235063
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1679235063
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1679235063
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1679235063
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1679235063
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1679235063
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1679235063
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1679235063
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1679235063
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1679235063
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1679235063
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1679235063
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1679235063
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1679235063
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1679235063
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1679235063
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_23
timestamp 1679235063
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_35
timestamp 1679235063
transform 1 0 4324 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_42
timestamp 1679235063
transform 1 0 4968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1679235063
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1679235063
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1679235063
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1679235063
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1679235063
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1679235063
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_143
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1679235063
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1679235063
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1679235063
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1679235063
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_191
timestamp 1679235063
transform 1 0 18676 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1679235063
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1679235063
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_255
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_267
timestamp 1679235063
transform 1 0 25668 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_279
timestamp 1679235063
transform 1 0 26772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_291
timestamp 1679235063
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1679235063
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1679235063
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1679235063
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1679235063
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1679235063
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1679235063
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1679235063
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1679235063
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1679235063
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1679235063
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1679235063
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1679235063
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1679235063
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1679235063
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1679235063
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1679235063
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1679235063
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1679235063
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1679235063
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1679235063
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1679235063
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1679235063
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1679235063
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1679235063
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1679235063
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_31
timestamp 1679235063
transform 1 0 3956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1679235063
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1679235063
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1679235063
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_60
timestamp 1679235063
transform 1 0 6624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1679235063
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1679235063
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_105
timestamp 1679235063
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_120
timestamp 1679235063
transform 1 0 12144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_133
timestamp 1679235063
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1679235063
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1679235063
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1679235063
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_174
timestamp 1679235063
transform 1 0 17112 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_180
timestamp 1679235063
transform 1 0 17664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1679235063
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_205
timestamp 1679235063
transform 1 0 19964 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_231
timestamp 1679235063
transform 1 0 22356 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1679235063
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1679235063
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1679235063
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1679235063
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1679235063
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1679235063
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1679235063
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1679235063
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1679235063
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1679235063
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1679235063
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1679235063
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1679235063
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1679235063
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1679235063
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1679235063
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1679235063
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1679235063
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1679235063
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1679235063
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1679235063
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1679235063
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1679235063
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1679235063
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1679235063
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1679235063
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1679235063
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1679235063
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1679235063
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1679235063
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1679235063
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1679235063
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_31
timestamp 1679235063
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1679235063
transform 1 0 6532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1679235063
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1679235063
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1679235063
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1679235063
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1679235063
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_201
timestamp 1679235063
transform 1 0 19596 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_229
timestamp 1679235063
transform 1 0 22172 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_234
timestamp 1679235063
transform 1 0 22632 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_245
timestamp 1679235063
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_266
timestamp 1679235063
transform 1 0 25576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_278
timestamp 1679235063
transform 1 0 26680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1679235063
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1679235063
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1679235063
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1679235063
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1679235063
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1679235063
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1679235063
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1679235063
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1679235063
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1679235063
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1679235063
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1679235063
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1679235063
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1679235063
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1679235063
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1679235063
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1679235063
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1679235063
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1679235063
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1679235063
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1679235063
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1679235063
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1679235063
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1679235063
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1679235063
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_28
timestamp 1679235063
transform 1 0 3680 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1679235063
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1679235063
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1679235063
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1679235063
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1679235063
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1679235063
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1679235063
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1679235063
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1679235063
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_171
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1679235063
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1679235063
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1679235063
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1679235063
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1679235063
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_227
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1679235063
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1679235063
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1679235063
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1679235063
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1679235063
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1679235063
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1679235063
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1679235063
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1679235063
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1679235063
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1679235063
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1679235063
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1679235063
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1679235063
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1679235063
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1679235063
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1679235063
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1679235063
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1679235063
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1679235063
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1679235063
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1679235063
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1679235063
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1679235063
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1679235063
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1679235063
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1679235063
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1679235063
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1679235063
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1679235063
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_21
timestamp 1679235063
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1679235063
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1679235063
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1679235063
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_72
timestamp 1679235063
transform 1 0 7728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1679235063
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1679235063
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1679235063
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1679235063
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1679235063
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_191
timestamp 1679235063
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1679235063
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1679235063
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_210
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_220
timestamp 1679235063
transform 1 0 21344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1679235063
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1679235063
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_277
timestamp 1679235063
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_283
timestamp 1679235063
transform 1 0 27140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_295
timestamp 1679235063
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1679235063
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1679235063
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1679235063
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1679235063
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1679235063
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1679235063
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1679235063
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1679235063
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1679235063
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1679235063
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1679235063
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1679235063
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1679235063
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1679235063
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1679235063
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1679235063
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1679235063
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1679235063
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1679235063
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1679235063
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1679235063
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1679235063
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1679235063
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1679235063
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1679235063
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1679235063
transform 1 0 3404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1679235063
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1679235063
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_63
timestamp 1679235063
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1679235063
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1679235063
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1679235063
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1679235063
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1679235063
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_171
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1679235063
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1679235063
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_211
timestamp 1679235063
transform 1 0 20516 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1679235063
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1679235063
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1679235063
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_257
timestamp 1679235063
transform 1 0 24748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1679235063
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_283
timestamp 1679235063
transform 1 0 27140 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_295
timestamp 1679235063
transform 1 0 28244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_307
timestamp 1679235063
transform 1 0 29348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_319
timestamp 1679235063
transform 1 0 30452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 1679235063
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1679235063
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1679235063
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1679235063
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1679235063
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1679235063
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1679235063
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1679235063
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1679235063
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1679235063
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1679235063
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1679235063
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1679235063
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1679235063
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1679235063
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1679235063
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1679235063
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1679235063
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1679235063
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1679235063
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1679235063
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1679235063
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1679235063
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_21
timestamp 1679235063
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1679235063
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1679235063
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1679235063
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1679235063
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1679235063
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1679235063
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1679235063
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_128
timestamp 1679235063
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1679235063
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1679235063
transform 1 0 15272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1679235063
transform 1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1679235063
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1679235063
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_202
timestamp 1679235063
transform 1 0 19688 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1679235063
transform 1 0 20056 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1679235063
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_234
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_237
timestamp 1679235063
transform 1 0 22908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_255
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1679235063
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_271
timestamp 1679235063
transform 1 0 26036 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1679235063
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1679235063
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1679235063
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1679235063
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1679235063
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1679235063
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1679235063
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1679235063
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1679235063
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1679235063
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1679235063
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1679235063
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1679235063
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1679235063
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1679235063
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1679235063
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1679235063
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1679235063
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1679235063
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1679235063
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1679235063
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1679235063
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1679235063
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1679235063
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1679235063
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1679235063
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1679235063
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1679235063
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1679235063
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_63
timestamp 1679235063
transform 1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1679235063
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1679235063
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1679235063
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1679235063
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1679235063
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1679235063
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1679235063
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1679235063
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1679235063
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1679235063
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1679235063
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1679235063
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1679235063
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1679235063
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_250
timestamp 1679235063
transform 1 0 24104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_256
timestamp 1679235063
transform 1 0 24656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1679235063
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_283
timestamp 1679235063
transform 1 0 27140 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_295
timestamp 1679235063
transform 1 0 28244 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_307
timestamp 1679235063
transform 1 0 29348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_319
timestamp 1679235063
transform 1 0 30452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1679235063
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1679235063
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1679235063
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1679235063
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1679235063
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1679235063
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1679235063
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1679235063
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1679235063
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1679235063
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1679235063
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1679235063
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1679235063
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1679235063
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1679235063
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1679235063
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1679235063
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1679235063
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1679235063
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1679235063
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1679235063
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1679235063
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1679235063
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1679235063
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1679235063
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_59
timestamp 1679235063
transform 1 0 6532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1679235063
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_91
timestamp 1679235063
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_95
timestamp 1679235063
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1679235063
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1679235063
transform 1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1679235063
transform 1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1679235063
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1679235063
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1679235063
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1679235063
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1679235063
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1679235063
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1679235063
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_226
timestamp 1679235063
transform 1 0 21896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1679235063
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1679235063
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_265
timestamp 1679235063
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_271
timestamp 1679235063
transform 1 0 26036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1679235063
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_299
timestamp 1679235063
transform 1 0 28612 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1679235063
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1679235063
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1679235063
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1679235063
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1679235063
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1679235063
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1679235063
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1679235063
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1679235063
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1679235063
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1679235063
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1679235063
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1679235063
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1679235063
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1679235063
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1679235063
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1679235063
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1679235063
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1679235063
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1679235063
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1679235063
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1679235063
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1679235063
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1679235063
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1679235063
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1679235063
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1679235063
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1679235063
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1679235063
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_84
timestamp 1679235063
transform 1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1679235063
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1679235063
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1679235063
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1679235063
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1679235063
transform 1 0 12420 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_133
timestamp 1679235063
transform 1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1679235063
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp 1679235063
transform 1 0 15272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1679235063
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1679235063
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1679235063
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1679235063
transform 1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1679235063
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1679235063
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_240
timestamp 1679235063
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_250
timestamp 1679235063
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1679235063
transform 1 0 24472 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_276
timestamp 1679235063
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1679235063
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1679235063
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_310
timestamp 1679235063
transform 1 0 29624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_314
timestamp 1679235063
transform 1 0 29992 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_324
timestamp 1679235063
transform 1 0 30912 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1679235063
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1679235063
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1679235063
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1679235063
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1679235063
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1679235063
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1679235063
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1679235063
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1679235063
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1679235063
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1679235063
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1679235063
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1679235063
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1679235063
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1679235063
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1679235063
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1679235063
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1679235063
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1679235063
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1679235063
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1679235063
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1679235063
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1679235063
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1679235063
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1679235063
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1679235063
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1679235063
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1679235063
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1679235063
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1679235063
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1679235063
transform 1 0 14628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1679235063
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_158
timestamp 1679235063
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1679235063
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1679235063
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_189
timestamp 1679235063
transform 1 0 18492 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1679235063
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_222
timestamp 1679235063
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1679235063
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_255
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1679235063
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1679235063
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1679235063
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1679235063
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1679235063
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_333
timestamp 1679235063
transform 1 0 31740 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_337
timestamp 1679235063
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_349
timestamp 1679235063
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1679235063
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1679235063
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1679235063
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1679235063
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1679235063
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1679235063
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1679235063
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1679235063
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1679235063
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1679235063
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1679235063
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1679235063
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1679235063
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1679235063
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1679235063
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1679235063
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1679235063
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1679235063
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1679235063
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1679235063
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_79
timestamp 1679235063
transform 1 0 8372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1679235063
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1679235063
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1679235063
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_127
timestamp 1679235063
transform 1 0 12788 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_134
timestamp 1679235063
transform 1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1679235063
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1679235063
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1679235063
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1679235063
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_192
timestamp 1679235063
transform 1 0 18768 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1679235063
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1679235063
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_230
timestamp 1679235063
transform 1 0 22264 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_234
timestamp 1679235063
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1679235063
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1679235063
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1679235063
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1679235063
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_286
timestamp 1679235063
transform 1 0 27416 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_292
timestamp 1679235063
transform 1 0 27968 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1679235063
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_326
timestamp 1679235063
transform 1 0 31096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1679235063
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1679235063
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1679235063
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1679235063
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1679235063
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1679235063
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1679235063
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1679235063
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1679235063
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1679235063
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1679235063
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1679235063
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1679235063
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1679235063
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1679235063
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1679235063
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1679235063
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1679235063
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1679235063
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1679235063
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1679235063
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1679235063
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1679235063
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1679235063
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_99
timestamp 1679235063
transform 1 0 10212 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp 1679235063
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1679235063
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1679235063
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1679235063
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_177
timestamp 1679235063
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1679235063
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1679235063
transform 1 0 20608 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_216
timestamp 1679235063
transform 1 0 20976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1679235063
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_245
timestamp 1679235063
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1679235063
transform 1 0 24840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_262
timestamp 1679235063
transform 1 0 25208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1679235063
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1679235063
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1679235063
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1679235063
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1679235063
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_324
timestamp 1679235063
transform 1 0 30912 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_336
timestamp 1679235063
transform 1 0 32016 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_348
timestamp 1679235063
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1679235063
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1679235063
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1679235063
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1679235063
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1679235063
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1679235063
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1679235063
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1679235063
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1679235063
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1679235063
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1679235063
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1679235063
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1679235063
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1679235063
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1679235063
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1679235063
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1679235063
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1679235063
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1679235063
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1679235063
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1679235063
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1679235063
transform 1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_135
timestamp 1679235063
transform 1 0 13524 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_161
timestamp 1679235063
transform 1 0 15916 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1679235063
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1679235063
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1679235063
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1679235063
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_243
timestamp 1679235063
transform 1 0 23460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1679235063
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1679235063
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1679235063
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_274
timestamp 1679235063
transform 1 0 26312 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1679235063
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_283
timestamp 1679235063
transform 1 0 27140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_288
timestamp 1679235063
transform 1 0 27600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_293
timestamp 1679235063
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_315
timestamp 1679235063
transform 1 0 30084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_322
timestamp 1679235063
transform 1 0 30728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1679235063
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1679235063
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1679235063
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1679235063
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1679235063
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1679235063
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1679235063
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1679235063
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1679235063
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1679235063
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1679235063
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1679235063
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1679235063
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1679235063
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1679235063
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1679235063
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1679235063
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1679235063
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1679235063
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1679235063
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1679235063
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1679235063
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_21
timestamp 1679235063
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_35
timestamp 1679235063
transform 1 0 4324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1679235063
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1679235063
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_107
timestamp 1679235063
transform 1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1679235063
transform 1 0 11592 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1679235063
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_166
timestamp 1679235063
transform 1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1679235063
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_184
timestamp 1679235063
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1679235063
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1679235063
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1679235063
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1679235063
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1679235063
transform 1 0 23184 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_289
timestamp 1679235063
transform 1 0 27692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_293
timestamp 1679235063
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1679235063
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1679235063
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_314
timestamp 1679235063
transform 1 0 29992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_320
timestamp 1679235063
transform 1 0 30544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_331
timestamp 1679235063
transform 1 0 31556 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_335
timestamp 1679235063
transform 1 0 31924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_347
timestamp 1679235063
transform 1 0 33028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1679235063
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1679235063
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1679235063
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1679235063
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1679235063
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1679235063
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1679235063
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1679235063
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1679235063
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1679235063
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1679235063
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1679235063
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1679235063
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1679235063
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1679235063
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1679235063
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1679235063
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1679235063
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1679235063
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1679235063
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1679235063
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_75
timestamp 1679235063
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_80
timestamp 1679235063
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1679235063
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1679235063
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_123
timestamp 1679235063
transform 1 0 12420 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1679235063
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_182
timestamp 1679235063
transform 1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1679235063
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1679235063
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1679235063
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_245
timestamp 1679235063
transform 1 0 23644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_250
timestamp 1679235063
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_272
timestamp 1679235063
transform 1 0 26128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1679235063
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1679235063
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1679235063
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1679235063
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1679235063
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_347
timestamp 1679235063
transform 1 0 33028 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_359
timestamp 1679235063
transform 1 0 34132 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_371
timestamp 1679235063
transform 1 0 35236 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_383
timestamp 1679235063
transform 1 0 36340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1679235063
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1679235063
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1679235063
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1679235063
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1679235063
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1679235063
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1679235063
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1679235063
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1679235063
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1679235063
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1679235063
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1679235063
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1679235063
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1679235063
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1679235063
transform 1 0 48668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1679235063
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1679235063
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_45
timestamp 1679235063
transform 1 0 5244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1679235063
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_103
timestamp 1679235063
transform 1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_108
timestamp 1679235063
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_114
timestamp 1679235063
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_144
timestamp 1679235063
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1679235063
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1679235063
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1679235063
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_219
timestamp 1679235063
transform 1 0 21252 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_226
timestamp 1679235063
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1679235063
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_269
timestamp 1679235063
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1679235063
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1679235063
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1679235063
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_321
timestamp 1679235063
transform 1 0 30636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1679235063
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_337
timestamp 1679235063
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_344
timestamp 1679235063
transform 1 0 32752 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_350
timestamp 1679235063
transform 1 0 33304 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_356
timestamp 1679235063
transform 1 0 33856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1679235063
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1679235063
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1679235063
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1679235063
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1679235063
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1679235063
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1679235063
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1679235063
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1679235063
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1679235063
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1679235063
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1679235063
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1679235063
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1679235063
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1679235063
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1679235063
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1679235063
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_41
timestamp 1679235063
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_61
timestamp 1679235063
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_67
timestamp 1679235063
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_91
timestamp 1679235063
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_104
timestamp 1679235063
transform 1 0 10672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1679235063
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_129
timestamp 1679235063
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_150
timestamp 1679235063
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1679235063
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1679235063
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_211
timestamp 1679235063
transform 1 0 20516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_217
timestamp 1679235063
transform 1 0 21068 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_275
timestamp 1679235063
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1679235063
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1679235063
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1679235063
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_330
timestamp 1679235063
transform 1 0 31464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1679235063
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1679235063
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_350
timestamp 1679235063
transform 1 0 33304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_354
timestamp 1679235063
transform 1 0 33672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_360
timestamp 1679235063
transform 1 0 34224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_368
timestamp 1679235063
transform 1 0 34960 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_372
timestamp 1679235063
transform 1 0 35328 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_375
timestamp 1679235063
transform 1 0 35604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1679235063
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1679235063
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1679235063
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1679235063
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1679235063
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1679235063
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1679235063
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1679235063
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1679235063
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1679235063
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1679235063
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1679235063
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1679235063
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1679235063
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_507
timestamp 1679235063
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1679235063
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_47
timestamp 1679235063
transform 1 0 5428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1679235063
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_57
timestamp 1679235063
transform 1 0 6348 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1679235063
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_78
timestamp 1679235063
transform 1 0 8280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1679235063
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_147
timestamp 1679235063
transform 1 0 14628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1679235063
transform 1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1679235063
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_173
timestamp 1679235063
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1679235063
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1679235063
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_225
timestamp 1679235063
transform 1 0 21804 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_229
timestamp 1679235063
transform 1 0 22172 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_232
timestamp 1679235063
transform 1 0 22448 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1679235063
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1679235063
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1679235063
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_302
timestamp 1679235063
transform 1 0 28888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_313
timestamp 1679235063
transform 1 0 29900 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_324
timestamp 1679235063
transform 1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_332
timestamp 1679235063
transform 1 0 31648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_340
timestamp 1679235063
transform 1 0 32384 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_352
timestamp 1679235063
transform 1 0 33488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_360
timestamp 1679235063
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1679235063
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_371
timestamp 1679235063
transform 1 0 35236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_378
timestamp 1679235063
transform 1 0 35880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_385
timestamp 1679235063
transform 1 0 36524 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_393
timestamp 1679235063
transform 1 0 37260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_398
timestamp 1679235063
transform 1 0 37720 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_402
timestamp 1679235063
transform 1 0 38088 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_408
timestamp 1679235063
transform 1 0 38640 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_412
timestamp 1679235063
transform 1 0 39008 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1679235063
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1679235063
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1679235063
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1679235063
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1679235063
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1679235063
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1679235063
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1679235063
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1679235063
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1679235063
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_513
timestamp 1679235063
transform 1 0 48300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_517
timestamp 1679235063
transform 1 0 48668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1679235063
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1679235063
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1679235063
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1679235063
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1679235063
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1679235063
transform 1 0 14260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1679235063
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1679235063
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_230
timestamp 1679235063
transform 1 0 22264 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1679235063
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1679235063
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1679235063
transform 1 0 26128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1679235063
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1679235063
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1679235063
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_329
timestamp 1679235063
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1679235063
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1679235063
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_343
timestamp 1679235063
transform 1 0 32660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_351
timestamp 1679235063
transform 1 0 33396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_357
timestamp 1679235063
transform 1 0 33948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_370
timestamp 1679235063
transform 1 0 35144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_378
timestamp 1679235063
transform 1 0 35880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_386
timestamp 1679235063
transform 1 0 36616 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1679235063
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_397
timestamp 1679235063
transform 1 0 37628 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_419
timestamp 1679235063
transform 1 0 39652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_427
timestamp 1679235063
transform 1 0 40388 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_433
timestamp 1679235063
transform 1 0 40940 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_440
timestamp 1679235063
transform 1 0 41584 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1679235063
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1679235063
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_459
timestamp 1679235063
transform 1 0 43332 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1679235063
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1679235063
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1679235063
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1679235063
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1679235063
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_517
timestamp 1679235063
transform 1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1679235063
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp 1679235063
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1679235063
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_87
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1679235063
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_133
timestamp 1679235063
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_147
timestamp 1679235063
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_152
timestamp 1679235063
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1679235063
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1679235063
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_277
timestamp 1679235063
transform 1 0 26588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_281
timestamp 1679235063
transform 1 0 26956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_304
timestamp 1679235063
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1679235063
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_331
timestamp 1679235063
transform 1 0 31556 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_338
timestamp 1679235063
transform 1 0 32200 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_344
timestamp 1679235063
transform 1 0 32752 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_349
timestamp 1679235063
transform 1 0 33212 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_355
timestamp 1679235063
transform 1 0 33764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1679235063
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1679235063
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_371
timestamp 1679235063
transform 1 0 35236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_378
timestamp 1679235063
transform 1 0 35880 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_382
timestamp 1679235063
transform 1 0 36248 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_405
timestamp 1679235063
transform 1 0 38364 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_412
timestamp 1679235063
transform 1 0 39008 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_416
timestamp 1679235063
transform 1 0 39376 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1679235063
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1679235063
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_445
timestamp 1679235063
transform 1 0 42044 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_451
timestamp 1679235063
transform 1 0 42596 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_455
timestamp 1679235063
transform 1 0 42964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_467
timestamp 1679235063
transform 1 0 44068 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1679235063
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1679235063
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_489
timestamp 1679235063
transform 1 0 46092 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_498
timestamp 1679235063
transform 1 0 46920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_502
timestamp 1679235063
transform 1 0 47288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_507
timestamp 1679235063
transform 1 0 47748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_513
timestamp 1679235063
transform 1 0 48300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1679235063
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_8
timestamp 1679235063
transform 1 0 1840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1679235063
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_115
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1679235063
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1679235063
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1679235063
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_219
timestamp 1679235063
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1679235063
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1679235063
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1679235063
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1679235063
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1679235063
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_310
timestamp 1679235063
transform 1 0 29624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_318
timestamp 1679235063
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_324
timestamp 1679235063
transform 1 0 30912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_331
timestamp 1679235063
transform 1 0 31556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1679235063
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1679235063
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_347
timestamp 1679235063
transform 1 0 33028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_355
timestamp 1679235063
transform 1 0 33764 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_362
timestamp 1679235063
transform 1 0 34408 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_374
timestamp 1679235063
transform 1 0 35512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_382
timestamp 1679235063
transform 1 0 36248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1679235063
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1679235063
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_398
timestamp 1679235063
transform 1 0 37720 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_402
timestamp 1679235063
transform 1 0 38088 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_409
timestamp 1679235063
transform 1 0 38732 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_417
timestamp 1679235063
transform 1 0 39468 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_421
timestamp 1679235063
transform 1 0 39836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_430
timestamp 1679235063
transform 1 0 40664 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_436
timestamp 1679235063
transform 1 0 41216 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1679235063
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1679235063
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_459
timestamp 1679235063
transform 1 0 43332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_471
timestamp 1679235063
transform 1 0 44436 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_479
timestamp 1679235063
transform 1 0 45172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_487
timestamp 1679235063
transform 1 0 45908 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_493
timestamp 1679235063
transform 1 0 46460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1679235063
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_507
timestamp 1679235063
transform 1 0 47748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_513
timestamp 1679235063
transform 1 0 48300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1679235063
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1679235063
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1679235063
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_191
timestamp 1679235063
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1679235063
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_277
timestamp 1679235063
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1679235063
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_292
timestamp 1679235063
transform 1 0 27968 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_296
timestamp 1679235063
transform 1 0 28336 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1679235063
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1679235063
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1679235063
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_333
timestamp 1679235063
transform 1 0 31740 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1679235063
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_347
timestamp 1679235063
transform 1 0 33028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_359
timestamp 1679235063
transform 1 0 34132 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1679235063
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1679235063
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_375
timestamp 1679235063
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_387
timestamp 1679235063
transform 1 0 36708 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_391
timestamp 1679235063
transform 1 0 37076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1679235063
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_398
timestamp 1679235063
transform 1 0 37720 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_404
timestamp 1679235063
transform 1 0 38272 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_414
timestamp 1679235063
transform 1 0 39192 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1679235063
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_431
timestamp 1679235063
transform 1 0 40756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_443
timestamp 1679235063
transform 1 0 41860 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_447
timestamp 1679235063
transform 1 0 42228 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_451
timestamp 1679235063
transform 1 0 42596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_463
timestamp 1679235063
transform 1 0 43700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_467
timestamp 1679235063
transform 1 0 44068 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_471
timestamp 1679235063
transform 1 0 44436 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1679235063
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1679235063
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1679235063
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1679235063
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1679235063
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1679235063
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1679235063
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_515
timestamp 1679235063
transform 1 0 48484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_524
timestamp 1679235063
transform 1 0 49312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 43700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold2
timestamp 1679235063
transform 1 0 42688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 41400 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 43332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 42596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold6
timestamp 1679235063
transform 1 0 36524 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 42596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 48576 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 43884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 2944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 6532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 28244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 37444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold15
timestamp 1679235063
transform 1 0 35236 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 25576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold17
timestamp 1679235063
transform 1 0 37812 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 30912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold19
timestamp 1679235063
transform 1 0 35696 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 28520 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 32292 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 2852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 35972 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 33396 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 34776 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 41124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 34868 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 38456 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 39928 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 40020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 2668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 31004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 32292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 1564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 48668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 48668 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 46184 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 1840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 4600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 48392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1679235063
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1679235063
transform 1 0 1564 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 3496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 2852 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1679235063
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1679235063
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1679235063
transform 1 0 1564 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1679235063
transform 1 0 1564 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1679235063
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1679235063
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1679235063
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1679235063
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1679235063
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1679235063
transform 1 0 33028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1679235063
transform 1 0 29716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1679235063
transform 1 0 30544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 32936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 35604 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1679235063
transform 1 0 36616 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 37444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1679235063
transform 1 0 33396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1679235063
transform 1 0 33948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1679235063
transform 1 0 34868 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1679235063
transform 1 0 35880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1679235063
transform 1 0 38732 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 37444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 37444 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 38732 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1679235063
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1679235063
transform 1 0 39100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1679235063
transform 1 0 40020 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 40664 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1679235063
transform 1 0 41308 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 31924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1679235063
transform 1 0 34132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1679235063
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1679235063
transform 1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 33488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 36064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1679235063
transform 1 0 44160 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1679235063
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1679235063
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1679235063
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1679235063
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1679235063
transform 1 0 47932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1679235063
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1679235063
transform 1 0 45540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1679235063
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1679235063
transform 1 0 49036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1679235063
transform 1 0 48300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1679235063
transform 1 0 47932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 8372 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 3404 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 10488 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 11960 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 15180 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 7912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 4140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 6808 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 12144 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 14812 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform 1 0 17480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18676 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20240 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21160 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18676 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20056 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24288 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25852 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 26036 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27232 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28336 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28336 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28244 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28060 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37812 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27784 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24840 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20884 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20332 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 20240 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 20056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16008 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14444 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14720 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16284 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14536 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14628 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12052 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11500 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11960 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6716 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 4876 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 4600 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 4508 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7636 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11500 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12420 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13708 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15180 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18124 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30728 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 27784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__194
timestamp 1679235063
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17204 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__160
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11224 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__162
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18492 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6808 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__195
timestamp 1679235063
transform 1 0 35604 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__196
timestamp 1679235063
transform 1 0 36248 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 31004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__197
timestamp 1679235063
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 28336 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25760 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15732 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__198
timestamp 1679235063
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__151
timestamp 1679235063
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__152
timestamp 1679235063
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27232 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__154
timestamp 1679235063
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30544 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__156
timestamp 1679235063
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30084 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__157
timestamp 1679235063
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25576 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__158
timestamp 1679235063
transform 1 0 26404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30544 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__159
timestamp 1679235063
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30912 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__161
timestamp 1679235063
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 26588 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__164
timestamp 1679235063
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23644 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23368 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__170
timestamp 1679235063
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 22172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17756 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__181
timestamp 1679235063
transform 1 0 12604 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12144 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__188
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24656 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__189
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__165
timestamp 1679235063
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20516 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__166
timestamp 1679235063
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14260 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__167
timestamp 1679235063
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10120 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__168
timestamp 1679235063
transform 1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__169
timestamp 1679235063
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15824 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__171
timestamp 1679235063
transform 1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__172
timestamp 1679235063
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13708 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__173
timestamp 1679235063
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__174
timestamp 1679235063
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10304 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__175
timestamp 1679235063
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11316 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__176
timestamp 1679235063
transform 1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__177
timestamp 1679235063
transform 1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 32476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12512 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__178
timestamp 1679235063
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 30452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11592 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__179
timestamp 1679235063
transform 1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 4140 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__180
timestamp 1679235063
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 6716 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__182
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__183
timestamp 1679235063
transform 1 0 33580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17848 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 9844 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__184
timestamp 1679235063
transform 1 0 4140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__185
timestamp 1679235063
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 32568 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13708 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__186
timestamp 1679235063
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 27600 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__187
timestamp 1679235063
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40866 26200 40922 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 41510 26200 41566 27000 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 test_enable
port 142 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 22856 51000 22976 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 24760 51000 24880 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 17526 6188 17526 6188 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 12466 6188 12466 6188 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 14812 5746 14812 5746 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 9614 7956 9614 7956 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20884 17714 20884 17714 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 8694 9894 8694 9894 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal2 21482 15912 21482 15912 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 10948 13838 10948 13838 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 8602 9010 8602 9010 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 5704 12138 5704 12138 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal2 10074 17884 10074 17884 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 6670 12750 6670 12750 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 5842 13804 5842 13804 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal2 9660 12580 9660 12580 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal2 6532 21420 6532 21420 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 12650 15589 12650 15589 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 9752 13430 9752 13430 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 5842 17136 5842 17136 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 13662 17578 13662 17578 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 9384 18870 9384 18870 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 8832 14382 8832 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8786 9146 8786 9146 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13570 9384 13570 9384 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 8234 14450 8234 14450 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9062 15776 9062 15776 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10442 15130 10442 15130 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11546 14042 11546 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8096 11186 8096 11186 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8878 14858 8878 14858 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8970 8058 8970 8058 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 8234 9316 8234 9316 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10396 9622 10396 9622 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4416 14042 4416 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4876 11866 4876 11866 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 10810 7412 10810 7412 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 4922 14382 4922 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6808 15538 6808 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7544 15402 7544 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8970 12954 8970 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5566 13974 5566 13974 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6026 14042 6026 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 6302 11798 6302 11798 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 5382 12614 5382 12614 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 4922 11730 4922 11730 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 5612 15538 5612 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9522 11458 9522 11458 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 11362 9350 11362 9350 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 4784 15402 4784 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6348 13906 6348 13906 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7314 14416 7314 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9384 12206 9384 12206 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 8602 14229 8602 14229 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6946 14008 6946 14008 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9384 12410 9384 12410 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 12742 13634 12742 13634 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8694 14042 8694 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 8464 17578 8464 17578 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10488 17850 10488 17850 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 7084 13396 7084 13396 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 6302 20230 6302 20230 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6302 17306 6302 17306 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7866 16388 7866 16388 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10120 14382 10120 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7544 22610 7544 22610 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6992 22610 6992 22610 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 9430 15912 9430 15912 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 14398 18462 14398 18462 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 6256 22474 6256 22474 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 17434 4284 17434 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal2 17710 4114 17710 4114 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 20562 4012 20562 4012 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 26795 4794 26795 4794 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 19964 5882 19964 5882 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 15686 5134 15686 5134 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 18124 3026 18124 3026 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 25047 5338 25047 5338 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25806 7514 25806 7514 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 16468 5678 16468 5678 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 17066 4284 17066 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 24380 4522 24380 4522 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 15456 7854 15456 7854 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 15226 6052 15226 6052 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal2 24886 5916 24886 5916 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 1656 4114 1656 4114 0 ccff_head
rlabel metal1 48622 23086 48622 23086 0 ccff_head_1
rlabel metal2 49174 21233 49174 21233 0 ccff_tail
rlabel metal2 2254 24252 2254 24252 0 ccff_tail_0
rlabel metal3 1786 1564 1786 1564 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal3 1004 6052 1004 6052 0 chanx_left_in[11]
rlabel metal1 1794 5712 1794 5712 0 chanx_left_in[12]
rlabel metal1 4140 6766 4140 6766 0 chanx_left_in[13]
rlabel metal1 2944 6290 2944 6290 0 chanx_left_in[14]
rlabel metal2 3726 6987 3726 6987 0 chanx_left_in[15]
rlabel metal2 1334 7769 1334 7769 0 chanx_left_in[16]
rlabel metal1 4554 7854 4554 7854 0 chanx_left_in[17]
rlabel metal1 4554 7378 4554 7378 0 chanx_left_in[18]
rlabel metal3 1119 9316 1119 9316 0 chanx_left_in[19]
rlabel metal1 3082 2380 3082 2380 0 chanx_left_in[1]
rlabel metal2 2898 9095 2898 9095 0 chanx_left_in[20]
rlabel metal3 2254 10064 2254 10064 0 chanx_left_in[21]
rlabel metal1 2162 6800 2162 6800 0 chanx_left_in[22]
rlabel metal2 1610 9163 1610 9163 0 chanx_left_in[23]
rlabel metal1 1564 7922 1564 7922 0 chanx_left_in[24]
rlabel metal3 1004 11764 1004 11764 0 chanx_left_in[25]
rlabel metal1 1380 11730 1380 11730 0 chanx_left_in[26]
rlabel metal3 1717 12580 1717 12580 0 chanx_left_in[27]
rlabel metal2 1334 12937 1334 12937 0 chanx_left_in[28]
rlabel metal1 1656 12750 1656 12750 0 chanx_left_in[29]
rlabel metal1 2714 2482 2714 2482 0 chanx_left_in[2]
rlabel metal1 3174 2550 3174 2550 0 chanx_left_in[3]
rlabel metal3 1004 3196 1004 3196 0 chanx_left_in[4]
rlabel metal1 2990 4590 2990 4590 0 chanx_left_in[5]
rlabel metal1 4140 3502 4140 3502 0 chanx_left_in[6]
rlabel metal1 4232 4114 4232 4114 0 chanx_left_in[7]
rlabel metal1 1472 4658 1472 4658 0 chanx_left_in[8]
rlabel metal1 1472 5202 1472 5202 0 chanx_left_in[9]
rlabel metal3 1372 13804 1372 13804 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal2 2806 18819 2806 18819 0 chanx_left_out[11]
rlabel metal2 2898 19227 2898 19227 0 chanx_left_out[12]
rlabel metal3 1372 19108 1372 19108 0 chanx_left_out[13]
rlabel metal2 2806 20179 2806 20179 0 chanx_left_out[14]
rlabel metal3 1326 19924 1326 19924 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal2 2852 21148 2852 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal2 4094 22015 4094 22015 0 chanx_left_out[20]
rlabel metal3 1487 22372 1487 22372 0 chanx_left_out[21]
rlabel metal1 5842 20502 5842 20502 0 chanx_left_out[22]
rlabel metal1 3772 19754 3772 19754 0 chanx_left_out[23]
rlabel metal2 3818 23545 3818 23545 0 chanx_left_out[24]
rlabel metal2 4094 23800 4094 23800 0 chanx_left_out[25]
rlabel metal2 5198 19319 5198 19319 0 chanx_left_out[26]
rlabel metal1 8050 20026 8050 20026 0 chanx_left_out[27]
rlabel metal1 8924 19414 8924 19414 0 chanx_left_out[28]
rlabel metal2 3864 20468 3864 20468 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 912 15028 912 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal3 1372 17476 1372 17476 0 chanx_left_out[9]
rlabel via2 5382 7395 5382 7395 0 chany_top_in[0]
rlabel metal1 32568 20570 32568 20570 0 chany_top_in[10]
rlabel metal2 31050 24276 31050 24276 0 chany_top_in[11]
rlabel metal1 32338 24208 32338 24208 0 chany_top_in[12]
rlabel metal2 33166 23188 33166 23188 0 chany_top_in[13]
rlabel metal1 35650 21998 35650 21998 0 chany_top_in[14]
rlabel metal2 36846 23426 36846 23426 0 chany_top_in[15]
rlabel metal1 37398 23698 37398 23698 0 chany_top_in[16]
rlabel metal1 33810 21114 33810 21114 0 chany_top_in[17]
rlabel metal1 34868 24174 34868 24174 0 chany_top_in[18]
rlabel metal1 34684 23698 34684 23698 0 chany_top_in[19]
rlabel metal1 30590 22066 30590 22066 0 chany_top_in[1]
rlabel metal1 35558 24174 35558 24174 0 chany_top_in[20]
rlabel metal1 37352 23086 37352 23086 0 chany_top_in[21]
rlabel metal1 37030 24174 37030 24174 0 chany_top_in[22]
rlabel metal1 37490 21998 37490 21998 0 chany_top_in[23]
rlabel metal1 39100 22066 39100 22066 0 chany_top_in[24]
rlabel metal2 38502 25245 38502 25245 0 chany_top_in[25]
rlabel metal1 39514 24174 39514 24174 0 chany_top_in[26]
rlabel metal1 39790 23698 39790 23698 0 chany_top_in[27]
rlabel metal2 40250 25238 40250 25238 0 chany_top_in[28]
rlabel metal1 41538 22644 41538 22644 0 chany_top_in[29]
rlabel metal3 17204 23256 17204 23256 0 chany_top_in[2]
rlabel metal2 598 20468 598 20468 0 chany_top_in[3]
rlabel metal1 14536 24174 14536 24174 0 chany_top_in[4]
rlabel metal2 20746 22780 20746 22780 0 chany_top_in[5]
rlabel metal1 32338 20434 32338 20434 0 chany_top_in[6]
rlabel metal1 29532 23698 29532 23698 0 chany_top_in[7]
rlabel metal2 32062 23936 32062 23936 0 chany_top_in[8]
rlabel metal2 32246 23494 32246 23494 0 chany_top_in[9]
rlabel metal1 3818 22134 3818 22134 0 chany_top_out[0]
rlabel metal1 8786 24242 8786 24242 0 chany_top_out[10]
rlabel metal1 9568 23766 9568 23766 0 chany_top_out[11]
rlabel metal2 10718 24497 10718 24497 0 chany_top_out[12]
rlabel metal2 11270 24184 11270 24184 0 chany_top_out[13]
rlabel metal2 12650 21964 12650 21964 0 chany_top_out[14]
rlabel metal2 12558 25034 12558 25034 0 chany_top_out[15]
rlabel metal2 13301 26316 13301 26316 0 chany_top_out[16]
rlabel metal2 13846 25204 13846 25204 0 chany_top_out[17]
rlabel metal1 13984 24242 13984 24242 0 chany_top_out[18]
rlabel metal1 15410 22066 15410 22066 0 chany_top_out[19]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[1]
rlabel metal1 15042 23766 15042 23766 0 chany_top_out[20]
rlabel metal2 16146 24497 16146 24497 0 chany_top_out[21]
rlabel metal2 17211 26316 17211 26316 0 chany_top_out[22]
rlabel metal1 16974 23154 16974 23154 0 chany_top_out[23]
rlabel metal1 17250 23630 17250 23630 0 chany_top_out[24]
rlabel metal1 16468 24242 16468 24242 0 chany_top_out[25]
rlabel metal1 18584 23766 18584 23766 0 chany_top_out[26]
rlabel metal1 20792 21930 20792 21930 0 chany_top_out[27]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[28]
rlabel metal2 22034 25296 22034 25296 0 chany_top_out[29]
rlabel metal1 4094 23766 4094 23766 0 chany_top_out[2]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[3]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[4]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[5]
rlabel metal1 7038 22134 7038 22134 0 chany_top_out[6]
rlabel metal1 6624 24242 6624 24242 0 chany_top_out[7]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[8]
rlabel metal2 8694 24422 8694 24422 0 chany_top_out[9]
rlabel metal2 18446 17408 18446 17408 0 clknet_0_prog_clk
rlabel metal1 8004 9486 8004 9486 0 clknet_4_0_0_prog_clk
rlabel metal1 26174 13226 26174 13226 0 clknet_4_10_0_prog_clk
rlabel metal2 22034 16320 22034 16320 0 clknet_4_11_0_prog_clk
rlabel metal2 16330 18496 16330 18496 0 clknet_4_12_0_prog_clk
rlabel metal1 19734 20502 19734 20502 0 clknet_4_13_0_prog_clk
rlabel metal1 25852 19822 25852 19822 0 clknet_4_14_0_prog_clk
rlabel metal1 37628 22610 37628 22610 0 clknet_4_15_0_prog_clk
rlabel metal1 6762 13294 6762 13294 0 clknet_4_1_0_prog_clk
rlabel metal1 14536 10030 14536 10030 0 clknet_4_2_0_prog_clk
rlabel metal2 14306 13090 14306 13090 0 clknet_4_3_0_prog_clk
rlabel metal1 4554 17646 4554 17646 0 clknet_4_4_0_prog_clk
rlabel metal1 9430 20298 9430 20298 0 clknet_4_5_0_prog_clk
rlabel metal2 14582 19652 14582 19652 0 clknet_4_6_0_prog_clk
rlabel metal1 12834 21522 12834 21522 0 clknet_4_7_0_prog_clk
rlabel metal2 16882 7616 16882 7616 0 clknet_4_8_0_prog_clk
rlabel metal1 19964 12750 19964 12750 0 clknet_4_9_0_prog_clk
rlabel metal2 4094 1622 4094 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 1622 6762 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 9430 1622 9430 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12098 1622 12098 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 25392 2278 25392 2278 0 gfpga_pad_io_soc_in[0]
rlabel metal1 27876 2278 27876 2278 0 gfpga_pad_io_soc_in[1]
rlabel metal1 30728 2278 30728 2278 0 gfpga_pad_io_soc_in[2]
rlabel metal1 33396 2278 33396 2278 0 gfpga_pad_io_soc_in[3]
rlabel metal2 14766 1622 14766 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 17434 1622 17434 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 20102 959 20102 959 0 gfpga_pad_io_soc_out[2]
rlabel metal2 22770 1622 22770 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 36110 1588 36110 1588 0 isol_n
rlabel metal1 4646 3060 4646 3060 0 net1
rlabel metal2 12558 16966 12558 16966 0 net10
rlabel metal1 4462 17170 4462 17170 0 net100
rlabel metal1 4600 16558 4600 16558 0 net101
rlabel metal1 13570 18360 13570 18360 0 net102
rlabel metal1 8694 19346 8694 19346 0 net103
rlabel metal2 3542 15606 3542 15606 0 net104
rlabel metal2 1794 16609 1794 16609 0 net105
rlabel metal2 14490 17561 14490 17561 0 net106
rlabel metal2 3450 14756 3450 14756 0 net107
rlabel metal1 2277 16082 2277 16082 0 net108
rlabel metal1 2898 16558 2898 16558 0 net109
rlabel metal1 11546 16966 11546 16966 0 net11
rlabel metal1 2277 17170 2277 17170 0 net110
rlabel metal1 1794 17680 1794 17680 0 net111
rlabel metal1 2024 18258 2024 18258 0 net112
rlabel metal2 1196 16932 1196 16932 0 net113
rlabel metal1 7636 7922 7636 7922 0 net114
rlabel metal2 7728 17238 7728 17238 0 net115
rlabel metal2 20654 22168 20654 22168 0 net116
rlabel metal2 36570 23766 36570 23766 0 net117
rlabel metal1 34040 21318 34040 21318 0 net118
rlabel metal2 19596 18700 19596 18700 0 net119
rlabel metal1 6164 7514 6164 7514 0 net12
rlabel metal1 12558 21964 12558 21964 0 net120
rlabel metal1 27324 19278 27324 19278 0 net121
rlabel metal2 35098 21913 35098 21913 0 net122
rlabel metal1 33856 21862 33856 21862 0 net123
rlabel metal1 1564 24174 1564 24174 0 net124
rlabel metal2 13294 23647 13294 23647 0 net125
rlabel metal2 15042 23800 15042 23800 0 net126
rlabel metal2 14674 21726 14674 21726 0 net127
rlabel metal2 15502 24157 15502 24157 0 net128
rlabel metal2 17250 19244 17250 19244 0 net129
rlabel metal1 2668 6970 2668 6970 0 net13
rlabel metal1 18722 17782 18722 17782 0 net130
rlabel metal1 17296 23698 17296 23698 0 net131
rlabel metal1 20286 22406 20286 22406 0 net132
rlabel metal1 19320 20026 19320 20026 0 net133
rlabel metal1 21988 24174 21988 24174 0 net134
rlabel metal1 4324 10098 4324 10098 0 net135
rlabel via2 16146 20587 16146 20587 0 net136
rlabel metal2 21206 24650 21206 24650 0 net137
rlabel metal2 4784 13940 4784 13940 0 net138
rlabel metal3 6739 12444 6739 12444 0 net139
rlabel metal1 6256 2618 6256 2618 0 net14
rlabel metal1 1564 10642 1564 10642 0 net140
rlabel metal3 6739 10812 6739 10812 0 net141
rlabel metal2 6992 13498 6992 13498 0 net142
rlabel metal1 4784 2414 4784 2414 0 net143
rlabel metal1 7682 2414 7682 2414 0 net144
rlabel metal1 9706 2414 9706 2414 0 net145
rlabel metal1 12420 2414 12420 2414 0 net146
rlabel metal2 15042 3162 15042 3162 0 net147
rlabel metal1 17204 2822 17204 2822 0 net148
rlabel metal1 19136 2822 19136 2822 0 net149
rlabel metal1 4600 21046 4600 21046 0 net15
rlabel metal1 22310 2414 22310 2414 0 net150
rlabel metal1 21850 21522 21850 21522 0 net151
rlabel metal2 23414 20706 23414 20706 0 net152
rlabel metal1 21574 18326 21574 18326 0 net153
rlabel metal2 24978 21879 24978 21879 0 net154
rlabel metal1 23644 21862 23644 21862 0 net155
rlabel metal1 24610 23834 24610 23834 0 net156
rlabel metal2 25990 21760 25990 21760 0 net157
rlabel metal1 26358 19482 26358 19482 0 net158
rlabel metal1 28658 18394 28658 18394 0 net159
rlabel metal1 10534 21658 10534 21658 0 net16
rlabel metal1 16744 20366 16744 20366 0 net160
rlabel metal1 20010 17578 20010 17578 0 net161
rlabel metal1 24150 18802 24150 18802 0 net162
rlabel via1 7590 20417 7590 20417 0 net163
rlabel metal1 19596 16218 19596 16218 0 net164
rlabel metal1 14122 8874 14122 8874 0 net165
rlabel metal1 14168 8466 14168 8466 0 net166
rlabel metal1 10580 6834 10580 6834 0 net167
rlabel metal1 11454 7514 11454 7514 0 net168
rlabel metal2 13570 12002 13570 12002 0 net169
rlabel metal2 5750 16609 5750 16609 0 net17
rlabel metal1 13524 7514 13524 7514 0 net170
rlabel metal1 17020 16626 17020 16626 0 net171
rlabel metal2 15410 17034 15410 17034 0 net172
rlabel metal1 14812 15470 14812 15470 0 net173
rlabel metal1 9568 11866 9568 11866 0 net174
rlabel metal1 9614 9010 9614 9010 0 net175
rlabel metal2 6670 15742 6670 15742 0 net176
rlabel metal1 12098 18190 12098 18190 0 net177
rlabel metal1 20700 14926 20700 14926 0 net178
rlabel metal2 1978 12291 1978 12291 0 net179
rlabel metal1 2070 7378 2070 7378 0 net18
rlabel metal1 4646 9044 4646 9044 0 net180
rlabel metal2 12558 8704 12558 8704 0 net181
rlabel metal2 5842 9673 5842 9673 0 net182
rlabel metal1 33856 20978 33856 20978 0 net183
rlabel metal1 10258 21488 10258 21488 0 net184
rlabel metal2 9982 16847 9982 16847 0 net185
rlabel metal1 13800 17170 13800 17170 0 net186
rlabel metal2 12834 16082 12834 16082 0 net187
rlabel metal1 16100 12750 16100 12750 0 net188
rlabel metal1 16146 8602 16146 8602 0 net189
rlabel metal1 2208 7854 2208 7854 0 net19
rlabel metal1 7452 10778 7452 10778 0 net190
rlabel metal1 5750 10030 5750 10030 0 net191
rlabel metal2 16514 14756 16514 14756 0 net192
rlabel metal1 12650 12920 12650 12920 0 net193
rlabel metal1 27968 16558 27968 16558 0 net194
rlabel via2 35650 23035 35650 23035 0 net195
rlabel metal2 36294 21709 36294 21709 0 net196
rlabel metal1 18676 16422 18676 16422 0 net197
rlabel metal2 17526 19856 17526 19856 0 net198
rlabel metal1 43884 23086 43884 23086 0 net199
rlabel metal2 48438 22576 48438 22576 0 net2
rlabel metal1 1886 8364 1886 8364 0 net20
rlabel metal1 42734 22984 42734 22984 0 net200
rlabel metal1 43746 23664 43746 23664 0 net201
rlabel metal1 44114 23290 44114 23290 0 net202
rlabel metal2 43286 22916 43286 22916 0 net203
rlabel metal1 1656 24038 1656 24038 0 net204
rlabel metal1 41446 23732 41446 23732 0 net205
rlabel metal2 48714 23868 48714 23868 0 net206
rlabel metal1 41354 22542 41354 22542 0 net207
rlabel metal1 3128 3026 3128 3026 0 net208
rlabel metal1 8142 2958 8142 2958 0 net209
rlabel metal1 6578 16626 6578 16626 0 net21
rlabel metal1 28658 2618 28658 2618 0 net210
rlabel metal2 37490 3774 37490 3774 0 net211
rlabel metal1 33994 2618 33994 2618 0 net212
rlabel metal1 35282 3060 35282 3060 0 net213
rlabel metal1 25990 3026 25990 3026 0 net214
rlabel metal1 36869 3502 36869 3502 0 net215
rlabel metal1 31326 2618 31326 2618 0 net216
rlabel metal2 35742 4556 35742 4556 0 net217
rlabel metal1 34362 23766 34362 23766 0 net218
rlabel metal1 33028 21522 33028 21522 0 net219
rlabel metal1 2024 9486 2024 9486 0 net22
rlabel metal1 1840 8942 1840 8942 0 net220
rlabel metal2 36018 23902 36018 23902 0 net221
rlabel metal1 3450 6732 3450 6732 0 net222
rlabel metal2 33534 23902 33534 23902 0 net223
rlabel metal1 35236 23086 35236 23086 0 net224
rlabel metal2 41446 23324 41446 23324 0 net225
rlabel metal1 34132 23086 34132 23086 0 net226
rlabel metal2 38502 23902 38502 23902 0 net227
rlabel metal1 40342 23154 40342 23154 0 net228
rlabel metal1 39974 23766 39974 23766 0 net229
rlabel metal1 2300 8942 2300 8942 0 net23
rlabel metal2 2806 9996 2806 9996 0 net230
rlabel metal1 30728 24242 30728 24242 0 net231
rlabel metal2 30682 23902 30682 23902 0 net232
rlabel metal1 1932 11866 1932 11866 0 net233
rlabel metal1 48990 23290 48990 23290 0 net234
rlabel metal1 48668 21998 48668 21998 0 net235
rlabel metal2 46874 22780 46874 22780 0 net236
rlabel metal1 2760 4114 2760 4114 0 net237
rlabel metal1 3864 3026 3864 3026 0 net238
rlabel metal1 5934 3026 5934 3026 0 net239
rlabel metal2 19734 16422 19734 16422 0 net24
rlabel metal1 3933 2278 3933 2278 0 net25
rlabel metal2 15410 9605 15410 9605 0 net26
rlabel metal1 1288 3502 1288 3502 0 net27
rlabel metal2 14766 8058 14766 8058 0 net28
rlabel metal1 7314 3706 7314 3706 0 net29
rlabel metal2 13478 5746 13478 5746 0 net3
rlabel metal1 6900 3978 6900 3978 0 net30
rlabel metal1 10672 15334 10672 15334 0 net31
rlabel metal1 8970 14246 8970 14246 0 net32
rlabel via2 13938 20757 13938 20757 0 net33
rlabel metal1 32936 21318 32936 21318 0 net34
rlabel metal1 4554 21862 4554 21862 0 net35
rlabel metal2 9890 17119 9890 17119 0 net36
rlabel metal2 30866 21624 30866 21624 0 net37
rlabel metal2 35650 21760 35650 21760 0 net38
rlabel metal1 35742 23834 35742 23834 0 net39
rlabel via2 6394 13821 6394 13821 0 net4
rlabel metal2 31050 23154 31050 23154 0 net40
rlabel metal2 33718 24225 33718 24225 0 net41
rlabel metal1 15318 18054 15318 18054 0 net42
rlabel metal1 34362 23018 34362 23018 0 net43
rlabel metal1 17480 20978 17480 20978 0 net44
rlabel metal2 36202 24361 36202 24361 0 net45
rlabel metal1 31878 21930 31878 21930 0 net46
rlabel metal1 32338 21488 32338 21488 0 net47
rlabel metal2 37490 21182 37490 21182 0 net48
rlabel metal2 37582 19720 37582 19720 0 net49
rlabel metal1 1886 6324 1886 6324 0 net5
rlabel via2 16974 16133 16974 16133 0 net50
rlabel metal1 14398 18802 14398 18802 0 net51
rlabel metal2 36478 21199 36478 21199 0 net52
rlabel metal2 40710 21641 40710 21641 0 net53
rlabel metal2 41354 21114 41354 21114 0 net54
rlabel metal1 8142 24038 8142 24038 0 net55
rlabel metal2 14306 20077 14306 20077 0 net56
rlabel metal2 14306 24089 14306 24089 0 net57
rlabel metal1 27048 24174 27048 24174 0 net58
rlabel metal1 29394 22984 29394 22984 0 net59
rlabel metal1 6118 5814 6118 5814 0 net6
rlabel metal1 26680 23086 26680 23086 0 net60
rlabel metal1 26082 22746 26082 22746 0 net61
rlabel metal1 14490 21998 14490 21998 0 net62
rlabel metal2 25530 4352 25530 4352 0 net63
rlabel metal1 27876 3162 27876 3162 0 net64
rlabel metal1 30590 2890 30590 2890 0 net65
rlabel metal2 29670 4148 29670 4148 0 net66
rlabel metal1 33994 2482 33994 2482 0 net67
rlabel metal1 42734 22610 42734 22610 0 net68
rlabel metal2 45402 21437 45402 21437 0 net69
rlabel metal1 4462 6902 4462 6902 0 net7
rlabel metal2 43378 21216 43378 21216 0 net70
rlabel metal2 43470 21845 43470 21845 0 net71
rlabel metal2 46966 21216 46966 21216 0 net72
rlabel metal2 44942 23936 44942 23936 0 net73
rlabel metal1 46874 20774 46874 20774 0 net74
rlabel metal2 45034 20842 45034 20842 0 net75
rlabel metal2 45770 21097 45770 21097 0 net76
rlabel metal1 35880 19992 35880 19992 0 net77
rlabel metal2 42826 19584 42826 19584 0 net78
rlabel metal2 43470 17000 43470 17000 0 net79
rlabel metal3 3841 9452 3841 9452 0 net8
rlabel metal1 47932 23834 47932 23834 0 net80
rlabel metal1 47794 21522 47794 21522 0 net81
rlabel metal2 5934 20026 5934 20026 0 net82
rlabel via2 1794 13277 1794 13277 0 net83
rlabel metal2 15134 18819 15134 18819 0 net84
rlabel metal1 5704 19278 5704 19278 0 net85
rlabel metal2 4278 19873 4278 19873 0 net86
rlabel metal2 1794 21964 1794 21964 0 net87
rlabel metal1 1840 20910 1840 20910 0 net88
rlabel metal1 1610 21556 1610 21556 0 net89
rlabel metal2 13386 14790 13386 14790 0 net9
rlabel metal1 1426 20366 1426 20366 0 net90
rlabel metal1 2277 21998 2277 21998 0 net91
rlabel metal1 1794 22644 1794 22644 0 net92
rlabel metal1 2277 23086 2277 23086 0 net93
rlabel via2 1794 13923 1794 13923 0 net94
rlabel metal1 4140 21998 4140 21998 0 net95
rlabel metal1 4278 19346 4278 19346 0 net96
rlabel metal2 6118 21148 6118 21148 0 net97
rlabel metal1 6440 19346 6440 19346 0 net98
rlabel metal1 6026 12682 6026 12682 0 net99
rlabel metal2 38778 3458 38778 3458 0 prog_clk
rlabel metal1 41998 24378 41998 24378 0 prog_reset
rlabel metal1 18722 16966 18722 16966 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal1 25760 19890 25760 19890 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal2 29026 18224 29026 18224 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 16560 20434 16560 20434 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal1 17250 23018 17250 23018 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal2 17158 24378 17158 24378 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 16744 21454 16744 21454 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel metal1 19044 23630 19044 23630 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 15134 21012 15134 21012 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel metal1 20930 22746 20930 22746 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel metal2 16422 21590 16422 21590 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal2 23782 23358 23782 23358 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 23920 21454 23920 21454 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal1 23828 21590 23828 21590 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal1 26358 18938 26358 18938 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal1 26680 20366 26680 20366 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 18676 19890 18676 19890 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 20601 19142 20601 19142 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal2 26082 21658 26082 21658 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal1 27738 20026 27738 20026 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel via2 26634 23477 26634 23477 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal1 26910 22202 26910 22202 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal2 29026 23936 29026 23936 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal2 28934 23324 28934 23324 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal1 28152 21590 28152 21590 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel metal1 31142 23154 31142 23154 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 28372 19142 28372 19142 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal2 30222 20842 30222 20842 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel metal1 30084 18802 30084 18802 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal1 29348 19142 29348 19142 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal1 20102 19890 20102 19890 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel metal2 19734 21148 19734 21148 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 28842 17408 28842 17408 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal2 20654 19822 20654 19822 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal1 21804 19890 21804 19890 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 19090 20434 19090 20434 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal1 25070 15062 25070 15062 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal2 39606 20264 39606 20264 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 24978 16014 24978 16014 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 20654 13804 20654 13804 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal1 17250 9962 17250 9962 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal2 24058 14926 24058 14926 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 21436 12750 21436 12750 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 16284 8874 16284 8874 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal1 20470 14450 20470 14450 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 15548 10098 15548 10098 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel metal2 14766 9010 14766 9010 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 13202 12716 13202 12716 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal1 14628 11186 14628 11186 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 17480 13838 17480 13838 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal1 17250 13226 17250 13226 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 21206 9690 21206 9690 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 25162 14416 25162 14416 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 19504 9962 19504 9962 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 18124 15334 18124 15334 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal2 17342 14722 17342 14722 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal2 16330 14620 16330 14620 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal1 14904 15062 14904 15062 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 15548 13498 15548 13498 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal1 15502 13362 15502 13362 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal2 11822 10200 11822 10200 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal1 13110 11798 13110 11798 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 13432 9418 13432 9418 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal2 12006 9860 12006 9860 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12650 14178 12650 14178 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal1 12328 13226 12328 13226 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 12558 18156 12558 18156 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal2 13570 15470 13570 15470 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 10994 19822 10994 19822 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal1 13708 17782 13708 17782 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 9982 20026 9982 20026 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal2 11178 19941 11178 19941 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 4968 18666 4968 18666 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal1 7866 15980 7866 15980 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal1 19908 13498 19908 13498 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal2 22862 15232 22862 15232 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 17388 11050 17388 11050 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 7130 21590 7130 21590 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel metal1 7406 18598 7406 18598 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 8096 20978 8096 20978 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel metal1 9430 21624 9430 21624 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 13432 21590 13432 21590 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel metal1 17710 19278 17710 19278 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 15180 19890 15180 19890 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal1 14950 19346 14950 19346 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 16790 17714 16790 17714 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal2 20102 18428 20102 18428 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 18400 17238 18400 17238 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 21942 14824 21942 14824 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal1 21390 17068 21390 17068 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 19274 13226 19274 13226 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 23874 14518 23874 14518 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 20378 10268 20378 10268 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 3634 14994 3634 14994 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 26450 19686 26450 19686 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27278 16422 27278 16422 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21022 18768 21022 18768 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 4324 12886 4324 12886 0 sb_8__0_.mux_left_track_11.out
rlabel metal2 23966 23970 23966 23970 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 2231 11322 2231 11322 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 10212 17136 10212 17136 0 sb_8__0_.mux_left_track_13.out
rlabel metal2 16054 22559 16054 22559 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 15594 21403 15594 21403 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 17020 19992 17020 19992 0 sb_8__0_.mux_left_track_15.out
rlabel via2 17894 20859 17894 20859 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15594 21114 15594 21114 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 5612 14212 5612 14212 0 sb_8__0_.mux_left_track_17.out
rlabel metal2 16238 21318 16238 21318 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 15847 20740 15847 20740 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5520 17170 5520 17170 0 sb_8__0_.mux_left_track_19.out
rlabel metal2 22494 22015 22494 22015 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19918 15470 19918 15470 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7866 14994 7866 14994 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 27140 20570 27140 20570 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22126 13192 22126 13192 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32062 18139 32062 18139 0 sb_8__0_.mux_left_track_3.out
rlabel metal1 18032 19822 18032 19822 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 17250 19941 17250 19941 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16146 17442 16146 17442 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 26496 21318 26496 21318 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17158 17510 17158 17510 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1196 6834 1196 6834 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 24932 22202 24932 22202 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 23322 21845 23322 21845 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 9292 13668 9292 13668 0 sb_8__0_.mux_left_track_35.out
rlabel metal2 30590 23596 30590 23596 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12834 9435 12834 9435 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21298 16439 21298 16439 0 sb_8__0_.mux_left_track_45.out
rlabel metal1 26312 21522 26312 21522 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25438 21318 25438 21318 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9614 16201 9614 16201 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 26450 20774 26450 20774 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13754 15589 13754 15589 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13846 14977 13846 14977 0 sb_8__0_.mux_left_track_49.out
rlabel metal1 30406 18734 30406 18734 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17618 16524 17618 16524 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16836 21862 16836 21862 0 sb_8__0_.mux_left_track_5.out
rlabel metal1 17250 20570 17250 20570 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16790 19482 16790 19482 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14030 14280 14030 14280 0 sb_8__0_.mux_left_track_51.out
rlabel metal2 21206 17136 21206 17136 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16376 16082 16376 16082 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6992 16422 6992 16422 0 sb_8__0_.mux_left_track_7.out
rlabel metal1 22586 19414 22586 19414 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 19482 22862 19482 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14858 18734 14858 18734 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11592 17170 11592 17170 0 sb_8__0_.mux_left_track_9.out
rlabel metal1 18538 20536 18538 20536 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12512 17340 12512 17340 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16376 16762 16376 16762 0 sb_8__0_.mux_top_track_0.out
rlabel metal2 27094 17408 27094 17408 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27738 16490 27738 16490 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26634 16456 26634 16456 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23782 19414 23782 19414 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23598 18938 23598 18938 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18906 16082 18906 16082 0 sb_8__0_.mux_top_track_10.out
rlabel metal1 21643 12818 21643 12818 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21160 12954 21160 12954 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20102 12614 20102 12614 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15134 9146 15134 9146 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17388 11594 17388 11594 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 14398 16473 14398 16473 0 sb_8__0_.mux_top_track_12.out
rlabel metal1 16054 10540 16054 10540 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14628 8602 14628 8602 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15364 14212 15364 14212 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15640 16966 15640 16966 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 15916 10710 15916 10710 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 9588 12466 9588 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15042 10506 15042 10506 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 10994 15963 10994 15963 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 18032 11866 18032 11866 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12673 12818 12673 12818 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11776 12954 11776 12954 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21712 16014 21712 16014 0 sb_8__0_.mux_top_track_18.out
rlabel metal1 19228 16150 19228 16150 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13754 14042 13754 14042 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16974 15946 16974 15946 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19090 19652 19090 19652 0 sb_8__0_.mux_top_track_2.out
rlabel metal1 24840 13974 24840 13974 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25392 14042 25392 14042 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22080 9622 22080 9622 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13524 8058 13524 8058 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19182 19346 19182 19346 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 34040 21998 34040 21998 0 sb_8__0_.mux_top_track_20.out
rlabel metal2 15870 16388 15870 16388 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 14824 12926 14824 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34960 21318 34960 21318 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 14444 14042 14444 14042 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19044 14382 19044 14382 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 9430 13379 9430 13379 0 sb_8__0_.mux_top_track_24.out
rlabel metal2 13754 14144 13754 14144 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14214 14246 14214 14246 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 33074 21420 33074 21420 0 sb_8__0_.mux_top_track_26.out
rlabel metal2 10626 11934 10626 11934 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 3404 13940 3404 13940 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32522 14416 32522 14416 0 sb_8__0_.mux_top_track_28.out
rlabel metal1 10442 10234 10442 10234 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10856 8942 10856 8942 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 29762 20570 29762 20570 0 sb_8__0_.mux_top_track_30.out
rlabel metal2 12558 13872 12558 13872 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 12098 15589 12098 15589 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34132 21046 34132 21046 0 sb_8__0_.mux_top_track_32.out
rlabel metal1 12880 15130 12880 15130 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32430 20910 32430 20910 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35190 22610 35190 22610 0 sb_8__0_.mux_top_track_34.out
rlabel metal2 11638 18326 11638 18326 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11914 19431 11914 19431 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2300 10234 2300 10234 0 sb_8__0_.mux_top_track_36.out
rlabel metal1 11362 18938 11362 18938 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 2162 11866 2162 11866 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4784 9146 4784 9146 0 sb_8__0_.mux_top_track_38.out
rlabel metal1 7268 16218 7268 16218 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 5451 9588 5451 9588 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 16422 18308 16422 0 sb_8__0_.mux_top_track_4.out
rlabel metal1 21114 12852 21114 12852 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18630 12954 18630 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16928 12954 16928 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15778 13906 15778 13906 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16422 14042 16422 14042 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5566 8330 5566 8330 0 sb_8__0_.mux_top_track_40.out
rlabel metal1 7728 17306 7728 17306 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 1012 16762 1012 16762 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9154 8194 9154 8194 0 sb_8__0_.mux_top_track_42.out
rlabel metal1 8694 20910 8694 20910 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8924 18836 8924 18836 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2116 10574 2116 10574 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 17894 19448 17894 19448 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11730 19822 11730 19822 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32430 21471 32430 21471 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 32775 20740 32775 20740 0 sb_8__0_.mux_top_track_46.out
rlabel metal1 18078 18598 18078 18598 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12742 18904 12742 18904 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32614 21488 32614 21488 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 2622 10115 2622 10115 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 17526 18122 17526 18122 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13754 17850 13754 17850 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 15042 18139 15042 18139 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19596 13770 19596 13770 0 sb_8__0_.mux_top_track_50.out
rlabel metal1 19044 18394 19044 18394 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13662 16422 13662 16422 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19642 13872 19642 13872 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 34270 22899 34270 22899 0 sb_8__0_.mux_top_track_6.out
rlabel metal2 20746 16796 20746 16796 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 16558 22862 16558 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20470 15062 20470 15062 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19826 14994 19826 14994 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19780 14858 19780 14858 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18262 17714 18262 17714 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 23322 13396 23322 13396 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23276 13226 23276 13226 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21666 13668 21666 13668 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18032 8330 18032 8330 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19550 14042 19550 14042 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 44758 25340 44758 25340 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 45494 25296 45494 25296 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46368 24174 46368 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 46736 23698 46736 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47564 24174 47564 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 47932 23086 47932 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44344 23698 44344 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal2 44114 25034 44114 25034 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel via2 49082 21981 49082 21981 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 49082 22763 49082 22763 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 48346 22831 48346 22831 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 48162 23698 48162 23698 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 36478 2924 36478 2924 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 36938 3400 36938 3400 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 38594 3060 38594 3060 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 39054 3536 39054 3536 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
