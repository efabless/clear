VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2544.940 BY 2903.800 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 367.340 29.180 367.940 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 170.140 29.180 170.740 ;
    END
  END Test_en
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 4.500 2903.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 2544.940 4.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2899.300 2544.940 2903.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2540.440 0.000 2544.940 2903.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 140.950 2544.940 145.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 185.950 2544.940 190.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 230.950 2544.940 235.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 275.950 2544.940 280.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 320.950 2544.940 325.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 365.950 2544.940 370.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 410.950 2544.940 415.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 455.950 2544.940 460.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 500.950 2544.940 505.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 545.950 2544.940 550.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 590.950 2544.940 595.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 635.950 2544.940 640.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 680.950 2544.940 685.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 725.950 2544.940 730.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 770.950 2544.940 775.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 815.950 2544.940 820.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 860.950 2544.940 865.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 905.950 2544.940 910.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 950.950 2544.940 955.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 995.950 2544.940 1000.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1040.950 2544.940 1045.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1085.950 2544.940 1090.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1130.950 2544.940 1135.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1175.950 2544.940 1180.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1220.950 2544.940 1225.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1265.950 2544.940 1270.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1310.950 2544.940 1315.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1355.950 2544.940 1360.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1400.950 2544.940 1405.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1445.950 2544.940 1450.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1490.950 2544.940 1495.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1535.950 2544.940 1540.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1580.950 2544.940 1585.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1625.950 2544.940 1630.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1670.950 2544.940 1675.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1715.950 2544.940 1720.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1760.950 2544.940 1765.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1805.950 2544.940 1810.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1850.950 2544.940 1855.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1895.950 2544.940 1900.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1940.950 2544.940 1945.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1985.950 2544.940 1990.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2030.950 2544.940 2035.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2075.950 2544.940 2080.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2120.950 2544.940 2125.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2165.950 2544.940 2170.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2210.950 2544.940 2215.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2255.950 2544.940 2260.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2300.950 2544.940 2305.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2345.950 2544.940 2350.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2390.950 2544.940 2395.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2435.950 2544.940 2440.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2480.950 2544.940 2485.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2525.950 2544.940 2530.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2570.950 2544.940 2575.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2615.950 2544.940 2620.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2660.950 2544.940 2665.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2705.950 2544.940 2710.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2750.950 2544.940 2755.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2795.950 2544.940 2800.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2840.950 2544.940 2845.450 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.200 6.200 10.700 2897.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 6.200 6.200 2538.740 10.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 6.200 2893.100 2538.740 2897.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2534.240 6.200 2538.740 2897.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 118.450 2544.940 122.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 163.450 2544.940 167.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 208.450 2544.940 212.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 253.450 2544.940 257.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 298.450 2544.940 302.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 343.450 2544.940 347.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 388.450 2544.940 392.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 433.450 2544.940 437.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 478.450 2544.940 482.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 523.450 2544.940 527.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 568.450 2544.940 572.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 613.450 2544.940 617.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 658.450 2544.940 662.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 703.450 2544.940 707.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 748.450 2544.940 752.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 793.450 2544.940 797.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 838.450 2544.940 842.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 883.450 2544.940 887.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 928.450 2544.940 932.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 973.450 2544.940 977.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1018.450 2544.940 1022.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1063.450 2544.940 1067.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1108.450 2544.940 1112.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1153.450 2544.940 1157.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1198.450 2544.940 1202.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1243.450 2544.940 1247.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1288.450 2544.940 1292.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1333.450 2544.940 1337.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1378.450 2544.940 1382.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1423.450 2544.940 1427.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1468.450 2544.940 1472.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1513.450 2544.940 1517.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1558.450 2544.940 1562.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1603.450 2544.940 1607.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1648.450 2544.940 1652.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1693.450 2544.940 1697.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1738.450 2544.940 1742.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1783.450 2544.940 1787.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1828.450 2544.940 1832.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1873.450 2544.940 1877.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1918.450 2544.940 1922.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 1963.450 2544.940 1967.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2008.450 2544.940 2012.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2053.450 2544.940 2057.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2098.450 2544.940 2102.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2143.450 2544.940 2147.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2188.450 2544.940 2192.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2233.450 2544.940 2237.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2278.450 2544.940 2282.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2323.450 2544.940 2327.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2368.450 2544.940 2372.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2413.450 2544.940 2417.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2458.450 2544.940 2462.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2503.450 2544.940 2507.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2548.450 2544.940 2552.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2593.450 2544.940 2597.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2638.450 2544.940 2642.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2683.450 2544.940 2687.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2728.450 2544.940 2732.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2773.450 2544.940 2777.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2818.450 2544.940 2822.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2863.450 2544.940 2867.950 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 2701.100 2520.180 2701.700 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 71.540 29.180 72.140 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 268.740 29.180 269.340 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.330 2880.820 76.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 559.100 2520.180 559.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 916.100 2520.180 916.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1273.100 2520.180 1273.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1630.100 2520.180 1630.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1987.100 2520.180 1987.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 2344.100 2520.180 2344.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.810 19.820 2210.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.310 19.820 2221.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.810 19.820 2233.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.310 19.820 2244.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.330 2880.820 168.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2255.810 19.820 2256.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2267.310 19.820 2267.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.810 19.820 2279.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.310 19.820 2290.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.810 19.820 2302.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.310 19.820 1899.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.810 19.820 1911.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.310 19.820 1922.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.810 19.820 1934.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.310 19.820 1945.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.330 2880.820 260.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.810 19.820 1957.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.310 19.820 1968.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.810 19.820 1980.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.310 19.820 1991.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.810 19.820 1589.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.310 19.820 1600.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.810 19.820 1612.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.310 19.820 1623.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.810 19.820 1635.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.310 19.820 1646.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.330 2880.820 352.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.810 19.820 1658.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.310 19.820 1669.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.810 19.820 1681.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.310 19.820 1278.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.810 19.820 1290.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.310 19.820 1301.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.810 19.820 1313.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.310 19.820 1324.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.810 19.820 1336.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.310 19.820 1347.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.330 2880.820 444.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.810 19.820 1359.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.310 19.820 1370.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.810 19.820 968.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.310 19.820 979.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.810 19.820 991.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.310 19.820 1002.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.810 19.820 1014.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.310 19.820 1025.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.810 19.820 1037.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.310 19.820 1048.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.330 2880.820 536.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.810 19.820 1060.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.310 19.820 657.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.810 19.820 669.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.310 19.820 680.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.810 19.820 692.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.310 19.820 703.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.810 19.820 715.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.310 19.820 726.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.810 19.820 738.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.310 19.820 749.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.330 2880.820 628.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.810 19.820 347.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.310 19.820 358.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.810 19.820 370.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.310 19.820 381.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.810 19.820 393.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.310 19.820 404.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.810 19.820 416.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.310 19.820 427.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.810 19.820 439.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.310 19.820 36.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.330 2880.820 720.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.810 19.820 48.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.310 19.820 59.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.810 19.820 71.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.310 19.820 82.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.810 19.820 94.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.310 19.820 105.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.810 19.820 117.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.310 19.820 128.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 465.940 29.180 466.540 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 761.740 29.180 762.340 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.330 2880.820 812.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1057.540 29.180 1058.140 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1353.340 29.180 1353.940 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1649.140 29.180 1649.740 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1944.940 29.180 1945.540 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2240.740 29.180 2241.340 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2536.540 29.180 2537.140 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 202.100 2520.180 202.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.330 2880.820 904.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 678.100 2520.180 678.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1035.100 2520.180 1035.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1392.100 2520.180 1392.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1749.100 2520.180 1749.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 2106.100 2520.180 2106.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 2463.100 2520.180 2463.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.310 19.820 2313.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.810 19.820 2325.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2336.310 19.820 2336.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2347.810 19.820 2348.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.330 2880.820 996.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.310 19.820 2359.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.810 19.820 2371.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.310 19.820 2382.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.810 19.820 2394.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.310 19.820 2405.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.810 19.820 2003.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.310 19.820 2014.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.810 19.820 2026.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2037.310 19.820 2037.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.810 19.820 2049.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.330 2880.820 1088.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.310 19.820 2060.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.810 19.820 2072.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.310 19.820 2083.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.810 19.820 2095.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.310 19.820 1692.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.810 19.820 1704.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.310 19.820 1715.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.810 19.820 1727.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.310 19.820 1738.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.810 19.820 1750.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.330 2880.820 1180.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.310 19.820 1761.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.810 19.820 1773.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.310 19.820 1784.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.810 19.820 1382.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.310 19.820 1393.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.810 19.820 1405.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.310 19.820 1416.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.810 19.820 1428.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.310 19.820 1439.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.810 19.820 1451.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.330 2880.820 1272.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.310 19.820 1462.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.810 19.820 1474.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.310 19.820 1071.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.810 19.820 1083.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.310 19.820 1094.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.810 19.820 1106.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.310 19.820 1117.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.810 19.820 1129.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.310 19.820 1140.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.810 19.820 1152.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.330 2880.820 1364.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.310 19.820 1163.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.810 19.820 761.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.310 19.820 772.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.810 19.820 784.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.310 19.820 795.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.810 19.820 807.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.310 19.820 818.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.810 19.820 830.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.310 19.820 841.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.810 19.820 853.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.330 2880.820 1456.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.310 19.820 450.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.810 19.820 462.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.310 19.820 473.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.810 19.820 485.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.310 19.820 496.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.810 19.820 508.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.310 19.820 519.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.810 19.820 531.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.310 19.820 542.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.810 19.820 140.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.330 2880.820 1548.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.310 19.820 151.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.810 19.820 163.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.310 19.820 174.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.810 19.820 186.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.310 19.820 197.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.810 19.820 209.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.310 19.820 220.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.810 19.820 232.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 564.540 29.180 565.140 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 860.340 29.180 860.940 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.330 2880.820 1640.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1156.140 29.180 1156.740 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1451.940 29.180 1452.540 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1747.740 29.180 1748.340 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2043.540 29.180 2044.140 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2339.340 29.180 2339.940 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2635.140 29.180 2635.740 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 321.100 2520.180 321.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.330 2880.820 1732.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 797.100 2520.180 797.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1154.100 2520.180 1154.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1511.100 2520.180 1511.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 1868.100 2520.180 1868.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 2225.100 2520.180 2225.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 2582.100 2520.180 2582.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.810 19.820 2417.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.310 19.820 2428.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.810 19.820 2440.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2451.310 19.820 2451.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.330 2880.820 1824.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2462.810 19.820 2463.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2474.310 19.820 2474.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.810 19.820 2486.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2497.310 19.820 2497.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.810 19.820 2509.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.310 19.820 2106.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.810 19.820 2118.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.310 19.820 2129.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.810 19.820 2141.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.310 19.820 2152.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.330 2880.820 1916.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.810 19.820 2164.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.310 19.820 2175.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.810 19.820 2187.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.310 19.820 2198.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.810 19.820 1796.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.310 19.820 1807.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.810 19.820 1819.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.310 19.820 1830.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.810 19.820 1842.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.310 19.820 1853.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.330 2880.820 2008.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.810 19.820 1865.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.310 19.820 1876.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.810 19.820 1888.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.310 19.820 1485.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.810 19.820 1497.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.310 19.820 1508.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.810 19.820 1520.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.310 19.820 1531.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.810 19.820 1543.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.310 19.820 1554.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.330 2880.820 2100.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.810 19.820 1566.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.310 19.820 1577.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.810 19.820 1175.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.310 19.820 1186.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.810 19.820 1198.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.310 19.820 1209.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.810 19.820 1221.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.310 19.820 1232.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.810 19.820 1244.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.310 19.820 1255.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.330 2880.820 2192.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.810 19.820 1267.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.310 19.820 864.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.810 19.820 876.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.310 19.820 887.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.810 19.820 899.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.310 19.820 910.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.810 19.820 922.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.310 19.820 933.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.810 19.820 945.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.310 19.820 956.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.330 2880.820 2284.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.810 19.820 554.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.310 19.820 565.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.810 19.820 577.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.310 19.820 588.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.810 19.820 600.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.310 19.820 611.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.810 19.820 623.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.310 19.820 634.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.810 19.820 646.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.310 19.820 243.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.330 2880.820 2376.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.810 19.820 255.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.310 19.820 266.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.810 19.820 278.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.310 19.820 289.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.810 19.820 301.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.310 19.820 312.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.810 19.820 324.090 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.310 19.820 335.590 23.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 663.140 29.180 663.740 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 958.940 29.180 959.540 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2468.330 2880.820 2468.610 2884.820 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1254.740 29.180 1255.340 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1550.540 29.180 1551.140 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 1846.340 29.180 1846.940 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2142.140 29.180 2142.740 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2437.940 29.180 2438.540 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2733.740 29.180 2734.340 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 440.100 2520.180 440.700 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 83.100 2520.180 83.700 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.180 2832.340 29.180 2832.940 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.180 2820.100 2520.180 2820.700 ;
    END
  END sc_tail
  OBS
      LAYER li1 ;
        RECT 80.700 105.615 2464.660 2870.025 ;
      LAYER met1 ;
        RECT 36.290 25.980 2509.110 2870.180 ;
      LAYER met2 ;
        RECT 36.320 2880.540 76.050 2880.990 ;
        RECT 76.890 2880.540 168.050 2880.990 ;
        RECT 168.890 2880.540 260.050 2880.990 ;
        RECT 260.890 2880.540 352.050 2880.990 ;
        RECT 352.890 2880.540 444.050 2880.990 ;
        RECT 444.890 2880.540 536.050 2880.990 ;
        RECT 536.890 2880.540 628.050 2880.990 ;
        RECT 628.890 2880.540 720.050 2880.990 ;
        RECT 720.890 2880.540 812.050 2880.990 ;
        RECT 812.890 2880.540 904.050 2880.990 ;
        RECT 904.890 2880.540 996.050 2880.990 ;
        RECT 996.890 2880.540 1088.050 2880.990 ;
        RECT 1088.890 2880.540 1180.050 2880.990 ;
        RECT 1180.890 2880.540 1272.050 2880.990 ;
        RECT 1272.890 2880.540 1364.050 2880.990 ;
        RECT 1364.890 2880.540 1456.050 2880.990 ;
        RECT 1456.890 2880.540 1548.050 2880.990 ;
        RECT 1548.890 2880.540 1640.050 2880.990 ;
        RECT 1640.890 2880.540 1732.050 2880.990 ;
        RECT 1732.890 2880.540 1824.050 2880.990 ;
        RECT 1824.890 2880.540 1916.050 2880.990 ;
        RECT 1916.890 2880.540 2008.050 2880.990 ;
        RECT 2008.890 2880.540 2100.050 2880.990 ;
        RECT 2100.890 2880.540 2192.050 2880.990 ;
        RECT 2192.890 2880.540 2284.050 2880.990 ;
        RECT 2284.890 2880.540 2376.050 2880.990 ;
        RECT 2376.890 2880.540 2468.050 2880.990 ;
        RECT 2468.890 2880.540 2509.080 2880.990 ;
        RECT 36.320 24.100 2509.080 2880.540 ;
        RECT 36.870 23.490 47.530 24.100 ;
        RECT 48.370 23.490 59.030 24.100 ;
        RECT 59.870 23.490 70.530 24.100 ;
        RECT 71.370 23.490 82.030 24.100 ;
        RECT 82.870 23.490 93.530 24.100 ;
        RECT 94.370 23.490 105.030 24.100 ;
        RECT 105.870 23.490 116.530 24.100 ;
        RECT 117.370 23.490 128.030 24.100 ;
        RECT 128.870 23.490 139.530 24.100 ;
        RECT 140.370 23.490 151.030 24.100 ;
        RECT 151.870 23.490 162.530 24.100 ;
        RECT 163.370 23.490 174.030 24.100 ;
        RECT 174.870 23.490 185.530 24.100 ;
        RECT 186.370 23.490 197.030 24.100 ;
        RECT 197.870 23.490 208.530 24.100 ;
        RECT 209.370 23.490 220.030 24.100 ;
        RECT 220.870 23.490 231.530 24.100 ;
        RECT 232.370 23.490 243.030 24.100 ;
        RECT 243.870 23.490 254.530 24.100 ;
        RECT 255.370 23.490 266.030 24.100 ;
        RECT 266.870 23.490 277.530 24.100 ;
        RECT 278.370 23.490 289.030 24.100 ;
        RECT 289.870 23.490 300.530 24.100 ;
        RECT 301.370 23.490 312.030 24.100 ;
        RECT 312.870 23.490 323.530 24.100 ;
        RECT 324.370 23.490 335.030 24.100 ;
        RECT 335.870 23.490 346.530 24.100 ;
        RECT 347.370 23.490 358.030 24.100 ;
        RECT 358.870 23.490 369.530 24.100 ;
        RECT 370.370 23.490 381.030 24.100 ;
        RECT 381.870 23.490 392.530 24.100 ;
        RECT 393.370 23.490 404.030 24.100 ;
        RECT 404.870 23.490 415.530 24.100 ;
        RECT 416.370 23.490 427.030 24.100 ;
        RECT 427.870 23.490 438.530 24.100 ;
        RECT 439.370 23.490 450.030 24.100 ;
        RECT 450.870 23.490 461.530 24.100 ;
        RECT 462.370 23.490 473.030 24.100 ;
        RECT 473.870 23.490 484.530 24.100 ;
        RECT 485.370 23.490 496.030 24.100 ;
        RECT 496.870 23.490 507.530 24.100 ;
        RECT 508.370 23.490 519.030 24.100 ;
        RECT 519.870 23.490 530.530 24.100 ;
        RECT 531.370 23.490 542.030 24.100 ;
        RECT 542.870 23.490 553.530 24.100 ;
        RECT 554.370 23.490 565.030 24.100 ;
        RECT 565.870 23.490 576.530 24.100 ;
        RECT 577.370 23.490 588.030 24.100 ;
        RECT 588.870 23.490 599.530 24.100 ;
        RECT 600.370 23.490 611.030 24.100 ;
        RECT 611.870 23.490 622.530 24.100 ;
        RECT 623.370 23.490 634.030 24.100 ;
        RECT 634.870 23.490 645.530 24.100 ;
        RECT 646.370 23.490 657.030 24.100 ;
        RECT 657.870 23.490 668.530 24.100 ;
        RECT 669.370 23.490 680.030 24.100 ;
        RECT 680.870 23.490 691.530 24.100 ;
        RECT 692.370 23.490 703.030 24.100 ;
        RECT 703.870 23.490 714.530 24.100 ;
        RECT 715.370 23.490 726.030 24.100 ;
        RECT 726.870 23.490 737.530 24.100 ;
        RECT 738.370 23.490 749.030 24.100 ;
        RECT 749.870 23.490 760.530 24.100 ;
        RECT 761.370 23.490 772.030 24.100 ;
        RECT 772.870 23.490 783.530 24.100 ;
        RECT 784.370 23.490 795.030 24.100 ;
        RECT 795.870 23.490 806.530 24.100 ;
        RECT 807.370 23.490 818.030 24.100 ;
        RECT 818.870 23.490 829.530 24.100 ;
        RECT 830.370 23.490 841.030 24.100 ;
        RECT 841.870 23.490 852.530 24.100 ;
        RECT 853.370 23.490 864.030 24.100 ;
        RECT 864.870 23.490 875.530 24.100 ;
        RECT 876.370 23.490 887.030 24.100 ;
        RECT 887.870 23.490 898.530 24.100 ;
        RECT 899.370 23.490 910.030 24.100 ;
        RECT 910.870 23.490 921.530 24.100 ;
        RECT 922.370 23.490 933.030 24.100 ;
        RECT 933.870 23.490 944.530 24.100 ;
        RECT 945.370 23.490 956.030 24.100 ;
        RECT 956.870 23.490 967.530 24.100 ;
        RECT 968.370 23.490 979.030 24.100 ;
        RECT 979.870 23.490 990.530 24.100 ;
        RECT 991.370 23.490 1002.030 24.100 ;
        RECT 1002.870 23.490 1013.530 24.100 ;
        RECT 1014.370 23.490 1025.030 24.100 ;
        RECT 1025.870 23.490 1036.530 24.100 ;
        RECT 1037.370 23.490 1048.030 24.100 ;
        RECT 1048.870 23.490 1059.530 24.100 ;
        RECT 1060.370 23.490 1071.030 24.100 ;
        RECT 1071.870 23.490 1082.530 24.100 ;
        RECT 1083.370 23.490 1094.030 24.100 ;
        RECT 1094.870 23.490 1105.530 24.100 ;
        RECT 1106.370 23.490 1117.030 24.100 ;
        RECT 1117.870 23.490 1128.530 24.100 ;
        RECT 1129.370 23.490 1140.030 24.100 ;
        RECT 1140.870 23.490 1151.530 24.100 ;
        RECT 1152.370 23.490 1163.030 24.100 ;
        RECT 1163.870 23.490 1174.530 24.100 ;
        RECT 1175.370 23.490 1186.030 24.100 ;
        RECT 1186.870 23.490 1197.530 24.100 ;
        RECT 1198.370 23.490 1209.030 24.100 ;
        RECT 1209.870 23.490 1220.530 24.100 ;
        RECT 1221.370 23.490 1232.030 24.100 ;
        RECT 1232.870 23.490 1243.530 24.100 ;
        RECT 1244.370 23.490 1255.030 24.100 ;
        RECT 1255.870 23.490 1266.530 24.100 ;
        RECT 1267.370 23.490 1278.030 24.100 ;
        RECT 1278.870 23.490 1289.530 24.100 ;
        RECT 1290.370 23.490 1301.030 24.100 ;
        RECT 1301.870 23.490 1312.530 24.100 ;
        RECT 1313.370 23.490 1324.030 24.100 ;
        RECT 1324.870 23.490 1335.530 24.100 ;
        RECT 1336.370 23.490 1347.030 24.100 ;
        RECT 1347.870 23.490 1358.530 24.100 ;
        RECT 1359.370 23.490 1370.030 24.100 ;
        RECT 1370.870 23.490 1381.530 24.100 ;
        RECT 1382.370 23.490 1393.030 24.100 ;
        RECT 1393.870 23.490 1404.530 24.100 ;
        RECT 1405.370 23.490 1416.030 24.100 ;
        RECT 1416.870 23.490 1427.530 24.100 ;
        RECT 1428.370 23.490 1439.030 24.100 ;
        RECT 1439.870 23.490 1450.530 24.100 ;
        RECT 1451.370 23.490 1462.030 24.100 ;
        RECT 1462.870 23.490 1473.530 24.100 ;
        RECT 1474.370 23.490 1485.030 24.100 ;
        RECT 1485.870 23.490 1496.530 24.100 ;
        RECT 1497.370 23.490 1508.030 24.100 ;
        RECT 1508.870 23.490 1519.530 24.100 ;
        RECT 1520.370 23.490 1531.030 24.100 ;
        RECT 1531.870 23.490 1542.530 24.100 ;
        RECT 1543.370 23.490 1554.030 24.100 ;
        RECT 1554.870 23.490 1565.530 24.100 ;
        RECT 1566.370 23.490 1577.030 24.100 ;
        RECT 1577.870 23.490 1588.530 24.100 ;
        RECT 1589.370 23.490 1600.030 24.100 ;
        RECT 1600.870 23.490 1611.530 24.100 ;
        RECT 1612.370 23.490 1623.030 24.100 ;
        RECT 1623.870 23.490 1634.530 24.100 ;
        RECT 1635.370 23.490 1646.030 24.100 ;
        RECT 1646.870 23.490 1657.530 24.100 ;
        RECT 1658.370 23.490 1669.030 24.100 ;
        RECT 1669.870 23.490 1680.530 24.100 ;
        RECT 1681.370 23.490 1692.030 24.100 ;
        RECT 1692.870 23.490 1703.530 24.100 ;
        RECT 1704.370 23.490 1715.030 24.100 ;
        RECT 1715.870 23.490 1726.530 24.100 ;
        RECT 1727.370 23.490 1738.030 24.100 ;
        RECT 1738.870 23.490 1749.530 24.100 ;
        RECT 1750.370 23.490 1761.030 24.100 ;
        RECT 1761.870 23.490 1772.530 24.100 ;
        RECT 1773.370 23.490 1784.030 24.100 ;
        RECT 1784.870 23.490 1795.530 24.100 ;
        RECT 1796.370 23.490 1807.030 24.100 ;
        RECT 1807.870 23.490 1818.530 24.100 ;
        RECT 1819.370 23.490 1830.030 24.100 ;
        RECT 1830.870 23.490 1841.530 24.100 ;
        RECT 1842.370 23.490 1853.030 24.100 ;
        RECT 1853.870 23.490 1864.530 24.100 ;
        RECT 1865.370 23.490 1876.030 24.100 ;
        RECT 1876.870 23.490 1887.530 24.100 ;
        RECT 1888.370 23.490 1899.030 24.100 ;
        RECT 1899.870 23.490 1910.530 24.100 ;
        RECT 1911.370 23.490 1922.030 24.100 ;
        RECT 1922.870 23.490 1933.530 24.100 ;
        RECT 1934.370 23.490 1945.030 24.100 ;
        RECT 1945.870 23.490 1956.530 24.100 ;
        RECT 1957.370 23.490 1968.030 24.100 ;
        RECT 1968.870 23.490 1979.530 24.100 ;
        RECT 1980.370 23.490 1991.030 24.100 ;
        RECT 1991.870 23.490 2002.530 24.100 ;
        RECT 2003.370 23.490 2014.030 24.100 ;
        RECT 2014.870 23.490 2025.530 24.100 ;
        RECT 2026.370 23.490 2037.030 24.100 ;
        RECT 2037.870 23.490 2048.530 24.100 ;
        RECT 2049.370 23.490 2060.030 24.100 ;
        RECT 2060.870 23.490 2071.530 24.100 ;
        RECT 2072.370 23.490 2083.030 24.100 ;
        RECT 2083.870 23.490 2094.530 24.100 ;
        RECT 2095.370 23.490 2106.030 24.100 ;
        RECT 2106.870 23.490 2117.530 24.100 ;
        RECT 2118.370 23.490 2129.030 24.100 ;
        RECT 2129.870 23.490 2140.530 24.100 ;
        RECT 2141.370 23.490 2152.030 24.100 ;
        RECT 2152.870 23.490 2163.530 24.100 ;
        RECT 2164.370 23.490 2175.030 24.100 ;
        RECT 2175.870 23.490 2186.530 24.100 ;
        RECT 2187.370 23.490 2198.030 24.100 ;
        RECT 2198.870 23.490 2209.530 24.100 ;
        RECT 2210.370 23.490 2221.030 24.100 ;
        RECT 2221.870 23.490 2232.530 24.100 ;
        RECT 2233.370 23.490 2244.030 24.100 ;
        RECT 2244.870 23.490 2255.530 24.100 ;
        RECT 2256.370 23.490 2267.030 24.100 ;
        RECT 2267.870 23.490 2278.530 24.100 ;
        RECT 2279.370 23.490 2290.030 24.100 ;
        RECT 2290.870 23.490 2301.530 24.100 ;
        RECT 2302.370 23.490 2313.030 24.100 ;
        RECT 2313.870 23.490 2324.530 24.100 ;
        RECT 2325.370 23.490 2336.030 24.100 ;
        RECT 2336.870 23.490 2347.530 24.100 ;
        RECT 2348.370 23.490 2359.030 24.100 ;
        RECT 2359.870 23.490 2370.530 24.100 ;
        RECT 2371.370 23.490 2382.030 24.100 ;
        RECT 2382.870 23.490 2393.530 24.100 ;
        RECT 2394.370 23.490 2405.030 24.100 ;
        RECT 2405.870 23.490 2416.530 24.100 ;
        RECT 2417.370 23.490 2428.030 24.100 ;
        RECT 2428.870 23.490 2439.530 24.100 ;
        RECT 2440.370 23.490 2451.030 24.100 ;
        RECT 2451.870 23.490 2462.530 24.100 ;
        RECT 2463.370 23.490 2474.030 24.100 ;
        RECT 2474.870 23.490 2485.530 24.100 ;
        RECT 2486.370 23.490 2497.030 24.100 ;
        RECT 2497.870 23.490 2508.530 24.100 ;
      LAYER met3 ;
        RECT 29.180 2833.340 2516.180 2870.105 ;
        RECT 29.580 2831.940 2516.180 2833.340 ;
        RECT 29.180 2821.100 2516.180 2831.940 ;
        RECT 29.180 2819.700 2515.780 2821.100 ;
        RECT 29.180 2734.740 2516.180 2819.700 ;
        RECT 29.580 2733.340 2516.180 2734.740 ;
        RECT 29.180 2702.100 2516.180 2733.340 ;
        RECT 29.180 2700.700 2515.780 2702.100 ;
        RECT 29.180 2636.140 2516.180 2700.700 ;
        RECT 29.580 2634.740 2516.180 2636.140 ;
        RECT 29.180 2583.100 2516.180 2634.740 ;
        RECT 29.180 2581.700 2515.780 2583.100 ;
        RECT 29.180 2537.540 2516.180 2581.700 ;
        RECT 29.580 2536.140 2516.180 2537.540 ;
        RECT 29.180 2464.100 2516.180 2536.140 ;
        RECT 29.180 2462.700 2515.780 2464.100 ;
        RECT 29.180 2438.940 2516.180 2462.700 ;
        RECT 29.580 2437.540 2516.180 2438.940 ;
        RECT 29.180 2345.100 2516.180 2437.540 ;
        RECT 29.180 2343.700 2515.780 2345.100 ;
        RECT 29.180 2340.340 2516.180 2343.700 ;
        RECT 29.580 2338.940 2516.180 2340.340 ;
        RECT 29.180 2241.740 2516.180 2338.940 ;
        RECT 29.580 2240.340 2516.180 2241.740 ;
        RECT 29.180 2226.100 2516.180 2240.340 ;
        RECT 29.180 2224.700 2515.780 2226.100 ;
        RECT 29.180 2143.140 2516.180 2224.700 ;
        RECT 29.580 2141.740 2516.180 2143.140 ;
        RECT 29.180 2107.100 2516.180 2141.740 ;
        RECT 29.180 2105.700 2515.780 2107.100 ;
        RECT 29.180 2044.540 2516.180 2105.700 ;
        RECT 29.580 2043.140 2516.180 2044.540 ;
        RECT 29.180 1988.100 2516.180 2043.140 ;
        RECT 29.180 1986.700 2515.780 1988.100 ;
        RECT 29.180 1945.940 2516.180 1986.700 ;
        RECT 29.580 1944.540 2516.180 1945.940 ;
        RECT 29.180 1869.100 2516.180 1944.540 ;
        RECT 29.180 1867.700 2515.780 1869.100 ;
        RECT 29.180 1847.340 2516.180 1867.700 ;
        RECT 29.580 1845.940 2516.180 1847.340 ;
        RECT 29.180 1750.100 2516.180 1845.940 ;
        RECT 29.180 1748.740 2515.780 1750.100 ;
        RECT 29.580 1748.700 2515.780 1748.740 ;
        RECT 29.580 1747.340 2516.180 1748.700 ;
        RECT 29.180 1650.140 2516.180 1747.340 ;
        RECT 29.580 1648.740 2516.180 1650.140 ;
        RECT 29.180 1631.100 2516.180 1648.740 ;
        RECT 29.180 1629.700 2515.780 1631.100 ;
        RECT 29.180 1551.540 2516.180 1629.700 ;
        RECT 29.580 1550.140 2516.180 1551.540 ;
        RECT 29.180 1512.100 2516.180 1550.140 ;
        RECT 29.180 1510.700 2515.780 1512.100 ;
        RECT 29.180 1452.940 2516.180 1510.700 ;
        RECT 29.580 1451.540 2516.180 1452.940 ;
        RECT 29.180 1393.100 2516.180 1451.540 ;
        RECT 29.180 1391.700 2515.780 1393.100 ;
        RECT 29.180 1354.340 2516.180 1391.700 ;
        RECT 29.580 1352.940 2516.180 1354.340 ;
        RECT 29.180 1274.100 2516.180 1352.940 ;
        RECT 29.180 1272.700 2515.780 1274.100 ;
        RECT 29.180 1255.740 2516.180 1272.700 ;
        RECT 29.580 1254.340 2516.180 1255.740 ;
        RECT 29.180 1157.140 2516.180 1254.340 ;
        RECT 29.580 1155.740 2516.180 1157.140 ;
        RECT 29.180 1155.100 2516.180 1155.740 ;
        RECT 29.180 1153.700 2515.780 1155.100 ;
        RECT 29.180 1058.540 2516.180 1153.700 ;
        RECT 29.580 1057.140 2516.180 1058.540 ;
        RECT 29.180 1036.100 2516.180 1057.140 ;
        RECT 29.180 1034.700 2515.780 1036.100 ;
        RECT 29.180 959.940 2516.180 1034.700 ;
        RECT 29.580 958.540 2516.180 959.940 ;
        RECT 29.180 917.100 2516.180 958.540 ;
        RECT 29.180 915.700 2515.780 917.100 ;
        RECT 29.180 861.340 2516.180 915.700 ;
        RECT 29.580 859.940 2516.180 861.340 ;
        RECT 29.180 798.100 2516.180 859.940 ;
        RECT 29.180 796.700 2515.780 798.100 ;
        RECT 29.180 762.740 2516.180 796.700 ;
        RECT 29.580 761.340 2516.180 762.740 ;
        RECT 29.180 679.100 2516.180 761.340 ;
        RECT 29.180 677.700 2515.780 679.100 ;
        RECT 29.180 664.140 2516.180 677.700 ;
        RECT 29.580 662.740 2516.180 664.140 ;
        RECT 29.180 565.540 2516.180 662.740 ;
        RECT 29.580 564.140 2516.180 565.540 ;
        RECT 29.180 560.100 2516.180 564.140 ;
        RECT 29.180 558.700 2515.780 560.100 ;
        RECT 29.180 466.940 2516.180 558.700 ;
        RECT 29.580 465.540 2516.180 466.940 ;
        RECT 29.180 441.100 2516.180 465.540 ;
        RECT 29.180 439.700 2515.780 441.100 ;
        RECT 29.180 368.340 2516.180 439.700 ;
        RECT 29.580 366.940 2516.180 368.340 ;
        RECT 29.180 322.100 2516.180 366.940 ;
        RECT 29.180 320.700 2515.780 322.100 ;
        RECT 29.180 269.740 2516.180 320.700 ;
        RECT 29.580 268.340 2516.180 269.740 ;
        RECT 29.180 203.100 2516.180 268.340 ;
        RECT 29.180 201.700 2515.780 203.100 ;
        RECT 29.180 171.140 2516.180 201.700 ;
        RECT 29.580 169.740 2516.180 171.140 ;
        RECT 29.180 84.100 2516.180 169.740 ;
        RECT 29.180 82.700 2515.780 84.100 ;
        RECT 29.180 72.540 2516.180 82.700 ;
        RECT 29.580 71.675 2516.180 72.540 ;
      LAYER met4 ;
        RECT 92.895 105.460 2465.460 2870.180 ;
  END
END fpga_core
END LIBRARY

